`define iteration_times 40 module bp_256_128 #(	parameter integer BIT = 8)(	input clk,	input rst_n,	input start,	output reg en_busy,	input [BIT - 1:0] LLR_1,	input [BIT - 1:0] LLR_2,	input [BIT - 1:0] LLR_3,	input [BIT - 1:0] LLR_4,	input [BIT - 1:0] LLR_5,	input [BIT - 1:0] LLR_6,	input [BIT - 1:0] LLR_7,	input [BIT - 1:0] LLR_8,	input [BIT - 1:0] LLR_9,	input [BIT - 1:0] LLR_10,	input [BIT - 1:0] LLR_11,	input [BIT - 1:0] LLR_12,	input [BIT - 1:0] LLR_13,	input [BIT - 1:0] LLR_14,	input [BIT - 1:0] LLR_15,	input [BIT - 1:0] LLR_16,	input [BIT - 1:0] LLR_17,	input [BIT - 1:0] LLR_18,	input [BIT - 1:0] LLR_19,	input [BIT - 1:0] LLR_20,	input [BIT - 1:0] LLR_21,	input [BIT - 1:0] LLR_22,	input [BIT - 1:0] LLR_23,	input [BIT - 1:0] LLR_24,	input [BIT - 1:0] LLR_25,	input [BIT - 1:0] LLR_26,	input [BIT - 1:0] LLR_27,	input [BIT - 1:0] LLR_28,	input [BIT - 1:0] LLR_29,	input [BIT - 1:0] LLR_30,	input [BIT - 1:0] LLR_31,	input [BIT - 1:0] LLR_32,	input [BIT - 1:0] LLR_33,	input [BIT - 1:0] LLR_34,	input [BIT - 1:0] LLR_35,	input [BIT - 1:0] LLR_36,	input [BIT - 1:0] LLR_37,	input [BIT - 1:0] LLR_38,	input [BIT - 1:0] LLR_39,	input [BIT - 1:0] LLR_40,	input [BIT - 1:0] LLR_41,	input [BIT - 1:0] LLR_42,	input [BIT - 1:0] LLR_43,	input [BIT - 1:0] LLR_44,	input [BIT - 1:0] LLR_45,	input [BIT - 1:0] LLR_46,	input [BIT - 1:0] LLR_47,	input [BIT - 1:0] LLR_48,	input [BIT - 1:0] LLR_49,	input [BIT - 1:0] LLR_50,	input [BIT - 1:0] LLR_51,	input [BIT - 1:0] LLR_52,	input [BIT - 1:0] LLR_53,	input [BIT - 1:0] LLR_54,	input [BIT - 1:0] LLR_55,	input [BIT - 1:0] LLR_56,	input [BIT - 1:0] LLR_57,	input [BIT - 1:0] LLR_58,	input [BIT - 1:0] LLR_59,	input [BIT - 1:0] LLR_60,	input [BIT - 1:0] LLR_61,	input [BIT - 1:0] LLR_62,	input [BIT - 1:0] LLR_63,	input [BIT - 1:0] LLR_64,	input [BIT - 1:0] LLR_65,	input [BIT - 1:0] LLR_66,	input [BIT - 1:0] LLR_67,	input [BIT - 1:0] LLR_68,	input [BIT - 1:0] LLR_69,	input [BIT - 1:0] LLR_70,	input [BIT - 1:0] LLR_71,	input [BIT - 1:0] LLR_72,	input [BIT - 1:0] LLR_73,	input [BIT - 1:0] LLR_74,	input [BIT - 1:0] LLR_75,	input [BIT - 1:0] LLR_76,	input [BIT - 1:0] LLR_77,	input [BIT - 1:0] LLR_78,	input [BIT - 1:0] LLR_79,	input [BIT - 1:0] LLR_80,	input [BIT - 1:0] LLR_81,	input [BIT - 1:0] LLR_82,	input [BIT - 1:0] LLR_83,	input [BIT - 1:0] LLR_84,	input [BIT - 1:0] LLR_85,	input [BIT - 1:0] LLR_86,	input [BIT - 1:0] LLR_87,	input [BIT - 1:0] LLR_88,	input [BIT - 1:0] LLR_89,	input [BIT - 1:0] LLR_90,	input [BIT - 1:0] LLR_91,	input [BIT - 1:0] LLR_92,	input [BIT - 1:0] LLR_93,	input [BIT - 1:0] LLR_94,	input [BIT - 1:0] LLR_95,	input [BIT - 1:0] LLR_96,	input [BIT - 1:0] LLR_97,	input [BIT - 1:0] LLR_98,	input [BIT - 1:0] LLR_99,	input [BIT - 1:0] LLR_100,	input [BIT - 1:0] LLR_101,	input [BIT - 1:0] LLR_102,	input [BIT - 1:0] LLR_103,	input [BIT - 1:0] LLR_104,	input [BIT - 1:0] LLR_105,	input [BIT - 1:0] LLR_106,	input [BIT - 1:0] LLR_107,	input [BIT - 1:0] LLR_108,	input [BIT - 1:0] LLR_109,	input [BIT - 1:0] LLR_110,	input [BIT - 1:0] LLR_111,	input [BIT - 1:0] LLR_112,	input [BIT - 1:0] LLR_113,	input [BIT - 1:0] LLR_114,	input [BIT - 1:0] LLR_115,	input [BIT - 1:0] LLR_116,	input [BIT - 1:0] LLR_117,	input [BIT - 1:0] LLR_118,	input [BIT - 1:0] LLR_119,	input [BIT - 1:0] LLR_120,	input [BIT - 1:0] LLR_121,	input [BIT - 1:0] LLR_122,	input [BIT - 1:0] LLR_123,	input [BIT - 1:0] LLR_124,	input [BIT - 1:0] LLR_125,	input [BIT - 1:0] LLR_126,	input [BIT - 1:0] LLR_127,	input [BIT - 1:0] LLR_128,	input [BIT - 1:0] LLR_129,	input [BIT - 1:0] LLR_130,	input [BIT - 1:0] LLR_131,	input [BIT - 1:0] LLR_132,	input [BIT - 1:0] LLR_133,	input [BIT - 1:0] LLR_134,	input [BIT - 1:0] LLR_135,	input [BIT - 1:0] LLR_136,	input [BIT - 1:0] LLR_137,	input [BIT - 1:0] LLR_138,	input [BIT - 1:0] LLR_139,	input [BIT - 1:0] LLR_140,	input [BIT - 1:0] LLR_141,	input [BIT - 1:0] LLR_142,	input [BIT - 1:0] LLR_143,	input [BIT - 1:0] LLR_144,	input [BIT - 1:0] LLR_145,	input [BIT - 1:0] LLR_146,	input [BIT - 1:0] LLR_147,	input [BIT - 1:0] LLR_148,	input [BIT - 1:0] LLR_149,	input [BIT - 1:0] LLR_150,	input [BIT - 1:0] LLR_151,	input [BIT - 1:0] LLR_152,	input [BIT - 1:0] LLR_153,	input [BIT - 1:0] LLR_154,	input [BIT - 1:0] LLR_155,	input [BIT - 1:0] LLR_156,	input [BIT - 1:0] LLR_157,	input [BIT - 1:0] LLR_158,	input [BIT - 1:0] LLR_159,	input [BIT - 1:0] LLR_160,	input [BIT - 1:0] LLR_161,	input [BIT - 1:0] LLR_162,	input [BIT - 1:0] LLR_163,	input [BIT - 1:0] LLR_164,	input [BIT - 1:0] LLR_165,	input [BIT - 1:0] LLR_166,	input [BIT - 1:0] LLR_167,	input [BIT - 1:0] LLR_168,	input [BIT - 1:0] LLR_169,	input [BIT - 1:0] LLR_170,	input [BIT - 1:0] LLR_171,	input [BIT - 1:0] LLR_172,	input [BIT - 1:0] LLR_173,	input [BIT - 1:0] LLR_174,	input [BIT - 1:0] LLR_175,	input [BIT - 1:0] LLR_176,	input [BIT - 1:0] LLR_177,	input [BIT - 1:0] LLR_178,	input [BIT - 1:0] LLR_179,	input [BIT - 1:0] LLR_180,	input [BIT - 1:0] LLR_181,	input [BIT - 1:0] LLR_182,	input [BIT - 1:0] LLR_183,	input [BIT - 1:0] LLR_184,	input [BIT - 1:0] LLR_185,	input [BIT - 1:0] LLR_186,	input [BIT - 1:0] LLR_187,	input [BIT - 1:0] LLR_188,	input [BIT - 1:0] LLR_189,	input [BIT - 1:0] LLR_190,	input [BIT - 1:0] LLR_191,	input [BIT - 1:0] LLR_192,	input [BIT - 1:0] LLR_193,	input [BIT - 1:0] LLR_194,	input [BIT - 1:0] LLR_195,	input [BIT - 1:0] LLR_196,	input [BIT - 1:0] LLR_197,	input [BIT - 1:0] LLR_198,	input [BIT - 1:0] LLR_199,	input [BIT - 1:0] LLR_200,	input [BIT - 1:0] LLR_201,	input [BIT - 1:0] LLR_202,	input [BIT - 1:0] LLR_203,	input [BIT - 1:0] LLR_204,	input [BIT - 1:0] LLR_205,	input [BIT - 1:0] LLR_206,	input [BIT - 1:0] LLR_207,	input [BIT - 1:0] LLR_208,	input [BIT - 1:0] LLR_209,	input [BIT - 1:0] LLR_210,	input [BIT - 1:0] LLR_211,	input [BIT - 1:0] LLR_212,	input [BIT - 1:0] LLR_213,	input [BIT - 1:0] LLR_214,	input [BIT - 1:0] LLR_215,	input [BIT - 1:0] LLR_216,	input [BIT - 1:0] LLR_217,	input [BIT - 1:0] LLR_218,	input [BIT - 1:0] LLR_219,	input [BIT - 1:0] LLR_220,	input [BIT - 1:0] LLR_221,	input [BIT - 1:0] LLR_222,	input [BIT - 1:0] LLR_223,	input [BIT - 1:0] LLR_224,	input [BIT - 1:0] LLR_225,	input [BIT - 1:0] LLR_226,	input [BIT - 1:0] LLR_227,	input [BIT - 1:0] LLR_228,	input [BIT - 1:0] LLR_229,	input [BIT - 1:0] LLR_230,	input [BIT - 1:0] LLR_231,	input [BIT - 1:0] LLR_232,	input [BIT - 1:0] LLR_233,	input [BIT - 1:0] LLR_234,	input [BIT - 1:0] LLR_235,	input [BIT - 1:0] LLR_236,	input [BIT - 1:0] LLR_237,	input [BIT - 1:0] LLR_238,	input [BIT - 1:0] LLR_239,	input [BIT - 1:0] LLR_240,	input [BIT - 1:0] LLR_241,	input [BIT - 1:0] LLR_242,	input [BIT - 1:0] LLR_243,	input [BIT - 1:0] LLR_244,	input [BIT - 1:0] LLR_245,	input [BIT - 1:0] LLR_246,	input [BIT - 1:0] LLR_247,	input [BIT - 1:0] LLR_248,	input [BIT - 1:0] LLR_249,	input [BIT - 1:0] LLR_250,	input [BIT - 1:0] LLR_251,	input [BIT - 1:0] LLR_252,	input [BIT - 1:0] LLR_253,	input [BIT - 1:0] LLR_254,	input [BIT - 1:0] LLR_255,	input [BIT - 1:0] LLR_256,	output reg [BIT - 1:0] OUT_1,	output reg [BIT - 1:0] OUT_2,	output reg [BIT - 1:0] OUT_3,	output reg [BIT - 1:0] OUT_4,	output reg [BIT - 1:0] OUT_5,	output reg [BIT - 1:0] OUT_6,	output reg [BIT - 1:0] OUT_7,	output reg [BIT - 1:0] OUT_8,	output reg [BIT - 1:0] OUT_9,	output reg [BIT - 1:0] OUT_10,	output reg [BIT - 1:0] OUT_11,	output reg [BIT - 1:0] OUT_12,	output reg [BIT - 1:0] OUT_13,	output reg [BIT - 1:0] OUT_14,	output reg [BIT - 1:0] OUT_15,	output reg [BIT - 1:0] OUT_16,	output reg [BIT - 1:0] OUT_17,	output reg [BIT - 1:0] OUT_18,	output reg [BIT - 1:0] OUT_19,	output reg [BIT - 1:0] OUT_20,	output reg [BIT - 1:0] OUT_21,	output reg [BIT - 1:0] OUT_22,	output reg [BIT - 1:0] OUT_23,	output reg [BIT - 1:0] OUT_24,	output reg [BIT - 1:0] OUT_25,	output reg [BIT - 1:0] OUT_26,	output reg [BIT - 1:0] OUT_27,	output reg [BIT - 1:0] OUT_28,	output reg [BIT - 1:0] OUT_29,	output reg [BIT - 1:0] OUT_30,	output reg [BIT - 1:0] OUT_31,	output reg [BIT - 1:0] OUT_32,	output reg [BIT - 1:0] OUT_33,	output reg [BIT - 1:0] OUT_34,	output reg [BIT - 1:0] OUT_35,	output reg [BIT - 1:0] OUT_36,	output reg [BIT - 1:0] OUT_37,	output reg [BIT - 1:0] OUT_38,	output reg [BIT - 1:0] OUT_39,	output reg [BIT - 1:0] OUT_40,	output reg [BIT - 1:0] OUT_41,	output reg [BIT - 1:0] OUT_42,	output reg [BIT - 1:0] OUT_43,	output reg [BIT - 1:0] OUT_44,	output reg [BIT - 1:0] OUT_45,	output reg [BIT - 1:0] OUT_46,	output reg [BIT - 1:0] OUT_47,	output reg [BIT - 1:0] OUT_48,	output reg [BIT - 1:0] OUT_49,	output reg [BIT - 1:0] OUT_50,	output reg [BIT - 1:0] OUT_51,	output reg [BIT - 1:0] OUT_52,	output reg [BIT - 1:0] OUT_53,	output reg [BIT - 1:0] OUT_54,	output reg [BIT - 1:0] OUT_55,	output reg [BIT - 1:0] OUT_56,	output reg [BIT - 1:0] OUT_57,	output reg [BIT - 1:0] OUT_58,	output reg [BIT - 1:0] OUT_59,	output reg [BIT - 1:0] OUT_60,	output reg [BIT - 1:0] OUT_61,	output reg [BIT - 1:0] OUT_62,	output reg [BIT - 1:0] OUT_63,	output reg [BIT - 1:0] OUT_64,	output reg [BIT - 1:0] OUT_65,	output reg [BIT - 1:0] OUT_66,	output reg [BIT - 1:0] OUT_67,	output reg [BIT - 1:0] OUT_68,	output reg [BIT - 1:0] OUT_69,	output reg [BIT - 1:0] OUT_70,	output reg [BIT - 1:0] OUT_71,	output reg [BIT - 1:0] OUT_72,	output reg [BIT - 1:0] OUT_73,	output reg [BIT - 1:0] OUT_74,	output reg [BIT - 1:0] OUT_75,	output reg [BIT - 1:0] OUT_76,	output reg [BIT - 1:0] OUT_77,	output reg [BIT - 1:0] OUT_78,	output reg [BIT - 1:0] OUT_79,	output reg [BIT - 1:0] OUT_80,	output reg [BIT - 1:0] OUT_81,	output reg [BIT - 1:0] OUT_82,	output reg [BIT - 1:0] OUT_83,	output reg [BIT - 1:0] OUT_84,	output reg [BIT - 1:0] OUT_85,	output reg [BIT - 1:0] OUT_86,	output reg [BIT - 1:0] OUT_87,	output reg [BIT - 1:0] OUT_88,	output reg [BIT - 1:0] OUT_89,	output reg [BIT - 1:0] OUT_90,	output reg [BIT - 1:0] OUT_91,	output reg [BIT - 1:0] OUT_92,	output reg [BIT - 1:0] OUT_93,	output reg [BIT - 1:0] OUT_94,	output reg [BIT - 1:0] OUT_95,	output reg [BIT - 1:0] OUT_96,	output reg [BIT - 1:0] OUT_97,	output reg [BIT - 1:0] OUT_98,	output reg [BIT - 1:0] OUT_99,	output reg [BIT - 1:0] OUT_100,	output reg [BIT - 1:0] OUT_101,	output reg [BIT - 1:0] OUT_102,	output reg [BIT - 1:0] OUT_103,	output reg [BIT - 1:0] OUT_104,	output reg [BIT - 1:0] OUT_105,	output reg [BIT - 1:0] OUT_106,	output reg [BIT - 1:0] OUT_107,	output reg [BIT - 1:0] OUT_108,	output reg [BIT - 1:0] OUT_109,	output reg [BIT - 1:0] OUT_110,	output reg [BIT - 1:0] OUT_111,	output reg [BIT - 1:0] OUT_112,	output reg [BIT - 1:0] OUT_113,	output reg [BIT - 1:0] OUT_114,	output reg [BIT - 1:0] OUT_115,	output reg [BIT - 1:0] OUT_116,	output reg [BIT - 1:0] OUT_117,	output reg [BIT - 1:0] OUT_118,	output reg [BIT - 1:0] OUT_119,	output reg [BIT - 1:0] OUT_120,	output reg [BIT - 1:0] OUT_121,	output reg [BIT - 1:0] OUT_122,	output reg [BIT - 1:0] OUT_123,	output reg [BIT - 1:0] OUT_124,	output reg [BIT - 1:0] OUT_125,	output reg [BIT - 1:0] OUT_126,	output reg [BIT - 1:0] OUT_127,	output reg [BIT - 1:0] OUT_128,	output reg [BIT - 1:0] OUT_129,	output reg [BIT - 1:0] OUT_130,	output reg [BIT - 1:0] OUT_131,	output reg [BIT - 1:0] OUT_132,	output reg [BIT - 1:0] OUT_133,	output reg [BIT - 1:0] OUT_134,	output reg [BIT - 1:0] OUT_135,	output reg [BIT - 1:0] OUT_136,	output reg [BIT - 1:0] OUT_137,	output reg [BIT - 1:0] OUT_138,	output reg [BIT - 1:0] OUT_139,	output reg [BIT - 1:0] OUT_140,	output reg [BIT - 1:0] OUT_141,	output reg [BIT - 1:0] OUT_142,	output reg [BIT - 1:0] OUT_143,	output reg [BIT - 1:0] OUT_144,	output reg [BIT - 1:0] OUT_145,	output reg [BIT - 1:0] OUT_146,	output reg [BIT - 1:0] OUT_147,	output reg [BIT - 1:0] OUT_148,	output reg [BIT - 1:0] OUT_149,	output reg [BIT - 1:0] OUT_150,	output reg [BIT - 1:0] OUT_151,	output reg [BIT - 1:0] OUT_152,	output reg [BIT - 1:0] OUT_153,	output reg [BIT - 1:0] OUT_154,	output reg [BIT - 1:0] OUT_155,	output reg [BIT - 1:0] OUT_156,	output reg [BIT - 1:0] OUT_157,	output reg [BIT - 1:0] OUT_158,	output reg [BIT - 1:0] OUT_159,	output reg [BIT - 1:0] OUT_160,	output reg [BIT - 1:0] OUT_161,	output reg [BIT - 1:0] OUT_162,	output reg [BIT - 1:0] OUT_163,	output reg [BIT - 1:0] OUT_164,	output reg [BIT - 1:0] OUT_165,	output reg [BIT - 1:0] OUT_166,	output reg [BIT - 1:0] OUT_167,	output reg [BIT - 1:0] OUT_168,	output reg [BIT - 1:0] OUT_169,	output reg [BIT - 1:0] OUT_170,	output reg [BIT - 1:0] OUT_171,	output reg [BIT - 1:0] OUT_172,	output reg [BIT - 1:0] OUT_173,	output reg [BIT - 1:0] OUT_174,	output reg [BIT - 1:0] OUT_175,	output reg [BIT - 1:0] OUT_176,	output reg [BIT - 1:0] OUT_177,	output reg [BIT - 1:0] OUT_178,	output reg [BIT - 1:0] OUT_179,	output reg [BIT - 1:0] OUT_180,	output reg [BIT - 1:0] OUT_181,	output reg [BIT - 1:0] OUT_182,	output reg [BIT - 1:0] OUT_183,	output reg [BIT - 1:0] OUT_184,	output reg [BIT - 1:0] OUT_185,	output reg [BIT - 1:0] OUT_186,	output reg [BIT - 1:0] OUT_187,	output reg [BIT - 1:0] OUT_188,	output reg [BIT - 1:0] OUT_189,	output reg [BIT - 1:0] OUT_190,	output reg [BIT - 1:0] OUT_191,	output reg [BIT - 1:0] OUT_192,	output reg [BIT - 1:0] OUT_193,	output reg [BIT - 1:0] OUT_194,	output reg [BIT - 1:0] OUT_195,	output reg [BIT - 1:0] OUT_196,	output reg [BIT - 1:0] OUT_197,	output reg [BIT - 1:0] OUT_198,	output reg [BIT - 1:0] OUT_199,	output reg [BIT - 1:0] OUT_200,	output reg [BIT - 1:0] OUT_201,	output reg [BIT - 1:0] OUT_202,	output reg [BIT - 1:0] OUT_203,	output reg [BIT - 1:0] OUT_204,	output reg [BIT - 1:0] OUT_205,	output reg [BIT - 1:0] OUT_206,	output reg [BIT - 1:0] OUT_207,	output reg [BIT - 1:0] OUT_208,	output reg [BIT - 1:0] OUT_209,	output reg [BIT - 1:0] OUT_210,	output reg [BIT - 1:0] OUT_211,	output reg [BIT - 1:0] OUT_212,	output reg [BIT - 1:0] OUT_213,	output reg [BIT - 1:0] OUT_214,	output reg [BIT - 1:0] OUT_215,	output reg [BIT - 1:0] OUT_216,	output reg [BIT - 1:0] OUT_217,	output reg [BIT - 1:0] OUT_218,	output reg [BIT - 1:0] OUT_219,	output reg [BIT - 1:0] OUT_220,	output reg [BIT - 1:0] OUT_221,	output reg [BIT - 1:0] OUT_222,	output reg [BIT - 1:0] OUT_223,	output reg [BIT - 1:0] OUT_224,	output reg [BIT - 1:0] OUT_225,	output reg [BIT - 1:0] OUT_226,	output reg [BIT - 1:0] OUT_227,	output reg [BIT - 1:0] OUT_228,	output reg [BIT - 1:0] OUT_229,	output reg [BIT - 1:0] OUT_230,	output reg [BIT - 1:0] OUT_231,	output reg [BIT - 1:0] OUT_232,	output reg [BIT - 1:0] OUT_233,	output reg [BIT - 1:0] OUT_234,	output reg [BIT - 1:0] OUT_235,	output reg [BIT - 1:0] OUT_236,	output reg [BIT - 1:0] OUT_237,	output reg [BIT - 1:0] OUT_238,	output reg [BIT - 1:0] OUT_239,	output reg [BIT - 1:0] OUT_240,	output reg [BIT - 1:0] OUT_241,	output reg [BIT - 1:0] OUT_242,	output reg [BIT - 1:0] OUT_243,	output reg [BIT - 1:0] OUT_244,	output reg [BIT - 1:0] OUT_245,	output reg [BIT - 1:0] OUT_246,	output reg [BIT - 1:0] OUT_247,	output reg [BIT - 1:0] OUT_248,	output reg [BIT - 1:0] OUT_249,	output reg [BIT - 1:0] OUT_250,	output reg [BIT - 1:0] OUT_251,	output reg [BIT - 1:0] OUT_252,	output reg [BIT - 1:0] OUT_253,	output reg [BIT - 1:0] OUT_254,	output reg [BIT - 1:0] OUT_255,	output reg [BIT - 1:0] OUT_256);	integer x, y;
	reg [BIT - 1:0] inform_R [256-1:0][9-1:0];	reg [BIT - 1:0] inform_L [256-1:0][9-1:0];	localparam IDLE = 2'b00;	localparam BUSY_LEFT = 2'b01;	localparam BUSY_RIGHT = 2'b10;	reg [1:0] bp_state,bp_next_state;	reg [8-1:0] cell_enable,w2r;	reg left_over_flag,right_over_flag,init_over_flag;	wire bp_over_flag;	reg [6:0]itera_time;
	always @(posedge clk or negedge rst_n) begin		if (!rst_n) begin			bp_state <= IDLE;		end		else begin			bp_state <= bp_next_state;		end	end
	always @(*) begin		case (bp_state)			IDLE:			if (init_over_flag) begin				bp_next_state <= BUSY_LEFT;			end			else begin				bp_next_state <= IDLE;			end
			BUSY_LEFT:			if (left_over_flag) begin				bp_next_state <= BUSY_RIGHT;			end			else begin				 bp_next_state <= BUSY_LEFT;			end
			BUSY_RIGHT:			if (bp_over_flag) begin				bp_next_state <= IDLE;			end			else if (right_over_flag) begin				bp_next_state <= BUSY_LEFT;			end			else begin				 bp_next_state <= BUSY_RIGHT;			end
			default: bp_next_state <= IDLE;		endcase	end
	reg [1:0] clk_counter;
	always @(posedge clk) begin		case (bp_next_state)			IDLE:			begin				left_over_flag <= 0;				right_over_flag <= 0;				itera_time <= 7'b0;				clk_counter <= 2'b0;				if (start) begin					cell_enable <=8'b1;					w2r <= 8;					init_over_flag <= 1;					en_busy <= 1;				end				else begin					cell_enable <=8'b0;					w2r <= 0;					init_over_flag <= 0;					en_busy <= 0;				end			end
			BUSY_LEFT:			begin				init_over_flag <= 0;				en_busy <= 1;				right_over_flag <= 0;				if (clk_counter == 2'b11) begin					clk_counter <= 2'b00;					if (cell_enable == 128) begin						left_over_flag <= 1;						cell_enable <= cell_enable >> 1;						w2r <= w2r + 1;					end					else begin						left_over_flag <= 0;						cell_enable <= cell_enable << 1;						w2r <= w2r - 1;					end				end				else begin					clk_counter <= clk_counter + 1;				end			end
			BUSY_RIGHT:			begin				en_busy <= 1;				left_over_flag <= 0;				if (clk_counter == 2'b11) begin					clk_counter <= 2'b00;					if (cell_enable == 1) begin						right_over_flag <= 1;						itera_time <= itera_time + 1;						cell_enable <= cell_enable << 1;						w2r <= w2r - 1;					end					else begin						right_over_flag <= 0;						cell_enable <= cell_enable >> 1;						w2r <= w2r + 1;					end				end				else begin					clk_counter <= clk_counter + 1;				end			end
			default:			begin				left_over_flag <= 0;				right_over_flag <= 0;				itera_time <= 7'b0;				clk_counter <= 2'b0;				if (start) begin					cell_enable <=8'b1;					w2r <= 8;					init_over_flag <= 1;					en_busy <= 1;				end				else begin					cell_enable <=8'b0;					w2r <= 0;					init_over_flag <= 0;					en_busy <= 0;				end			end
		endcase	end
	reg[BIT - 1:0] r_cell_reg[256-1:0];	reg[BIT - 1:0] l_cell_reg[256-1:0];	wire[BIT - 1:0] r_cell_wire[256-1:0];	wire[BIT - 1:0] l_cell_wire[256-1:0];
	always @(posedge clk) begin		case (bp_next_state)			IDLE:			begin				if (start) begin					inform_R [0][0] <= 8'b0111_1111;					inform_R [1][0] <= 8'b0111_1111;					inform_R [2][0] <= 8'b0111_1111;					inform_R [3][0] <= 8'b0111_1111;					inform_R [4][0] <= 8'b0111_1111;					inform_R [5][0] <= 8'b0111_1111;					inform_R [6][0] <= 8'b0111_1111;					inform_R [7][0] <= 8'b0111_1111;					inform_R [8][0] <= 8'b0111_1111;					inform_R [9][0] <= 8'b0111_1111;					inform_R [10][0] <= 8'b0111_1111;					inform_R [11][0] <= 8'b0111_1111;					inform_R [12][0] <= 8'b0111_1111;					inform_R [13][0] <= 8'b0111_1111;					inform_R [14][0] <= 8'b0111_1111;					inform_R [15][0] <= 8'b0111_1111;					inform_R [16][0] <= 8'b0111_1111;					inform_R [17][0] <= 8'b0111_1111;					inform_R [18][0] <= 8'b0111_1111;					inform_R [19][0] <= 8'b0111_1111;					inform_R [20][0] <= 8'b0111_1111;					inform_R [21][0] <= 8'b0111_1111;					inform_R [22][0] <= 8'b0111_1111;					inform_R [23][0] <= 8'b0111_1111;					inform_R [24][0] <= 8'b0111_1111;					inform_R [25][0] <= 8'b0111_1111;					inform_R [26][0] <= 8'b0111_1111;					inform_R [27][0] <= 8'b0111_1111;					inform_R [28][0] <= 8'b0111_1111;					inform_R [29][0] <= 8'b0111_1111;					inform_R [30][0] <= 8'b0111_1111;					inform_R [31][0] <= 8'b0111_1111;					inform_R [32][0] <= 8'b0111_1111;					inform_R [33][0] <= 8'b0111_1111;					inform_R [34][0] <= 8'b0111_1111;					inform_R [35][0] <= 8'b0111_1111;					inform_R [36][0] <= 8'b0111_1111;					inform_R [37][0] <= 8'b0111_1111;					inform_R [38][0] <= 8'b0111_1111;					inform_R [39][0] <= 8'b0111_1111;					inform_R [40][0] <= 8'b0111_1111;					inform_R [41][0] <= 8'b0111_1111;					inform_R [42][0] <= 8'b0111_1111;					inform_R [43][0] <= 8'b0111_1111;					inform_R [44][0] <= 8'b0111_1111;					inform_R [45][0] <= 8'b0111_1111;					inform_R [46][0] <= 8'b0111_1111;					inform_R [47][0] <= 8'b0111_1111;					inform_R [48][0] <= 8'b0111_1111;					inform_R [49][0] <= 8'b0111_1111;					inform_R [50][0] <= 8'b0111_1111;					inform_R [51][0] <= 8'b0111_1111;					inform_R [52][0] <= 8'b0111_1111;					inform_R [53][0] <= 8'b0111_1111;					inform_R [54][0] <= 8'b0111_1111;					inform_R [55][0] <= 8'b0111_1111;					inform_R [56][0] <= 8'b0111_1111;					inform_R [57][0] <= 8'b0111_1111;					inform_R [58][0] <= 8'b0111_1111;					inform_R [59][0] <= 8'b0000_0000;					inform_R [60][0] <= 8'b0111_1111;					inform_R [61][0] <= 8'b0000_0000;					inform_R [62][0] <= 8'b0000_0000;					inform_R [63][0] <= 8'b0000_0000;					inform_R [64][0] <= 8'b0111_1111;					inform_R [65][0] <= 8'b0111_1111;					inform_R [66][0] <= 8'b0111_1111;					inform_R [67][0] <= 8'b0111_1111;					inform_R [68][0] <= 8'b0111_1111;					inform_R [69][0] <= 8'b0111_1111;					inform_R [70][0] <= 8'b0111_1111;					inform_R [71][0] <= 8'b0111_1111;					inform_R [72][0] <= 8'b0111_1111;					inform_R [73][0] <= 8'b0111_1111;					inform_R [74][0] <= 8'b0111_1111;					inform_R [75][0] <= 8'b0111_1111;					inform_R [76][0] <= 8'b0111_1111;					inform_R [77][0] <= 8'b0111_1111;					inform_R [78][0] <= 8'b0111_1111;					inform_R [79][0] <= 8'b0111_1111;					inform_R [80][0] <= 8'b0111_1111;					inform_R [81][0] <= 8'b0111_1111;					inform_R [82][0] <= 8'b0111_1111;					inform_R [83][0] <= 8'b0111_1111;					inform_R [84][0] <= 8'b0111_1111;					inform_R [85][0] <= 8'b0111_1111;					inform_R [86][0] <= 8'b0111_1111;					inform_R [87][0] <= 8'b0000_0000;					inform_R [88][0] <= 8'b0111_1111;					inform_R [89][0] <= 8'b0111_1111;					inform_R [90][0] <= 8'b0111_1111;					inform_R [91][0] <= 8'b0000_0000;					inform_R [92][0] <= 8'b0111_1111;					inform_R [93][0] <= 8'b0000_0000;					inform_R [94][0] <= 8'b0000_0000;					inform_R [95][0] <= 8'b0000_0000;					inform_R [96][0] <= 8'b0111_1111;					inform_R [97][0] <= 8'b0111_1111;					inform_R [98][0] <= 8'b0111_1111;					inform_R [99][0] <= 8'b0111_1111;					inform_R [100][0] <= 8'b0111_1111;					inform_R [101][0] <= 8'b0111_1111;					inform_R [102][0] <= 8'b0111_1111;					inform_R [103][0] <= 8'b0000_0000;					inform_R [104][0] <= 8'b0111_1111;					inform_R [105][0] <= 8'b0111_1111;					inform_R [106][0] <= 8'b0000_0000;					inform_R [107][0] <= 8'b0000_0000;					inform_R [108][0] <= 8'b0000_0000;					inform_R [109][0] <= 8'b0000_0000;					inform_R [110][0] <= 8'b0000_0000;					inform_R [111][0] <= 8'b0000_0000;					inform_R [112][0] <= 8'b0111_1111;					inform_R [113][0] <= 8'b0000_0000;					inform_R [114][0] <= 8'b0000_0000;					inform_R [115][0] <= 8'b0000_0000;					inform_R [116][0] <= 8'b0000_0000;					inform_R [117][0] <= 8'b0000_0000;					inform_R [118][0] <= 8'b0000_0000;					inform_R [119][0] <= 8'b0000_0000;					inform_R [120][0] <= 8'b0000_0000;					inform_R [121][0] <= 8'b0000_0000;					inform_R [122][0] <= 8'b0000_0000;					inform_R [123][0] <= 8'b0000_0000;					inform_R [124][0] <= 8'b0000_0000;					inform_R [125][0] <= 8'b0000_0000;					inform_R [126][0] <= 8'b0000_0000;					inform_R [127][0] <= 8'b0000_0000;					inform_R [128][0] <= 8'b0111_1111;					inform_R [129][0] <= 8'b0111_1111;					inform_R [130][0] <= 8'b0111_1111;					inform_R [131][0] <= 8'b0111_1111;					inform_R [132][0] <= 8'b0111_1111;					inform_R [133][0] <= 8'b0111_1111;					inform_R [134][0] <= 8'b0111_1111;					inform_R [135][0] <= 8'b0111_1111;					inform_R [136][0] <= 8'b0111_1111;					inform_R [137][0] <= 8'b0111_1111;					inform_R [138][0] <= 8'b0111_1111;					inform_R [139][0] <= 8'b0111_1111;					inform_R [140][0] <= 8'b0111_1111;					inform_R [141][0] <= 8'b0111_1111;					inform_R [142][0] <= 8'b0111_1111;					inform_R [143][0] <= 8'b0000_0000;					inform_R [144][0] <= 8'b0111_1111;					inform_R [145][0] <= 8'b0111_1111;					inform_R [146][0] <= 8'b0111_1111;					inform_R [147][0] <= 8'b0111_1111;					inform_R [148][0] <= 8'b0111_1111;					inform_R [149][0] <= 8'b0111_1111;					inform_R [150][0] <= 8'b0000_0000;					inform_R [151][0] <= 8'b0000_0000;					inform_R [152][0] <= 8'b0111_1111;					inform_R [153][0] <= 8'b0000_0000;					inform_R [154][0] <= 8'b0000_0000;					inform_R [155][0] <= 8'b0000_0000;					inform_R [156][0] <= 8'b0000_0000;					inform_R [157][0] <= 8'b0000_0000;					inform_R [158][0] <= 8'b0000_0000;					inform_R [159][0] <= 8'b0000_0000;					inform_R [160][0] <= 8'b0111_1111;					inform_R [161][0] <= 8'b0111_1111;					inform_R [162][0] <= 8'b0111_1111;					inform_R [163][0] <= 8'b0000_0000;					inform_R [164][0] <= 8'b0111_1111;					inform_R [165][0] <= 8'b0000_0000;					inform_R [166][0] <= 8'b0000_0000;					inform_R [167][0] <= 8'b0000_0000;					inform_R [168][0] <= 8'b0111_1111;					inform_R [169][0] <= 8'b0000_0000;					inform_R [170][0] <= 8'b0000_0000;					inform_R [171][0] <= 8'b0000_0000;					inform_R [172][0] <= 8'b0000_0000;					inform_R [173][0] <= 8'b0000_0000;					inform_R [174][0] <= 8'b0000_0000;					inform_R [175][0] <= 8'b0000_0000;					inform_R [176][0] <= 8'b0000_0000;					inform_R [177][0] <= 8'b0000_0000;					inform_R [178][0] <= 8'b0000_0000;					inform_R [179][0] <= 8'b0000_0000;					inform_R [180][0] <= 8'b0000_0000;					inform_R [181][0] <= 8'b0000_0000;					inform_R [182][0] <= 8'b0000_0000;					inform_R [183][0] <= 8'b0000_0000;					inform_R [184][0] <= 8'b0000_0000;					inform_R [185][0] <= 8'b0000_0000;					inform_R [186][0] <= 8'b0000_0000;					inform_R [187][0] <= 8'b0000_0000;					inform_R [188][0] <= 8'b0000_0000;					inform_R [189][0] <= 8'b0000_0000;					inform_R [190][0] <= 8'b0000_0000;					inform_R [191][0] <= 8'b0000_0000;					inform_R [192][0] <= 8'b0111_1111;					inform_R [193][0] <= 8'b0111_1111;					inform_R [194][0] <= 8'b0111_1111;					inform_R [195][0] <= 8'b0000_0000;					inform_R [196][0] <= 8'b0111_1111;					inform_R [197][0] <= 8'b0000_0000;					inform_R [198][0] <= 8'b0000_0000;					inform_R [199][0] <= 8'b0000_0000;					inform_R [200][0] <= 8'b0000_0000;					inform_R [201][0] <= 8'b0000_0000;					inform_R [202][0] <= 8'b0000_0000;					inform_R [203][0] <= 8'b0000_0000;					inform_R [204][0] <= 8'b0000_0000;					inform_R [205][0] <= 8'b0000_0000;					inform_R [206][0] <= 8'b0000_0000;					inform_R [207][0] <= 8'b0000_0000;					inform_R [208][0] <= 8'b0000_0000;					inform_R [209][0] <= 8'b0000_0000;					inform_R [210][0] <= 8'b0000_0000;					inform_R [211][0] <= 8'b0000_0000;					inform_R [212][0] <= 8'b0000_0000;					inform_R [213][0] <= 8'b0000_0000;					inform_R [214][0] <= 8'b0000_0000;					inform_R [215][0] <= 8'b0000_0000;					inform_R [216][0] <= 8'b0000_0000;					inform_R [217][0] <= 8'b0000_0000;					inform_R [218][0] <= 8'b0000_0000;					inform_R [219][0] <= 8'b0000_0000;					inform_R [220][0] <= 8'b0000_0000;					inform_R [221][0] <= 8'b0000_0000;					inform_R [222][0] <= 8'b0000_0000;					inform_R [223][0] <= 8'b0000_0000;					inform_R [224][0] <= 8'b0000_0000;					inform_R [225][0] <= 8'b0000_0000;					inform_R [226][0] <= 8'b0000_0000;					inform_R [227][0] <= 8'b0000_0000;					inform_R [228][0] <= 8'b0000_0000;					inform_R [229][0] <= 8'b0000_0000;					inform_R [230][0] <= 8'b0000_0000;					inform_R [231][0] <= 8'b0000_0000;					inform_R [232][0] <= 8'b0000_0000;					inform_R [233][0] <= 8'b0000_0000;					inform_R [234][0] <= 8'b0000_0000;					inform_R [235][0] <= 8'b0000_0000;					inform_R [236][0] <= 8'b0000_0000;					inform_R [237][0] <= 8'b0000_0000;					inform_R [238][0] <= 8'b0000_0000;					inform_R [239][0] <= 8'b0000_0000;					inform_R [240][0] <= 8'b0000_0000;					inform_R [241][0] <= 8'b0000_0000;					inform_R [242][0] <= 8'b0000_0000;					inform_R [243][0] <= 8'b0000_0000;					inform_R [244][0] <= 8'b0000_0000;					inform_R [245][0] <= 8'b0000_0000;					inform_R [246][0] <= 8'b0000_0000;					inform_R [247][0] <= 8'b0000_0000;					inform_R [248][0] <= 8'b0000_0000;					inform_R [249][0] <= 8'b0000_0000;					inform_R [250][0] <= 8'b0000_0000;					inform_R [251][0] <= 8'b0000_0000;					inform_R [252][0] <= 8'b0000_0000;					inform_R [253][0] <= 8'b0000_0000;					inform_R [254][0] <= 8'b0000_0000;					inform_R [255][0] <= 8'b0000_0000;					inform_L [0][8] <= LLR_1;					inform_L [1][8] <= LLR_2;					inform_L [2][8] <= LLR_3;					inform_L [3][8] <= LLR_4;					inform_L [4][8] <= LLR_5;					inform_L [5][8] <= LLR_6;					inform_L [6][8] <= LLR_7;					inform_L [7][8] <= LLR_8;					inform_L [8][8] <= LLR_9;					inform_L [9][8] <= LLR_10;					inform_L [10][8] <= LLR_11;					inform_L [11][8] <= LLR_12;					inform_L [12][8] <= LLR_13;					inform_L [13][8] <= LLR_14;					inform_L [14][8] <= LLR_15;					inform_L [15][8] <= LLR_16;					inform_L [16][8] <= LLR_17;					inform_L [17][8] <= LLR_18;					inform_L [18][8] <= LLR_19;					inform_L [19][8] <= LLR_20;					inform_L [20][8] <= LLR_21;					inform_L [21][8] <= LLR_22;					inform_L [22][8] <= LLR_23;					inform_L [23][8] <= LLR_24;					inform_L [24][8] <= LLR_25;					inform_L [25][8] <= LLR_26;					inform_L [26][8] <= LLR_27;					inform_L [27][8] <= LLR_28;					inform_L [28][8] <= LLR_29;					inform_L [29][8] <= LLR_30;					inform_L [30][8] <= LLR_31;					inform_L [31][8] <= LLR_32;					inform_L [32][8] <= LLR_33;					inform_L [33][8] <= LLR_34;					inform_L [34][8] <= LLR_35;					inform_L [35][8] <= LLR_36;					inform_L [36][8] <= LLR_37;					inform_L [37][8] <= LLR_38;					inform_L [38][8] <= LLR_39;					inform_L [39][8] <= LLR_40;					inform_L [40][8] <= LLR_41;					inform_L [41][8] <= LLR_42;					inform_L [42][8] <= LLR_43;					inform_L [43][8] <= LLR_44;					inform_L [44][8] <= LLR_45;					inform_L [45][8] <= LLR_46;					inform_L [46][8] <= LLR_47;					inform_L [47][8] <= LLR_48;					inform_L [48][8] <= LLR_49;					inform_L [49][8] <= LLR_50;					inform_L [50][8] <= LLR_51;					inform_L [51][8] <= LLR_52;					inform_L [52][8] <= LLR_53;					inform_L [53][8] <= LLR_54;					inform_L [54][8] <= LLR_55;					inform_L [55][8] <= LLR_56;					inform_L [56][8] <= LLR_57;					inform_L [57][8] <= LLR_58;					inform_L [58][8] <= LLR_59;					inform_L [59][8] <= LLR_60;					inform_L [60][8] <= LLR_61;					inform_L [61][8] <= LLR_62;					inform_L [62][8] <= LLR_63;					inform_L [63][8] <= LLR_64;					inform_L [64][8] <= LLR_65;					inform_L [65][8] <= LLR_66;					inform_L [66][8] <= LLR_67;					inform_L [67][8] <= LLR_68;					inform_L [68][8] <= LLR_69;					inform_L [69][8] <= LLR_70;					inform_L [70][8] <= LLR_71;					inform_L [71][8] <= LLR_72;					inform_L [72][8] <= LLR_73;					inform_L [73][8] <= LLR_74;					inform_L [74][8] <= LLR_75;					inform_L [75][8] <= LLR_76;					inform_L [76][8] <= LLR_77;					inform_L [77][8] <= LLR_78;					inform_L [78][8] <= LLR_79;					inform_L [79][8] <= LLR_80;					inform_L [80][8] <= LLR_81;					inform_L [81][8] <= LLR_82;					inform_L [82][8] <= LLR_83;					inform_L [83][8] <= LLR_84;					inform_L [84][8] <= LLR_85;					inform_L [85][8] <= LLR_86;					inform_L [86][8] <= LLR_87;					inform_L [87][8] <= LLR_88;					inform_L [88][8] <= LLR_89;					inform_L [89][8] <= LLR_90;					inform_L [90][8] <= LLR_91;					inform_L [91][8] <= LLR_92;					inform_L [92][8] <= LLR_93;					inform_L [93][8] <= LLR_94;					inform_L [94][8] <= LLR_95;					inform_L [95][8] <= LLR_96;					inform_L [96][8] <= LLR_97;					inform_L [97][8] <= LLR_98;					inform_L [98][8] <= LLR_99;					inform_L [99][8] <= LLR_100;					inform_L [100][8] <= LLR_101;					inform_L [101][8] <= LLR_102;					inform_L [102][8] <= LLR_103;					inform_L [103][8] <= LLR_104;					inform_L [104][8] <= LLR_105;					inform_L [105][8] <= LLR_106;					inform_L [106][8] <= LLR_107;					inform_L [107][8] <= LLR_108;					inform_L [108][8] <= LLR_109;					inform_L [109][8] <= LLR_110;					inform_L [110][8] <= LLR_111;					inform_L [111][8] <= LLR_112;					inform_L [112][8] <= LLR_113;					inform_L [113][8] <= LLR_114;					inform_L [114][8] <= LLR_115;					inform_L [115][8] <= LLR_116;					inform_L [116][8] <= LLR_117;					inform_L [117][8] <= LLR_118;					inform_L [118][8] <= LLR_119;					inform_L [119][8] <= LLR_120;					inform_L [120][8] <= LLR_121;					inform_L [121][8] <= LLR_122;					inform_L [122][8] <= LLR_123;					inform_L [123][8] <= LLR_124;					inform_L [124][8] <= LLR_125;					inform_L [125][8] <= LLR_126;					inform_L [126][8] <= LLR_127;					inform_L [127][8] <= LLR_128;					inform_L [128][8] <= LLR_129;					inform_L [129][8] <= LLR_130;					inform_L [130][8] <= LLR_131;					inform_L [131][8] <= LLR_132;					inform_L [132][8] <= LLR_133;					inform_L [133][8] <= LLR_134;					inform_L [134][8] <= LLR_135;					inform_L [135][8] <= LLR_136;					inform_L [136][8] <= LLR_137;					inform_L [137][8] <= LLR_138;					inform_L [138][8] <= LLR_139;					inform_L [139][8] <= LLR_140;					inform_L [140][8] <= LLR_141;					inform_L [141][8] <= LLR_142;					inform_L [142][8] <= LLR_143;					inform_L [143][8] <= LLR_144;					inform_L [144][8] <= LLR_145;					inform_L [145][8] <= LLR_146;					inform_L [146][8] <= LLR_147;					inform_L [147][8] <= LLR_148;					inform_L [148][8] <= LLR_149;					inform_L [149][8] <= LLR_150;					inform_L [150][8] <= LLR_151;					inform_L [151][8] <= LLR_152;					inform_L [152][8] <= LLR_153;					inform_L [153][8] <= LLR_154;					inform_L [154][8] <= LLR_155;					inform_L [155][8] <= LLR_156;					inform_L [156][8] <= LLR_157;					inform_L [157][8] <= LLR_158;					inform_L [158][8] <= LLR_159;					inform_L [159][8] <= LLR_160;					inform_L [160][8] <= LLR_161;					inform_L [161][8] <= LLR_162;					inform_L [162][8] <= LLR_163;					inform_L [163][8] <= LLR_164;					inform_L [164][8] <= LLR_165;					inform_L [165][8] <= LLR_166;					inform_L [166][8] <= LLR_167;					inform_L [167][8] <= LLR_168;					inform_L [168][8] <= LLR_169;					inform_L [169][8] <= LLR_170;					inform_L [170][8] <= LLR_171;					inform_L [171][8] <= LLR_172;					inform_L [172][8] <= LLR_173;					inform_L [173][8] <= LLR_174;					inform_L [174][8] <= LLR_175;					inform_L [175][8] <= LLR_176;					inform_L [176][8] <= LLR_177;					inform_L [177][8] <= LLR_178;					inform_L [178][8] <= LLR_179;					inform_L [179][8] <= LLR_180;					inform_L [180][8] <= LLR_181;					inform_L [181][8] <= LLR_182;					inform_L [182][8] <= LLR_183;					inform_L [183][8] <= LLR_184;					inform_L [184][8] <= LLR_185;					inform_L [185][8] <= LLR_186;					inform_L [186][8] <= LLR_187;					inform_L [187][8] <= LLR_188;					inform_L [188][8] <= LLR_189;					inform_L [189][8] <= LLR_190;					inform_L [190][8] <= LLR_191;					inform_L [191][8] <= LLR_192;					inform_L [192][8] <= LLR_193;					inform_L [193][8] <= LLR_194;					inform_L [194][8] <= LLR_195;					inform_L [195][8] <= LLR_196;					inform_L [196][8] <= LLR_197;					inform_L [197][8] <= LLR_198;					inform_L [198][8] <= LLR_199;					inform_L [199][8] <= LLR_200;					inform_L [200][8] <= LLR_201;					inform_L [201][8] <= LLR_202;					inform_L [202][8] <= LLR_203;					inform_L [203][8] <= LLR_204;					inform_L [204][8] <= LLR_205;					inform_L [205][8] <= LLR_206;					inform_L [206][8] <= LLR_207;					inform_L [207][8] <= LLR_208;					inform_L [208][8] <= LLR_209;					inform_L [209][8] <= LLR_210;					inform_L [210][8] <= LLR_211;					inform_L [211][8] <= LLR_212;					inform_L [212][8] <= LLR_213;					inform_L [213][8] <= LLR_214;					inform_L [214][8] <= LLR_215;					inform_L [215][8] <= LLR_216;					inform_L [216][8] <= LLR_217;					inform_L [217][8] <= LLR_218;					inform_L [218][8] <= LLR_219;					inform_L [219][8] <= LLR_220;					inform_L [220][8] <= LLR_221;					inform_L [221][8] <= LLR_222;					inform_L [222][8] <= LLR_223;					inform_L [223][8] <= LLR_224;					inform_L [224][8] <= LLR_225;					inform_L [225][8] <= LLR_226;					inform_L [226][8] <= LLR_227;					inform_L [227][8] <= LLR_228;					inform_L [228][8] <= LLR_229;					inform_L [229][8] <= LLR_230;					inform_L [230][8] <= LLR_231;					inform_L [231][8] <= LLR_232;					inform_L [232][8] <= LLR_233;					inform_L [233][8] <= LLR_234;					inform_L [234][8] <= LLR_235;					inform_L [235][8] <= LLR_236;					inform_L [236][8] <= LLR_237;					inform_L [237][8] <= LLR_238;					inform_L [238][8] <= LLR_239;					inform_L [239][8] <= LLR_240;					inform_L [240][8] <= LLR_241;					inform_L [241][8] <= LLR_242;					inform_L [242][8] <= LLR_243;					inform_L [243][8] <= LLR_244;					inform_L [244][8] <= LLR_245;					inform_L [245][8] <= LLR_246;					inform_L [246][8] <= LLR_247;					inform_L [247][8] <= LLR_248;					inform_L [248][8] <= LLR_249;					inform_L [249][8] <= LLR_250;					inform_L [250][8] <= LLR_251;					inform_L [251][8] <= LLR_252;					inform_L [252][8] <= LLR_253;					inform_L [253][8] <= LLR_254;					inform_L [254][8] <= LLR_255;					inform_L [255][8] <= LLR_256;				end				for (x = 0; x < 256; x = x + 1)					for (y = 0; y < 8; y = y + 1)					begin						inform_R[x][y+1] <= 8'd0;						inform_L[x][y] <= 8'd0;					end			end
			BUSY_LEFT:			begin				if(clk_counter == 2'b11)begin					case (w2r)						1:						begin							inform_R[0][1] = r_cell_wire[0];							inform_R[1][1] = r_cell_wire[1];							inform_R[2][1] = r_cell_wire[2];							inform_R[3][1] = r_cell_wire[3];							inform_R[4][1] = r_cell_wire[4];							inform_R[5][1] = r_cell_wire[5];							inform_R[6][1] = r_cell_wire[6];							inform_R[7][1] = r_cell_wire[7];							inform_R[8][1] = r_cell_wire[8];							inform_R[9][1] = r_cell_wire[9];							inform_R[10][1] = r_cell_wire[10];							inform_R[11][1] = r_cell_wire[11];							inform_R[12][1] = r_cell_wire[12];							inform_R[13][1] = r_cell_wire[13];							inform_R[14][1] = r_cell_wire[14];							inform_R[15][1] = r_cell_wire[15];							inform_R[16][1] = r_cell_wire[16];							inform_R[17][1] = r_cell_wire[17];							inform_R[18][1] = r_cell_wire[18];							inform_R[19][1] = r_cell_wire[19];							inform_R[20][1] = r_cell_wire[20];							inform_R[21][1] = r_cell_wire[21];							inform_R[22][1] = r_cell_wire[22];							inform_R[23][1] = r_cell_wire[23];							inform_R[24][1] = r_cell_wire[24];							inform_R[25][1] = r_cell_wire[25];							inform_R[26][1] = r_cell_wire[26];							inform_R[27][1] = r_cell_wire[27];							inform_R[28][1] = r_cell_wire[28];							inform_R[29][1] = r_cell_wire[29];							inform_R[30][1] = r_cell_wire[30];							inform_R[31][1] = r_cell_wire[31];							inform_R[32][1] = r_cell_wire[32];							inform_R[33][1] = r_cell_wire[33];							inform_R[34][1] = r_cell_wire[34];							inform_R[35][1] = r_cell_wire[35];							inform_R[36][1] = r_cell_wire[36];							inform_R[37][1] = r_cell_wire[37];							inform_R[38][1] = r_cell_wire[38];							inform_R[39][1] = r_cell_wire[39];							inform_R[40][1] = r_cell_wire[40];							inform_R[41][1] = r_cell_wire[41];							inform_R[42][1] = r_cell_wire[42];							inform_R[43][1] = r_cell_wire[43];							inform_R[44][1] = r_cell_wire[44];							inform_R[45][1] = r_cell_wire[45];							inform_R[46][1] = r_cell_wire[46];							inform_R[47][1] = r_cell_wire[47];							inform_R[48][1] = r_cell_wire[48];							inform_R[49][1] = r_cell_wire[49];							inform_R[50][1] = r_cell_wire[50];							inform_R[51][1] = r_cell_wire[51];							inform_R[52][1] = r_cell_wire[52];							inform_R[53][1] = r_cell_wire[53];							inform_R[54][1] = r_cell_wire[54];							inform_R[55][1] = r_cell_wire[55];							inform_R[56][1] = r_cell_wire[56];							inform_R[57][1] = r_cell_wire[57];							inform_R[58][1] = r_cell_wire[58];							inform_R[59][1] = r_cell_wire[59];							inform_R[60][1] = r_cell_wire[60];							inform_R[61][1] = r_cell_wire[61];							inform_R[62][1] = r_cell_wire[62];							inform_R[63][1] = r_cell_wire[63];							inform_R[64][1] = r_cell_wire[64];							inform_R[65][1] = r_cell_wire[65];							inform_R[66][1] = r_cell_wire[66];							inform_R[67][1] = r_cell_wire[67];							inform_R[68][1] = r_cell_wire[68];							inform_R[69][1] = r_cell_wire[69];							inform_R[70][1] = r_cell_wire[70];							inform_R[71][1] = r_cell_wire[71];							inform_R[72][1] = r_cell_wire[72];							inform_R[73][1] = r_cell_wire[73];							inform_R[74][1] = r_cell_wire[74];							inform_R[75][1] = r_cell_wire[75];							inform_R[76][1] = r_cell_wire[76];							inform_R[77][1] = r_cell_wire[77];							inform_R[78][1] = r_cell_wire[78];							inform_R[79][1] = r_cell_wire[79];							inform_R[80][1] = r_cell_wire[80];							inform_R[81][1] = r_cell_wire[81];							inform_R[82][1] = r_cell_wire[82];							inform_R[83][1] = r_cell_wire[83];							inform_R[84][1] = r_cell_wire[84];							inform_R[85][1] = r_cell_wire[85];							inform_R[86][1] = r_cell_wire[86];							inform_R[87][1] = r_cell_wire[87];							inform_R[88][1] = r_cell_wire[88];							inform_R[89][1] = r_cell_wire[89];							inform_R[90][1] = r_cell_wire[90];							inform_R[91][1] = r_cell_wire[91];							inform_R[92][1] = r_cell_wire[92];							inform_R[93][1] = r_cell_wire[93];							inform_R[94][1] = r_cell_wire[94];							inform_R[95][1] = r_cell_wire[95];							inform_R[96][1] = r_cell_wire[96];							inform_R[97][1] = r_cell_wire[97];							inform_R[98][1] = r_cell_wire[98];							inform_R[99][1] = r_cell_wire[99];							inform_R[100][1] = r_cell_wire[100];							inform_R[101][1] = r_cell_wire[101];							inform_R[102][1] = r_cell_wire[102];							inform_R[103][1] = r_cell_wire[103];							inform_R[104][1] = r_cell_wire[104];							inform_R[105][1] = r_cell_wire[105];							inform_R[106][1] = r_cell_wire[106];							inform_R[107][1] = r_cell_wire[107];							inform_R[108][1] = r_cell_wire[108];							inform_R[109][1] = r_cell_wire[109];							inform_R[110][1] = r_cell_wire[110];							inform_R[111][1] = r_cell_wire[111];							inform_R[112][1] = r_cell_wire[112];							inform_R[113][1] = r_cell_wire[113];							inform_R[114][1] = r_cell_wire[114];							inform_R[115][1] = r_cell_wire[115];							inform_R[116][1] = r_cell_wire[116];							inform_R[117][1] = r_cell_wire[117];							inform_R[118][1] = r_cell_wire[118];							inform_R[119][1] = r_cell_wire[119];							inform_R[120][1] = r_cell_wire[120];							inform_R[121][1] = r_cell_wire[121];							inform_R[122][1] = r_cell_wire[122];							inform_R[123][1] = r_cell_wire[123];							inform_R[124][1] = r_cell_wire[124];							inform_R[125][1] = r_cell_wire[125];							inform_R[126][1] = r_cell_wire[126];							inform_R[127][1] = r_cell_wire[127];							inform_R[128][1] = r_cell_wire[128];							inform_R[129][1] = r_cell_wire[129];							inform_R[130][1] = r_cell_wire[130];							inform_R[131][1] = r_cell_wire[131];							inform_R[132][1] = r_cell_wire[132];							inform_R[133][1] = r_cell_wire[133];							inform_R[134][1] = r_cell_wire[134];							inform_R[135][1] = r_cell_wire[135];							inform_R[136][1] = r_cell_wire[136];							inform_R[137][1] = r_cell_wire[137];							inform_R[138][1] = r_cell_wire[138];							inform_R[139][1] = r_cell_wire[139];							inform_R[140][1] = r_cell_wire[140];							inform_R[141][1] = r_cell_wire[141];							inform_R[142][1] = r_cell_wire[142];							inform_R[143][1] = r_cell_wire[143];							inform_R[144][1] = r_cell_wire[144];							inform_R[145][1] = r_cell_wire[145];							inform_R[146][1] = r_cell_wire[146];							inform_R[147][1] = r_cell_wire[147];							inform_R[148][1] = r_cell_wire[148];							inform_R[149][1] = r_cell_wire[149];							inform_R[150][1] = r_cell_wire[150];							inform_R[151][1] = r_cell_wire[151];							inform_R[152][1] = r_cell_wire[152];							inform_R[153][1] = r_cell_wire[153];							inform_R[154][1] = r_cell_wire[154];							inform_R[155][1] = r_cell_wire[155];							inform_R[156][1] = r_cell_wire[156];							inform_R[157][1] = r_cell_wire[157];							inform_R[158][1] = r_cell_wire[158];							inform_R[159][1] = r_cell_wire[159];							inform_R[160][1] = r_cell_wire[160];							inform_R[161][1] = r_cell_wire[161];							inform_R[162][1] = r_cell_wire[162];							inform_R[163][1] = r_cell_wire[163];							inform_R[164][1] = r_cell_wire[164];							inform_R[165][1] = r_cell_wire[165];							inform_R[166][1] = r_cell_wire[166];							inform_R[167][1] = r_cell_wire[167];							inform_R[168][1] = r_cell_wire[168];							inform_R[169][1] = r_cell_wire[169];							inform_R[170][1] = r_cell_wire[170];							inform_R[171][1] = r_cell_wire[171];							inform_R[172][1] = r_cell_wire[172];							inform_R[173][1] = r_cell_wire[173];							inform_R[174][1] = r_cell_wire[174];							inform_R[175][1] = r_cell_wire[175];							inform_R[176][1] = r_cell_wire[176];							inform_R[177][1] = r_cell_wire[177];							inform_R[178][1] = r_cell_wire[178];							inform_R[179][1] = r_cell_wire[179];							inform_R[180][1] = r_cell_wire[180];							inform_R[181][1] = r_cell_wire[181];							inform_R[182][1] = r_cell_wire[182];							inform_R[183][1] = r_cell_wire[183];							inform_R[184][1] = r_cell_wire[184];							inform_R[185][1] = r_cell_wire[185];							inform_R[186][1] = r_cell_wire[186];							inform_R[187][1] = r_cell_wire[187];							inform_R[188][1] = r_cell_wire[188];							inform_R[189][1] = r_cell_wire[189];							inform_R[190][1] = r_cell_wire[190];							inform_R[191][1] = r_cell_wire[191];							inform_R[192][1] = r_cell_wire[192];							inform_R[193][1] = r_cell_wire[193];							inform_R[194][1] = r_cell_wire[194];							inform_R[195][1] = r_cell_wire[195];							inform_R[196][1] = r_cell_wire[196];							inform_R[197][1] = r_cell_wire[197];							inform_R[198][1] = r_cell_wire[198];							inform_R[199][1] = r_cell_wire[199];							inform_R[200][1] = r_cell_wire[200];							inform_R[201][1] = r_cell_wire[201];							inform_R[202][1] = r_cell_wire[202];							inform_R[203][1] = r_cell_wire[203];							inform_R[204][1] = r_cell_wire[204];							inform_R[205][1] = r_cell_wire[205];							inform_R[206][1] = r_cell_wire[206];							inform_R[207][1] = r_cell_wire[207];							inform_R[208][1] = r_cell_wire[208];							inform_R[209][1] = r_cell_wire[209];							inform_R[210][1] = r_cell_wire[210];							inform_R[211][1] = r_cell_wire[211];							inform_R[212][1] = r_cell_wire[212];							inform_R[213][1] = r_cell_wire[213];							inform_R[214][1] = r_cell_wire[214];							inform_R[215][1] = r_cell_wire[215];							inform_R[216][1] = r_cell_wire[216];							inform_R[217][1] = r_cell_wire[217];							inform_R[218][1] = r_cell_wire[218];							inform_R[219][1] = r_cell_wire[219];							inform_R[220][1] = r_cell_wire[220];							inform_R[221][1] = r_cell_wire[221];							inform_R[222][1] = r_cell_wire[222];							inform_R[223][1] = r_cell_wire[223];							inform_R[224][1] = r_cell_wire[224];							inform_R[225][1] = r_cell_wire[225];							inform_R[226][1] = r_cell_wire[226];							inform_R[227][1] = r_cell_wire[227];							inform_R[228][1] = r_cell_wire[228];							inform_R[229][1] = r_cell_wire[229];							inform_R[230][1] = r_cell_wire[230];							inform_R[231][1] = r_cell_wire[231];							inform_R[232][1] = r_cell_wire[232];							inform_R[233][1] = r_cell_wire[233];							inform_R[234][1] = r_cell_wire[234];							inform_R[235][1] = r_cell_wire[235];							inform_R[236][1] = r_cell_wire[236];							inform_R[237][1] = r_cell_wire[237];							inform_R[238][1] = r_cell_wire[238];							inform_R[239][1] = r_cell_wire[239];							inform_R[240][1] = r_cell_wire[240];							inform_R[241][1] = r_cell_wire[241];							inform_R[242][1] = r_cell_wire[242];							inform_R[243][1] = r_cell_wire[243];							inform_R[244][1] = r_cell_wire[244];							inform_R[245][1] = r_cell_wire[245];							inform_R[246][1] = r_cell_wire[246];							inform_R[247][1] = r_cell_wire[247];							inform_R[248][1] = r_cell_wire[248];							inform_R[249][1] = r_cell_wire[249];							inform_R[250][1] = r_cell_wire[250];							inform_R[251][1] = r_cell_wire[251];							inform_R[252][1] = r_cell_wire[252];							inform_R[253][1] = r_cell_wire[253];							inform_R[254][1] = r_cell_wire[254];							inform_R[255][1] = r_cell_wire[255];							inform_L[0][0] = l_cell_wire[0];							inform_L[1][0] = l_cell_wire[1];							inform_L[2][0] = l_cell_wire[2];							inform_L[3][0] = l_cell_wire[3];							inform_L[4][0] = l_cell_wire[4];							inform_L[5][0] = l_cell_wire[5];							inform_L[6][0] = l_cell_wire[6];							inform_L[7][0] = l_cell_wire[7];							inform_L[8][0] = l_cell_wire[8];							inform_L[9][0] = l_cell_wire[9];							inform_L[10][0] = l_cell_wire[10];							inform_L[11][0] = l_cell_wire[11];							inform_L[12][0] = l_cell_wire[12];							inform_L[13][0] = l_cell_wire[13];							inform_L[14][0] = l_cell_wire[14];							inform_L[15][0] = l_cell_wire[15];							inform_L[16][0] = l_cell_wire[16];							inform_L[17][0] = l_cell_wire[17];							inform_L[18][0] = l_cell_wire[18];							inform_L[19][0] = l_cell_wire[19];							inform_L[20][0] = l_cell_wire[20];							inform_L[21][0] = l_cell_wire[21];							inform_L[22][0] = l_cell_wire[22];							inform_L[23][0] = l_cell_wire[23];							inform_L[24][0] = l_cell_wire[24];							inform_L[25][0] = l_cell_wire[25];							inform_L[26][0] = l_cell_wire[26];							inform_L[27][0] = l_cell_wire[27];							inform_L[28][0] = l_cell_wire[28];							inform_L[29][0] = l_cell_wire[29];							inform_L[30][0] = l_cell_wire[30];							inform_L[31][0] = l_cell_wire[31];							inform_L[32][0] = l_cell_wire[32];							inform_L[33][0] = l_cell_wire[33];							inform_L[34][0] = l_cell_wire[34];							inform_L[35][0] = l_cell_wire[35];							inform_L[36][0] = l_cell_wire[36];							inform_L[37][0] = l_cell_wire[37];							inform_L[38][0] = l_cell_wire[38];							inform_L[39][0] = l_cell_wire[39];							inform_L[40][0] = l_cell_wire[40];							inform_L[41][0] = l_cell_wire[41];							inform_L[42][0] = l_cell_wire[42];							inform_L[43][0] = l_cell_wire[43];							inform_L[44][0] = l_cell_wire[44];							inform_L[45][0] = l_cell_wire[45];							inform_L[46][0] = l_cell_wire[46];							inform_L[47][0] = l_cell_wire[47];							inform_L[48][0] = l_cell_wire[48];							inform_L[49][0] = l_cell_wire[49];							inform_L[50][0] = l_cell_wire[50];							inform_L[51][0] = l_cell_wire[51];							inform_L[52][0] = l_cell_wire[52];							inform_L[53][0] = l_cell_wire[53];							inform_L[54][0] = l_cell_wire[54];							inform_L[55][0] = l_cell_wire[55];							inform_L[56][0] = l_cell_wire[56];							inform_L[57][0] = l_cell_wire[57];							inform_L[58][0] = l_cell_wire[58];							inform_L[59][0] = l_cell_wire[59];							inform_L[60][0] = l_cell_wire[60];							inform_L[61][0] = l_cell_wire[61];							inform_L[62][0] = l_cell_wire[62];							inform_L[63][0] = l_cell_wire[63];							inform_L[64][0] = l_cell_wire[64];							inform_L[65][0] = l_cell_wire[65];							inform_L[66][0] = l_cell_wire[66];							inform_L[67][0] = l_cell_wire[67];							inform_L[68][0] = l_cell_wire[68];							inform_L[69][0] = l_cell_wire[69];							inform_L[70][0] = l_cell_wire[70];							inform_L[71][0] = l_cell_wire[71];							inform_L[72][0] = l_cell_wire[72];							inform_L[73][0] = l_cell_wire[73];							inform_L[74][0] = l_cell_wire[74];							inform_L[75][0] = l_cell_wire[75];							inform_L[76][0] = l_cell_wire[76];							inform_L[77][0] = l_cell_wire[77];							inform_L[78][0] = l_cell_wire[78];							inform_L[79][0] = l_cell_wire[79];							inform_L[80][0] = l_cell_wire[80];							inform_L[81][0] = l_cell_wire[81];							inform_L[82][0] = l_cell_wire[82];							inform_L[83][0] = l_cell_wire[83];							inform_L[84][0] = l_cell_wire[84];							inform_L[85][0] = l_cell_wire[85];							inform_L[86][0] = l_cell_wire[86];							inform_L[87][0] = l_cell_wire[87];							inform_L[88][0] = l_cell_wire[88];							inform_L[89][0] = l_cell_wire[89];							inform_L[90][0] = l_cell_wire[90];							inform_L[91][0] = l_cell_wire[91];							inform_L[92][0] = l_cell_wire[92];							inform_L[93][0] = l_cell_wire[93];							inform_L[94][0] = l_cell_wire[94];							inform_L[95][0] = l_cell_wire[95];							inform_L[96][0] = l_cell_wire[96];							inform_L[97][0] = l_cell_wire[97];							inform_L[98][0] = l_cell_wire[98];							inform_L[99][0] = l_cell_wire[99];							inform_L[100][0] = l_cell_wire[100];							inform_L[101][0] = l_cell_wire[101];							inform_L[102][0] = l_cell_wire[102];							inform_L[103][0] = l_cell_wire[103];							inform_L[104][0] = l_cell_wire[104];							inform_L[105][0] = l_cell_wire[105];							inform_L[106][0] = l_cell_wire[106];							inform_L[107][0] = l_cell_wire[107];							inform_L[108][0] = l_cell_wire[108];							inform_L[109][0] = l_cell_wire[109];							inform_L[110][0] = l_cell_wire[110];							inform_L[111][0] = l_cell_wire[111];							inform_L[112][0] = l_cell_wire[112];							inform_L[113][0] = l_cell_wire[113];							inform_L[114][0] = l_cell_wire[114];							inform_L[115][0] = l_cell_wire[115];							inform_L[116][0] = l_cell_wire[116];							inform_L[117][0] = l_cell_wire[117];							inform_L[118][0] = l_cell_wire[118];							inform_L[119][0] = l_cell_wire[119];							inform_L[120][0] = l_cell_wire[120];							inform_L[121][0] = l_cell_wire[121];							inform_L[122][0] = l_cell_wire[122];							inform_L[123][0] = l_cell_wire[123];							inform_L[124][0] = l_cell_wire[124];							inform_L[125][0] = l_cell_wire[125];							inform_L[126][0] = l_cell_wire[126];							inform_L[127][0] = l_cell_wire[127];							inform_L[128][0] = l_cell_wire[128];							inform_L[129][0] = l_cell_wire[129];							inform_L[130][0] = l_cell_wire[130];							inform_L[131][0] = l_cell_wire[131];							inform_L[132][0] = l_cell_wire[132];							inform_L[133][0] = l_cell_wire[133];							inform_L[134][0] = l_cell_wire[134];							inform_L[135][0] = l_cell_wire[135];							inform_L[136][0] = l_cell_wire[136];							inform_L[137][0] = l_cell_wire[137];							inform_L[138][0] = l_cell_wire[138];							inform_L[139][0] = l_cell_wire[139];							inform_L[140][0] = l_cell_wire[140];							inform_L[141][0] = l_cell_wire[141];							inform_L[142][0] = l_cell_wire[142];							inform_L[143][0] = l_cell_wire[143];							inform_L[144][0] = l_cell_wire[144];							inform_L[145][0] = l_cell_wire[145];							inform_L[146][0] = l_cell_wire[146];							inform_L[147][0] = l_cell_wire[147];							inform_L[148][0] = l_cell_wire[148];							inform_L[149][0] = l_cell_wire[149];							inform_L[150][0] = l_cell_wire[150];							inform_L[151][0] = l_cell_wire[151];							inform_L[152][0] = l_cell_wire[152];							inform_L[153][0] = l_cell_wire[153];							inform_L[154][0] = l_cell_wire[154];							inform_L[155][0] = l_cell_wire[155];							inform_L[156][0] = l_cell_wire[156];							inform_L[157][0] = l_cell_wire[157];							inform_L[158][0] = l_cell_wire[158];							inform_L[159][0] = l_cell_wire[159];							inform_L[160][0] = l_cell_wire[160];							inform_L[161][0] = l_cell_wire[161];							inform_L[162][0] = l_cell_wire[162];							inform_L[163][0] = l_cell_wire[163];							inform_L[164][0] = l_cell_wire[164];							inform_L[165][0] = l_cell_wire[165];							inform_L[166][0] = l_cell_wire[166];							inform_L[167][0] = l_cell_wire[167];							inform_L[168][0] = l_cell_wire[168];							inform_L[169][0] = l_cell_wire[169];							inform_L[170][0] = l_cell_wire[170];							inform_L[171][0] = l_cell_wire[171];							inform_L[172][0] = l_cell_wire[172];							inform_L[173][0] = l_cell_wire[173];							inform_L[174][0] = l_cell_wire[174];							inform_L[175][0] = l_cell_wire[175];							inform_L[176][0] = l_cell_wire[176];							inform_L[177][0] = l_cell_wire[177];							inform_L[178][0] = l_cell_wire[178];							inform_L[179][0] = l_cell_wire[179];							inform_L[180][0] = l_cell_wire[180];							inform_L[181][0] = l_cell_wire[181];							inform_L[182][0] = l_cell_wire[182];							inform_L[183][0] = l_cell_wire[183];							inform_L[184][0] = l_cell_wire[184];							inform_L[185][0] = l_cell_wire[185];							inform_L[186][0] = l_cell_wire[186];							inform_L[187][0] = l_cell_wire[187];							inform_L[188][0] = l_cell_wire[188];							inform_L[189][0] = l_cell_wire[189];							inform_L[190][0] = l_cell_wire[190];							inform_L[191][0] = l_cell_wire[191];							inform_L[192][0] = l_cell_wire[192];							inform_L[193][0] = l_cell_wire[193];							inform_L[194][0] = l_cell_wire[194];							inform_L[195][0] = l_cell_wire[195];							inform_L[196][0] = l_cell_wire[196];							inform_L[197][0] = l_cell_wire[197];							inform_L[198][0] = l_cell_wire[198];							inform_L[199][0] = l_cell_wire[199];							inform_L[200][0] = l_cell_wire[200];							inform_L[201][0] = l_cell_wire[201];							inform_L[202][0] = l_cell_wire[202];							inform_L[203][0] = l_cell_wire[203];							inform_L[204][0] = l_cell_wire[204];							inform_L[205][0] = l_cell_wire[205];							inform_L[206][0] = l_cell_wire[206];							inform_L[207][0] = l_cell_wire[207];							inform_L[208][0] = l_cell_wire[208];							inform_L[209][0] = l_cell_wire[209];							inform_L[210][0] = l_cell_wire[210];							inform_L[211][0] = l_cell_wire[211];							inform_L[212][0] = l_cell_wire[212];							inform_L[213][0] = l_cell_wire[213];							inform_L[214][0] = l_cell_wire[214];							inform_L[215][0] = l_cell_wire[215];							inform_L[216][0] = l_cell_wire[216];							inform_L[217][0] = l_cell_wire[217];							inform_L[218][0] = l_cell_wire[218];							inform_L[219][0] = l_cell_wire[219];							inform_L[220][0] = l_cell_wire[220];							inform_L[221][0] = l_cell_wire[221];							inform_L[222][0] = l_cell_wire[222];							inform_L[223][0] = l_cell_wire[223];							inform_L[224][0] = l_cell_wire[224];							inform_L[225][0] = l_cell_wire[225];							inform_L[226][0] = l_cell_wire[226];							inform_L[227][0] = l_cell_wire[227];							inform_L[228][0] = l_cell_wire[228];							inform_L[229][0] = l_cell_wire[229];							inform_L[230][0] = l_cell_wire[230];							inform_L[231][0] = l_cell_wire[231];							inform_L[232][0] = l_cell_wire[232];							inform_L[233][0] = l_cell_wire[233];							inform_L[234][0] = l_cell_wire[234];							inform_L[235][0] = l_cell_wire[235];							inform_L[236][0] = l_cell_wire[236];							inform_L[237][0] = l_cell_wire[237];							inform_L[238][0] = l_cell_wire[238];							inform_L[239][0] = l_cell_wire[239];							inform_L[240][0] = l_cell_wire[240];							inform_L[241][0] = l_cell_wire[241];							inform_L[242][0] = l_cell_wire[242];							inform_L[243][0] = l_cell_wire[243];							inform_L[244][0] = l_cell_wire[244];							inform_L[245][0] = l_cell_wire[245];							inform_L[246][0] = l_cell_wire[246];							inform_L[247][0] = l_cell_wire[247];							inform_L[248][0] = l_cell_wire[248];							inform_L[249][0] = l_cell_wire[249];							inform_L[250][0] = l_cell_wire[250];							inform_L[251][0] = l_cell_wire[251];							inform_L[252][0] = l_cell_wire[252];							inform_L[253][0] = l_cell_wire[253];							inform_L[254][0] = l_cell_wire[254];							inform_L[255][0] = l_cell_wire[255];						end
						2:						begin							inform_R[0][2] = r_cell_wire[0];							inform_R[2][2] = r_cell_wire[1];							inform_R[1][2] = r_cell_wire[2];							inform_R[3][2] = r_cell_wire[3];							inform_R[4][2] = r_cell_wire[4];							inform_R[6][2] = r_cell_wire[5];							inform_R[5][2] = r_cell_wire[6];							inform_R[7][2] = r_cell_wire[7];							inform_R[8][2] = r_cell_wire[8];							inform_R[10][2] = r_cell_wire[9];							inform_R[9][2] = r_cell_wire[10];							inform_R[11][2] = r_cell_wire[11];							inform_R[12][2] = r_cell_wire[12];							inform_R[14][2] = r_cell_wire[13];							inform_R[13][2] = r_cell_wire[14];							inform_R[15][2] = r_cell_wire[15];							inform_R[16][2] = r_cell_wire[16];							inform_R[18][2] = r_cell_wire[17];							inform_R[17][2] = r_cell_wire[18];							inform_R[19][2] = r_cell_wire[19];							inform_R[20][2] = r_cell_wire[20];							inform_R[22][2] = r_cell_wire[21];							inform_R[21][2] = r_cell_wire[22];							inform_R[23][2] = r_cell_wire[23];							inform_R[24][2] = r_cell_wire[24];							inform_R[26][2] = r_cell_wire[25];							inform_R[25][2] = r_cell_wire[26];							inform_R[27][2] = r_cell_wire[27];							inform_R[28][2] = r_cell_wire[28];							inform_R[30][2] = r_cell_wire[29];							inform_R[29][2] = r_cell_wire[30];							inform_R[31][2] = r_cell_wire[31];							inform_R[32][2] = r_cell_wire[32];							inform_R[34][2] = r_cell_wire[33];							inform_R[33][2] = r_cell_wire[34];							inform_R[35][2] = r_cell_wire[35];							inform_R[36][2] = r_cell_wire[36];							inform_R[38][2] = r_cell_wire[37];							inform_R[37][2] = r_cell_wire[38];							inform_R[39][2] = r_cell_wire[39];							inform_R[40][2] = r_cell_wire[40];							inform_R[42][2] = r_cell_wire[41];							inform_R[41][2] = r_cell_wire[42];							inform_R[43][2] = r_cell_wire[43];							inform_R[44][2] = r_cell_wire[44];							inform_R[46][2] = r_cell_wire[45];							inform_R[45][2] = r_cell_wire[46];							inform_R[47][2] = r_cell_wire[47];							inform_R[48][2] = r_cell_wire[48];							inform_R[50][2] = r_cell_wire[49];							inform_R[49][2] = r_cell_wire[50];							inform_R[51][2] = r_cell_wire[51];							inform_R[52][2] = r_cell_wire[52];							inform_R[54][2] = r_cell_wire[53];							inform_R[53][2] = r_cell_wire[54];							inform_R[55][2] = r_cell_wire[55];							inform_R[56][2] = r_cell_wire[56];							inform_R[58][2] = r_cell_wire[57];							inform_R[57][2] = r_cell_wire[58];							inform_R[59][2] = r_cell_wire[59];							inform_R[60][2] = r_cell_wire[60];							inform_R[62][2] = r_cell_wire[61];							inform_R[61][2] = r_cell_wire[62];							inform_R[63][2] = r_cell_wire[63];							inform_R[64][2] = r_cell_wire[64];							inform_R[66][2] = r_cell_wire[65];							inform_R[65][2] = r_cell_wire[66];							inform_R[67][2] = r_cell_wire[67];							inform_R[68][2] = r_cell_wire[68];							inform_R[70][2] = r_cell_wire[69];							inform_R[69][2] = r_cell_wire[70];							inform_R[71][2] = r_cell_wire[71];							inform_R[72][2] = r_cell_wire[72];							inform_R[74][2] = r_cell_wire[73];							inform_R[73][2] = r_cell_wire[74];							inform_R[75][2] = r_cell_wire[75];							inform_R[76][2] = r_cell_wire[76];							inform_R[78][2] = r_cell_wire[77];							inform_R[77][2] = r_cell_wire[78];							inform_R[79][2] = r_cell_wire[79];							inform_R[80][2] = r_cell_wire[80];							inform_R[82][2] = r_cell_wire[81];							inform_R[81][2] = r_cell_wire[82];							inform_R[83][2] = r_cell_wire[83];							inform_R[84][2] = r_cell_wire[84];							inform_R[86][2] = r_cell_wire[85];							inform_R[85][2] = r_cell_wire[86];							inform_R[87][2] = r_cell_wire[87];							inform_R[88][2] = r_cell_wire[88];							inform_R[90][2] = r_cell_wire[89];							inform_R[89][2] = r_cell_wire[90];							inform_R[91][2] = r_cell_wire[91];							inform_R[92][2] = r_cell_wire[92];							inform_R[94][2] = r_cell_wire[93];							inform_R[93][2] = r_cell_wire[94];							inform_R[95][2] = r_cell_wire[95];							inform_R[96][2] = r_cell_wire[96];							inform_R[98][2] = r_cell_wire[97];							inform_R[97][2] = r_cell_wire[98];							inform_R[99][2] = r_cell_wire[99];							inform_R[100][2] = r_cell_wire[100];							inform_R[102][2] = r_cell_wire[101];							inform_R[101][2] = r_cell_wire[102];							inform_R[103][2] = r_cell_wire[103];							inform_R[104][2] = r_cell_wire[104];							inform_R[106][2] = r_cell_wire[105];							inform_R[105][2] = r_cell_wire[106];							inform_R[107][2] = r_cell_wire[107];							inform_R[108][2] = r_cell_wire[108];							inform_R[110][2] = r_cell_wire[109];							inform_R[109][2] = r_cell_wire[110];							inform_R[111][2] = r_cell_wire[111];							inform_R[112][2] = r_cell_wire[112];							inform_R[114][2] = r_cell_wire[113];							inform_R[113][2] = r_cell_wire[114];							inform_R[115][2] = r_cell_wire[115];							inform_R[116][2] = r_cell_wire[116];							inform_R[118][2] = r_cell_wire[117];							inform_R[117][2] = r_cell_wire[118];							inform_R[119][2] = r_cell_wire[119];							inform_R[120][2] = r_cell_wire[120];							inform_R[122][2] = r_cell_wire[121];							inform_R[121][2] = r_cell_wire[122];							inform_R[123][2] = r_cell_wire[123];							inform_R[124][2] = r_cell_wire[124];							inform_R[126][2] = r_cell_wire[125];							inform_R[125][2] = r_cell_wire[126];							inform_R[127][2] = r_cell_wire[127];							inform_R[128][2] = r_cell_wire[128];							inform_R[130][2] = r_cell_wire[129];							inform_R[129][2] = r_cell_wire[130];							inform_R[131][2] = r_cell_wire[131];							inform_R[132][2] = r_cell_wire[132];							inform_R[134][2] = r_cell_wire[133];							inform_R[133][2] = r_cell_wire[134];							inform_R[135][2] = r_cell_wire[135];							inform_R[136][2] = r_cell_wire[136];							inform_R[138][2] = r_cell_wire[137];							inform_R[137][2] = r_cell_wire[138];							inform_R[139][2] = r_cell_wire[139];							inform_R[140][2] = r_cell_wire[140];							inform_R[142][2] = r_cell_wire[141];							inform_R[141][2] = r_cell_wire[142];							inform_R[143][2] = r_cell_wire[143];							inform_R[144][2] = r_cell_wire[144];							inform_R[146][2] = r_cell_wire[145];							inform_R[145][2] = r_cell_wire[146];							inform_R[147][2] = r_cell_wire[147];							inform_R[148][2] = r_cell_wire[148];							inform_R[150][2] = r_cell_wire[149];							inform_R[149][2] = r_cell_wire[150];							inform_R[151][2] = r_cell_wire[151];							inform_R[152][2] = r_cell_wire[152];							inform_R[154][2] = r_cell_wire[153];							inform_R[153][2] = r_cell_wire[154];							inform_R[155][2] = r_cell_wire[155];							inform_R[156][2] = r_cell_wire[156];							inform_R[158][2] = r_cell_wire[157];							inform_R[157][2] = r_cell_wire[158];							inform_R[159][2] = r_cell_wire[159];							inform_R[160][2] = r_cell_wire[160];							inform_R[162][2] = r_cell_wire[161];							inform_R[161][2] = r_cell_wire[162];							inform_R[163][2] = r_cell_wire[163];							inform_R[164][2] = r_cell_wire[164];							inform_R[166][2] = r_cell_wire[165];							inform_R[165][2] = r_cell_wire[166];							inform_R[167][2] = r_cell_wire[167];							inform_R[168][2] = r_cell_wire[168];							inform_R[170][2] = r_cell_wire[169];							inform_R[169][2] = r_cell_wire[170];							inform_R[171][2] = r_cell_wire[171];							inform_R[172][2] = r_cell_wire[172];							inform_R[174][2] = r_cell_wire[173];							inform_R[173][2] = r_cell_wire[174];							inform_R[175][2] = r_cell_wire[175];							inform_R[176][2] = r_cell_wire[176];							inform_R[178][2] = r_cell_wire[177];							inform_R[177][2] = r_cell_wire[178];							inform_R[179][2] = r_cell_wire[179];							inform_R[180][2] = r_cell_wire[180];							inform_R[182][2] = r_cell_wire[181];							inform_R[181][2] = r_cell_wire[182];							inform_R[183][2] = r_cell_wire[183];							inform_R[184][2] = r_cell_wire[184];							inform_R[186][2] = r_cell_wire[185];							inform_R[185][2] = r_cell_wire[186];							inform_R[187][2] = r_cell_wire[187];							inform_R[188][2] = r_cell_wire[188];							inform_R[190][2] = r_cell_wire[189];							inform_R[189][2] = r_cell_wire[190];							inform_R[191][2] = r_cell_wire[191];							inform_R[192][2] = r_cell_wire[192];							inform_R[194][2] = r_cell_wire[193];							inform_R[193][2] = r_cell_wire[194];							inform_R[195][2] = r_cell_wire[195];							inform_R[196][2] = r_cell_wire[196];							inform_R[198][2] = r_cell_wire[197];							inform_R[197][2] = r_cell_wire[198];							inform_R[199][2] = r_cell_wire[199];							inform_R[200][2] = r_cell_wire[200];							inform_R[202][2] = r_cell_wire[201];							inform_R[201][2] = r_cell_wire[202];							inform_R[203][2] = r_cell_wire[203];							inform_R[204][2] = r_cell_wire[204];							inform_R[206][2] = r_cell_wire[205];							inform_R[205][2] = r_cell_wire[206];							inform_R[207][2] = r_cell_wire[207];							inform_R[208][2] = r_cell_wire[208];							inform_R[210][2] = r_cell_wire[209];							inform_R[209][2] = r_cell_wire[210];							inform_R[211][2] = r_cell_wire[211];							inform_R[212][2] = r_cell_wire[212];							inform_R[214][2] = r_cell_wire[213];							inform_R[213][2] = r_cell_wire[214];							inform_R[215][2] = r_cell_wire[215];							inform_R[216][2] = r_cell_wire[216];							inform_R[218][2] = r_cell_wire[217];							inform_R[217][2] = r_cell_wire[218];							inform_R[219][2] = r_cell_wire[219];							inform_R[220][2] = r_cell_wire[220];							inform_R[222][2] = r_cell_wire[221];							inform_R[221][2] = r_cell_wire[222];							inform_R[223][2] = r_cell_wire[223];							inform_R[224][2] = r_cell_wire[224];							inform_R[226][2] = r_cell_wire[225];							inform_R[225][2] = r_cell_wire[226];							inform_R[227][2] = r_cell_wire[227];							inform_R[228][2] = r_cell_wire[228];							inform_R[230][2] = r_cell_wire[229];							inform_R[229][2] = r_cell_wire[230];							inform_R[231][2] = r_cell_wire[231];							inform_R[232][2] = r_cell_wire[232];							inform_R[234][2] = r_cell_wire[233];							inform_R[233][2] = r_cell_wire[234];							inform_R[235][2] = r_cell_wire[235];							inform_R[236][2] = r_cell_wire[236];							inform_R[238][2] = r_cell_wire[237];							inform_R[237][2] = r_cell_wire[238];							inform_R[239][2] = r_cell_wire[239];							inform_R[240][2] = r_cell_wire[240];							inform_R[242][2] = r_cell_wire[241];							inform_R[241][2] = r_cell_wire[242];							inform_R[243][2] = r_cell_wire[243];							inform_R[244][2] = r_cell_wire[244];							inform_R[246][2] = r_cell_wire[245];							inform_R[245][2] = r_cell_wire[246];							inform_R[247][2] = r_cell_wire[247];							inform_R[248][2] = r_cell_wire[248];							inform_R[250][2] = r_cell_wire[249];							inform_R[249][2] = r_cell_wire[250];							inform_R[251][2] = r_cell_wire[251];							inform_R[252][2] = r_cell_wire[252];							inform_R[254][2] = r_cell_wire[253];							inform_R[253][2] = r_cell_wire[254];							inform_R[255][2] = r_cell_wire[255];							inform_L[0][1] = l_cell_wire[0];							inform_L[2][1] = l_cell_wire[1];							inform_L[1][1] = l_cell_wire[2];							inform_L[3][1] = l_cell_wire[3];							inform_L[4][1] = l_cell_wire[4];							inform_L[6][1] = l_cell_wire[5];							inform_L[5][1] = l_cell_wire[6];							inform_L[7][1] = l_cell_wire[7];							inform_L[8][1] = l_cell_wire[8];							inform_L[10][1] = l_cell_wire[9];							inform_L[9][1] = l_cell_wire[10];							inform_L[11][1] = l_cell_wire[11];							inform_L[12][1] = l_cell_wire[12];							inform_L[14][1] = l_cell_wire[13];							inform_L[13][1] = l_cell_wire[14];							inform_L[15][1] = l_cell_wire[15];							inform_L[16][1] = l_cell_wire[16];							inform_L[18][1] = l_cell_wire[17];							inform_L[17][1] = l_cell_wire[18];							inform_L[19][1] = l_cell_wire[19];							inform_L[20][1] = l_cell_wire[20];							inform_L[22][1] = l_cell_wire[21];							inform_L[21][1] = l_cell_wire[22];							inform_L[23][1] = l_cell_wire[23];							inform_L[24][1] = l_cell_wire[24];							inform_L[26][1] = l_cell_wire[25];							inform_L[25][1] = l_cell_wire[26];							inform_L[27][1] = l_cell_wire[27];							inform_L[28][1] = l_cell_wire[28];							inform_L[30][1] = l_cell_wire[29];							inform_L[29][1] = l_cell_wire[30];							inform_L[31][1] = l_cell_wire[31];							inform_L[32][1] = l_cell_wire[32];							inform_L[34][1] = l_cell_wire[33];							inform_L[33][1] = l_cell_wire[34];							inform_L[35][1] = l_cell_wire[35];							inform_L[36][1] = l_cell_wire[36];							inform_L[38][1] = l_cell_wire[37];							inform_L[37][1] = l_cell_wire[38];							inform_L[39][1] = l_cell_wire[39];							inform_L[40][1] = l_cell_wire[40];							inform_L[42][1] = l_cell_wire[41];							inform_L[41][1] = l_cell_wire[42];							inform_L[43][1] = l_cell_wire[43];							inform_L[44][1] = l_cell_wire[44];							inform_L[46][1] = l_cell_wire[45];							inform_L[45][1] = l_cell_wire[46];							inform_L[47][1] = l_cell_wire[47];							inform_L[48][1] = l_cell_wire[48];							inform_L[50][1] = l_cell_wire[49];							inform_L[49][1] = l_cell_wire[50];							inform_L[51][1] = l_cell_wire[51];							inform_L[52][1] = l_cell_wire[52];							inform_L[54][1] = l_cell_wire[53];							inform_L[53][1] = l_cell_wire[54];							inform_L[55][1] = l_cell_wire[55];							inform_L[56][1] = l_cell_wire[56];							inform_L[58][1] = l_cell_wire[57];							inform_L[57][1] = l_cell_wire[58];							inform_L[59][1] = l_cell_wire[59];							inform_L[60][1] = l_cell_wire[60];							inform_L[62][1] = l_cell_wire[61];							inform_L[61][1] = l_cell_wire[62];							inform_L[63][1] = l_cell_wire[63];							inform_L[64][1] = l_cell_wire[64];							inform_L[66][1] = l_cell_wire[65];							inform_L[65][1] = l_cell_wire[66];							inform_L[67][1] = l_cell_wire[67];							inform_L[68][1] = l_cell_wire[68];							inform_L[70][1] = l_cell_wire[69];							inform_L[69][1] = l_cell_wire[70];							inform_L[71][1] = l_cell_wire[71];							inform_L[72][1] = l_cell_wire[72];							inform_L[74][1] = l_cell_wire[73];							inform_L[73][1] = l_cell_wire[74];							inform_L[75][1] = l_cell_wire[75];							inform_L[76][1] = l_cell_wire[76];							inform_L[78][1] = l_cell_wire[77];							inform_L[77][1] = l_cell_wire[78];							inform_L[79][1] = l_cell_wire[79];							inform_L[80][1] = l_cell_wire[80];							inform_L[82][1] = l_cell_wire[81];							inform_L[81][1] = l_cell_wire[82];							inform_L[83][1] = l_cell_wire[83];							inform_L[84][1] = l_cell_wire[84];							inform_L[86][1] = l_cell_wire[85];							inform_L[85][1] = l_cell_wire[86];							inform_L[87][1] = l_cell_wire[87];							inform_L[88][1] = l_cell_wire[88];							inform_L[90][1] = l_cell_wire[89];							inform_L[89][1] = l_cell_wire[90];							inform_L[91][1] = l_cell_wire[91];							inform_L[92][1] = l_cell_wire[92];							inform_L[94][1] = l_cell_wire[93];							inform_L[93][1] = l_cell_wire[94];							inform_L[95][1] = l_cell_wire[95];							inform_L[96][1] = l_cell_wire[96];							inform_L[98][1] = l_cell_wire[97];							inform_L[97][1] = l_cell_wire[98];							inform_L[99][1] = l_cell_wire[99];							inform_L[100][1] = l_cell_wire[100];							inform_L[102][1] = l_cell_wire[101];							inform_L[101][1] = l_cell_wire[102];							inform_L[103][1] = l_cell_wire[103];							inform_L[104][1] = l_cell_wire[104];							inform_L[106][1] = l_cell_wire[105];							inform_L[105][1] = l_cell_wire[106];							inform_L[107][1] = l_cell_wire[107];							inform_L[108][1] = l_cell_wire[108];							inform_L[110][1] = l_cell_wire[109];							inform_L[109][1] = l_cell_wire[110];							inform_L[111][1] = l_cell_wire[111];							inform_L[112][1] = l_cell_wire[112];							inform_L[114][1] = l_cell_wire[113];							inform_L[113][1] = l_cell_wire[114];							inform_L[115][1] = l_cell_wire[115];							inform_L[116][1] = l_cell_wire[116];							inform_L[118][1] = l_cell_wire[117];							inform_L[117][1] = l_cell_wire[118];							inform_L[119][1] = l_cell_wire[119];							inform_L[120][1] = l_cell_wire[120];							inform_L[122][1] = l_cell_wire[121];							inform_L[121][1] = l_cell_wire[122];							inform_L[123][1] = l_cell_wire[123];							inform_L[124][1] = l_cell_wire[124];							inform_L[126][1] = l_cell_wire[125];							inform_L[125][1] = l_cell_wire[126];							inform_L[127][1] = l_cell_wire[127];							inform_L[128][1] = l_cell_wire[128];							inform_L[130][1] = l_cell_wire[129];							inform_L[129][1] = l_cell_wire[130];							inform_L[131][1] = l_cell_wire[131];							inform_L[132][1] = l_cell_wire[132];							inform_L[134][1] = l_cell_wire[133];							inform_L[133][1] = l_cell_wire[134];							inform_L[135][1] = l_cell_wire[135];							inform_L[136][1] = l_cell_wire[136];							inform_L[138][1] = l_cell_wire[137];							inform_L[137][1] = l_cell_wire[138];							inform_L[139][1] = l_cell_wire[139];							inform_L[140][1] = l_cell_wire[140];							inform_L[142][1] = l_cell_wire[141];							inform_L[141][1] = l_cell_wire[142];							inform_L[143][1] = l_cell_wire[143];							inform_L[144][1] = l_cell_wire[144];							inform_L[146][1] = l_cell_wire[145];							inform_L[145][1] = l_cell_wire[146];							inform_L[147][1] = l_cell_wire[147];							inform_L[148][1] = l_cell_wire[148];							inform_L[150][1] = l_cell_wire[149];							inform_L[149][1] = l_cell_wire[150];							inform_L[151][1] = l_cell_wire[151];							inform_L[152][1] = l_cell_wire[152];							inform_L[154][1] = l_cell_wire[153];							inform_L[153][1] = l_cell_wire[154];							inform_L[155][1] = l_cell_wire[155];							inform_L[156][1] = l_cell_wire[156];							inform_L[158][1] = l_cell_wire[157];							inform_L[157][1] = l_cell_wire[158];							inform_L[159][1] = l_cell_wire[159];							inform_L[160][1] = l_cell_wire[160];							inform_L[162][1] = l_cell_wire[161];							inform_L[161][1] = l_cell_wire[162];							inform_L[163][1] = l_cell_wire[163];							inform_L[164][1] = l_cell_wire[164];							inform_L[166][1] = l_cell_wire[165];							inform_L[165][1] = l_cell_wire[166];							inform_L[167][1] = l_cell_wire[167];							inform_L[168][1] = l_cell_wire[168];							inform_L[170][1] = l_cell_wire[169];							inform_L[169][1] = l_cell_wire[170];							inform_L[171][1] = l_cell_wire[171];							inform_L[172][1] = l_cell_wire[172];							inform_L[174][1] = l_cell_wire[173];							inform_L[173][1] = l_cell_wire[174];							inform_L[175][1] = l_cell_wire[175];							inform_L[176][1] = l_cell_wire[176];							inform_L[178][1] = l_cell_wire[177];							inform_L[177][1] = l_cell_wire[178];							inform_L[179][1] = l_cell_wire[179];							inform_L[180][1] = l_cell_wire[180];							inform_L[182][1] = l_cell_wire[181];							inform_L[181][1] = l_cell_wire[182];							inform_L[183][1] = l_cell_wire[183];							inform_L[184][1] = l_cell_wire[184];							inform_L[186][1] = l_cell_wire[185];							inform_L[185][1] = l_cell_wire[186];							inform_L[187][1] = l_cell_wire[187];							inform_L[188][1] = l_cell_wire[188];							inform_L[190][1] = l_cell_wire[189];							inform_L[189][1] = l_cell_wire[190];							inform_L[191][1] = l_cell_wire[191];							inform_L[192][1] = l_cell_wire[192];							inform_L[194][1] = l_cell_wire[193];							inform_L[193][1] = l_cell_wire[194];							inform_L[195][1] = l_cell_wire[195];							inform_L[196][1] = l_cell_wire[196];							inform_L[198][1] = l_cell_wire[197];							inform_L[197][1] = l_cell_wire[198];							inform_L[199][1] = l_cell_wire[199];							inform_L[200][1] = l_cell_wire[200];							inform_L[202][1] = l_cell_wire[201];							inform_L[201][1] = l_cell_wire[202];							inform_L[203][1] = l_cell_wire[203];							inform_L[204][1] = l_cell_wire[204];							inform_L[206][1] = l_cell_wire[205];							inform_L[205][1] = l_cell_wire[206];							inform_L[207][1] = l_cell_wire[207];							inform_L[208][1] = l_cell_wire[208];							inform_L[210][1] = l_cell_wire[209];							inform_L[209][1] = l_cell_wire[210];							inform_L[211][1] = l_cell_wire[211];							inform_L[212][1] = l_cell_wire[212];							inform_L[214][1] = l_cell_wire[213];							inform_L[213][1] = l_cell_wire[214];							inform_L[215][1] = l_cell_wire[215];							inform_L[216][1] = l_cell_wire[216];							inform_L[218][1] = l_cell_wire[217];							inform_L[217][1] = l_cell_wire[218];							inform_L[219][1] = l_cell_wire[219];							inform_L[220][1] = l_cell_wire[220];							inform_L[222][1] = l_cell_wire[221];							inform_L[221][1] = l_cell_wire[222];							inform_L[223][1] = l_cell_wire[223];							inform_L[224][1] = l_cell_wire[224];							inform_L[226][1] = l_cell_wire[225];							inform_L[225][1] = l_cell_wire[226];							inform_L[227][1] = l_cell_wire[227];							inform_L[228][1] = l_cell_wire[228];							inform_L[230][1] = l_cell_wire[229];							inform_L[229][1] = l_cell_wire[230];							inform_L[231][1] = l_cell_wire[231];							inform_L[232][1] = l_cell_wire[232];							inform_L[234][1] = l_cell_wire[233];							inform_L[233][1] = l_cell_wire[234];							inform_L[235][1] = l_cell_wire[235];							inform_L[236][1] = l_cell_wire[236];							inform_L[238][1] = l_cell_wire[237];							inform_L[237][1] = l_cell_wire[238];							inform_L[239][1] = l_cell_wire[239];							inform_L[240][1] = l_cell_wire[240];							inform_L[242][1] = l_cell_wire[241];							inform_L[241][1] = l_cell_wire[242];							inform_L[243][1] = l_cell_wire[243];							inform_L[244][1] = l_cell_wire[244];							inform_L[246][1] = l_cell_wire[245];							inform_L[245][1] = l_cell_wire[246];							inform_L[247][1] = l_cell_wire[247];							inform_L[248][1] = l_cell_wire[248];							inform_L[250][1] = l_cell_wire[249];							inform_L[249][1] = l_cell_wire[250];							inform_L[251][1] = l_cell_wire[251];							inform_L[252][1] = l_cell_wire[252];							inform_L[254][1] = l_cell_wire[253];							inform_L[253][1] = l_cell_wire[254];							inform_L[255][1] = l_cell_wire[255];						end
						3:						begin							inform_R[0][3] = r_cell_wire[0];							inform_R[4][3] = r_cell_wire[1];							inform_R[1][3] = r_cell_wire[2];							inform_R[5][3] = r_cell_wire[3];							inform_R[2][3] = r_cell_wire[4];							inform_R[6][3] = r_cell_wire[5];							inform_R[3][3] = r_cell_wire[6];							inform_R[7][3] = r_cell_wire[7];							inform_R[8][3] = r_cell_wire[8];							inform_R[12][3] = r_cell_wire[9];							inform_R[9][3] = r_cell_wire[10];							inform_R[13][3] = r_cell_wire[11];							inform_R[10][3] = r_cell_wire[12];							inform_R[14][3] = r_cell_wire[13];							inform_R[11][3] = r_cell_wire[14];							inform_R[15][3] = r_cell_wire[15];							inform_R[16][3] = r_cell_wire[16];							inform_R[20][3] = r_cell_wire[17];							inform_R[17][3] = r_cell_wire[18];							inform_R[21][3] = r_cell_wire[19];							inform_R[18][3] = r_cell_wire[20];							inform_R[22][3] = r_cell_wire[21];							inform_R[19][3] = r_cell_wire[22];							inform_R[23][3] = r_cell_wire[23];							inform_R[24][3] = r_cell_wire[24];							inform_R[28][3] = r_cell_wire[25];							inform_R[25][3] = r_cell_wire[26];							inform_R[29][3] = r_cell_wire[27];							inform_R[26][3] = r_cell_wire[28];							inform_R[30][3] = r_cell_wire[29];							inform_R[27][3] = r_cell_wire[30];							inform_R[31][3] = r_cell_wire[31];							inform_R[32][3] = r_cell_wire[32];							inform_R[36][3] = r_cell_wire[33];							inform_R[33][3] = r_cell_wire[34];							inform_R[37][3] = r_cell_wire[35];							inform_R[34][3] = r_cell_wire[36];							inform_R[38][3] = r_cell_wire[37];							inform_R[35][3] = r_cell_wire[38];							inform_R[39][3] = r_cell_wire[39];							inform_R[40][3] = r_cell_wire[40];							inform_R[44][3] = r_cell_wire[41];							inform_R[41][3] = r_cell_wire[42];							inform_R[45][3] = r_cell_wire[43];							inform_R[42][3] = r_cell_wire[44];							inform_R[46][3] = r_cell_wire[45];							inform_R[43][3] = r_cell_wire[46];							inform_R[47][3] = r_cell_wire[47];							inform_R[48][3] = r_cell_wire[48];							inform_R[52][3] = r_cell_wire[49];							inform_R[49][3] = r_cell_wire[50];							inform_R[53][3] = r_cell_wire[51];							inform_R[50][3] = r_cell_wire[52];							inform_R[54][3] = r_cell_wire[53];							inform_R[51][3] = r_cell_wire[54];							inform_R[55][3] = r_cell_wire[55];							inform_R[56][3] = r_cell_wire[56];							inform_R[60][3] = r_cell_wire[57];							inform_R[57][3] = r_cell_wire[58];							inform_R[61][3] = r_cell_wire[59];							inform_R[58][3] = r_cell_wire[60];							inform_R[62][3] = r_cell_wire[61];							inform_R[59][3] = r_cell_wire[62];							inform_R[63][3] = r_cell_wire[63];							inform_R[64][3] = r_cell_wire[64];							inform_R[68][3] = r_cell_wire[65];							inform_R[65][3] = r_cell_wire[66];							inform_R[69][3] = r_cell_wire[67];							inform_R[66][3] = r_cell_wire[68];							inform_R[70][3] = r_cell_wire[69];							inform_R[67][3] = r_cell_wire[70];							inform_R[71][3] = r_cell_wire[71];							inform_R[72][3] = r_cell_wire[72];							inform_R[76][3] = r_cell_wire[73];							inform_R[73][3] = r_cell_wire[74];							inform_R[77][3] = r_cell_wire[75];							inform_R[74][3] = r_cell_wire[76];							inform_R[78][3] = r_cell_wire[77];							inform_R[75][3] = r_cell_wire[78];							inform_R[79][3] = r_cell_wire[79];							inform_R[80][3] = r_cell_wire[80];							inform_R[84][3] = r_cell_wire[81];							inform_R[81][3] = r_cell_wire[82];							inform_R[85][3] = r_cell_wire[83];							inform_R[82][3] = r_cell_wire[84];							inform_R[86][3] = r_cell_wire[85];							inform_R[83][3] = r_cell_wire[86];							inform_R[87][3] = r_cell_wire[87];							inform_R[88][3] = r_cell_wire[88];							inform_R[92][3] = r_cell_wire[89];							inform_R[89][3] = r_cell_wire[90];							inform_R[93][3] = r_cell_wire[91];							inform_R[90][3] = r_cell_wire[92];							inform_R[94][3] = r_cell_wire[93];							inform_R[91][3] = r_cell_wire[94];							inform_R[95][3] = r_cell_wire[95];							inform_R[96][3] = r_cell_wire[96];							inform_R[100][3] = r_cell_wire[97];							inform_R[97][3] = r_cell_wire[98];							inform_R[101][3] = r_cell_wire[99];							inform_R[98][3] = r_cell_wire[100];							inform_R[102][3] = r_cell_wire[101];							inform_R[99][3] = r_cell_wire[102];							inform_R[103][3] = r_cell_wire[103];							inform_R[104][3] = r_cell_wire[104];							inform_R[108][3] = r_cell_wire[105];							inform_R[105][3] = r_cell_wire[106];							inform_R[109][3] = r_cell_wire[107];							inform_R[106][3] = r_cell_wire[108];							inform_R[110][3] = r_cell_wire[109];							inform_R[107][3] = r_cell_wire[110];							inform_R[111][3] = r_cell_wire[111];							inform_R[112][3] = r_cell_wire[112];							inform_R[116][3] = r_cell_wire[113];							inform_R[113][3] = r_cell_wire[114];							inform_R[117][3] = r_cell_wire[115];							inform_R[114][3] = r_cell_wire[116];							inform_R[118][3] = r_cell_wire[117];							inform_R[115][3] = r_cell_wire[118];							inform_R[119][3] = r_cell_wire[119];							inform_R[120][3] = r_cell_wire[120];							inform_R[124][3] = r_cell_wire[121];							inform_R[121][3] = r_cell_wire[122];							inform_R[125][3] = r_cell_wire[123];							inform_R[122][3] = r_cell_wire[124];							inform_R[126][3] = r_cell_wire[125];							inform_R[123][3] = r_cell_wire[126];							inform_R[127][3] = r_cell_wire[127];							inform_R[128][3] = r_cell_wire[128];							inform_R[132][3] = r_cell_wire[129];							inform_R[129][3] = r_cell_wire[130];							inform_R[133][3] = r_cell_wire[131];							inform_R[130][3] = r_cell_wire[132];							inform_R[134][3] = r_cell_wire[133];							inform_R[131][3] = r_cell_wire[134];							inform_R[135][3] = r_cell_wire[135];							inform_R[136][3] = r_cell_wire[136];							inform_R[140][3] = r_cell_wire[137];							inform_R[137][3] = r_cell_wire[138];							inform_R[141][3] = r_cell_wire[139];							inform_R[138][3] = r_cell_wire[140];							inform_R[142][3] = r_cell_wire[141];							inform_R[139][3] = r_cell_wire[142];							inform_R[143][3] = r_cell_wire[143];							inform_R[144][3] = r_cell_wire[144];							inform_R[148][3] = r_cell_wire[145];							inform_R[145][3] = r_cell_wire[146];							inform_R[149][3] = r_cell_wire[147];							inform_R[146][3] = r_cell_wire[148];							inform_R[150][3] = r_cell_wire[149];							inform_R[147][3] = r_cell_wire[150];							inform_R[151][3] = r_cell_wire[151];							inform_R[152][3] = r_cell_wire[152];							inform_R[156][3] = r_cell_wire[153];							inform_R[153][3] = r_cell_wire[154];							inform_R[157][3] = r_cell_wire[155];							inform_R[154][3] = r_cell_wire[156];							inform_R[158][3] = r_cell_wire[157];							inform_R[155][3] = r_cell_wire[158];							inform_R[159][3] = r_cell_wire[159];							inform_R[160][3] = r_cell_wire[160];							inform_R[164][3] = r_cell_wire[161];							inform_R[161][3] = r_cell_wire[162];							inform_R[165][3] = r_cell_wire[163];							inform_R[162][3] = r_cell_wire[164];							inform_R[166][3] = r_cell_wire[165];							inform_R[163][3] = r_cell_wire[166];							inform_R[167][3] = r_cell_wire[167];							inform_R[168][3] = r_cell_wire[168];							inform_R[172][3] = r_cell_wire[169];							inform_R[169][3] = r_cell_wire[170];							inform_R[173][3] = r_cell_wire[171];							inform_R[170][3] = r_cell_wire[172];							inform_R[174][3] = r_cell_wire[173];							inform_R[171][3] = r_cell_wire[174];							inform_R[175][3] = r_cell_wire[175];							inform_R[176][3] = r_cell_wire[176];							inform_R[180][3] = r_cell_wire[177];							inform_R[177][3] = r_cell_wire[178];							inform_R[181][3] = r_cell_wire[179];							inform_R[178][3] = r_cell_wire[180];							inform_R[182][3] = r_cell_wire[181];							inform_R[179][3] = r_cell_wire[182];							inform_R[183][3] = r_cell_wire[183];							inform_R[184][3] = r_cell_wire[184];							inform_R[188][3] = r_cell_wire[185];							inform_R[185][3] = r_cell_wire[186];							inform_R[189][3] = r_cell_wire[187];							inform_R[186][3] = r_cell_wire[188];							inform_R[190][3] = r_cell_wire[189];							inform_R[187][3] = r_cell_wire[190];							inform_R[191][3] = r_cell_wire[191];							inform_R[192][3] = r_cell_wire[192];							inform_R[196][3] = r_cell_wire[193];							inform_R[193][3] = r_cell_wire[194];							inform_R[197][3] = r_cell_wire[195];							inform_R[194][3] = r_cell_wire[196];							inform_R[198][3] = r_cell_wire[197];							inform_R[195][3] = r_cell_wire[198];							inform_R[199][3] = r_cell_wire[199];							inform_R[200][3] = r_cell_wire[200];							inform_R[204][3] = r_cell_wire[201];							inform_R[201][3] = r_cell_wire[202];							inform_R[205][3] = r_cell_wire[203];							inform_R[202][3] = r_cell_wire[204];							inform_R[206][3] = r_cell_wire[205];							inform_R[203][3] = r_cell_wire[206];							inform_R[207][3] = r_cell_wire[207];							inform_R[208][3] = r_cell_wire[208];							inform_R[212][3] = r_cell_wire[209];							inform_R[209][3] = r_cell_wire[210];							inform_R[213][3] = r_cell_wire[211];							inform_R[210][3] = r_cell_wire[212];							inform_R[214][3] = r_cell_wire[213];							inform_R[211][3] = r_cell_wire[214];							inform_R[215][3] = r_cell_wire[215];							inform_R[216][3] = r_cell_wire[216];							inform_R[220][3] = r_cell_wire[217];							inform_R[217][3] = r_cell_wire[218];							inform_R[221][3] = r_cell_wire[219];							inform_R[218][3] = r_cell_wire[220];							inform_R[222][3] = r_cell_wire[221];							inform_R[219][3] = r_cell_wire[222];							inform_R[223][3] = r_cell_wire[223];							inform_R[224][3] = r_cell_wire[224];							inform_R[228][3] = r_cell_wire[225];							inform_R[225][3] = r_cell_wire[226];							inform_R[229][3] = r_cell_wire[227];							inform_R[226][3] = r_cell_wire[228];							inform_R[230][3] = r_cell_wire[229];							inform_R[227][3] = r_cell_wire[230];							inform_R[231][3] = r_cell_wire[231];							inform_R[232][3] = r_cell_wire[232];							inform_R[236][3] = r_cell_wire[233];							inform_R[233][3] = r_cell_wire[234];							inform_R[237][3] = r_cell_wire[235];							inform_R[234][3] = r_cell_wire[236];							inform_R[238][3] = r_cell_wire[237];							inform_R[235][3] = r_cell_wire[238];							inform_R[239][3] = r_cell_wire[239];							inform_R[240][3] = r_cell_wire[240];							inform_R[244][3] = r_cell_wire[241];							inform_R[241][3] = r_cell_wire[242];							inform_R[245][3] = r_cell_wire[243];							inform_R[242][3] = r_cell_wire[244];							inform_R[246][3] = r_cell_wire[245];							inform_R[243][3] = r_cell_wire[246];							inform_R[247][3] = r_cell_wire[247];							inform_R[248][3] = r_cell_wire[248];							inform_R[252][3] = r_cell_wire[249];							inform_R[249][3] = r_cell_wire[250];							inform_R[253][3] = r_cell_wire[251];							inform_R[250][3] = r_cell_wire[252];							inform_R[254][3] = r_cell_wire[253];							inform_R[251][3] = r_cell_wire[254];							inform_R[255][3] = r_cell_wire[255];							inform_L[0][2] = l_cell_wire[0];							inform_L[4][2] = l_cell_wire[1];							inform_L[1][2] = l_cell_wire[2];							inform_L[5][2] = l_cell_wire[3];							inform_L[2][2] = l_cell_wire[4];							inform_L[6][2] = l_cell_wire[5];							inform_L[3][2] = l_cell_wire[6];							inform_L[7][2] = l_cell_wire[7];							inform_L[8][2] = l_cell_wire[8];							inform_L[12][2] = l_cell_wire[9];							inform_L[9][2] = l_cell_wire[10];							inform_L[13][2] = l_cell_wire[11];							inform_L[10][2] = l_cell_wire[12];							inform_L[14][2] = l_cell_wire[13];							inform_L[11][2] = l_cell_wire[14];							inform_L[15][2] = l_cell_wire[15];							inform_L[16][2] = l_cell_wire[16];							inform_L[20][2] = l_cell_wire[17];							inform_L[17][2] = l_cell_wire[18];							inform_L[21][2] = l_cell_wire[19];							inform_L[18][2] = l_cell_wire[20];							inform_L[22][2] = l_cell_wire[21];							inform_L[19][2] = l_cell_wire[22];							inform_L[23][2] = l_cell_wire[23];							inform_L[24][2] = l_cell_wire[24];							inform_L[28][2] = l_cell_wire[25];							inform_L[25][2] = l_cell_wire[26];							inform_L[29][2] = l_cell_wire[27];							inform_L[26][2] = l_cell_wire[28];							inform_L[30][2] = l_cell_wire[29];							inform_L[27][2] = l_cell_wire[30];							inform_L[31][2] = l_cell_wire[31];							inform_L[32][2] = l_cell_wire[32];							inform_L[36][2] = l_cell_wire[33];							inform_L[33][2] = l_cell_wire[34];							inform_L[37][2] = l_cell_wire[35];							inform_L[34][2] = l_cell_wire[36];							inform_L[38][2] = l_cell_wire[37];							inform_L[35][2] = l_cell_wire[38];							inform_L[39][2] = l_cell_wire[39];							inform_L[40][2] = l_cell_wire[40];							inform_L[44][2] = l_cell_wire[41];							inform_L[41][2] = l_cell_wire[42];							inform_L[45][2] = l_cell_wire[43];							inform_L[42][2] = l_cell_wire[44];							inform_L[46][2] = l_cell_wire[45];							inform_L[43][2] = l_cell_wire[46];							inform_L[47][2] = l_cell_wire[47];							inform_L[48][2] = l_cell_wire[48];							inform_L[52][2] = l_cell_wire[49];							inform_L[49][2] = l_cell_wire[50];							inform_L[53][2] = l_cell_wire[51];							inform_L[50][2] = l_cell_wire[52];							inform_L[54][2] = l_cell_wire[53];							inform_L[51][2] = l_cell_wire[54];							inform_L[55][2] = l_cell_wire[55];							inform_L[56][2] = l_cell_wire[56];							inform_L[60][2] = l_cell_wire[57];							inform_L[57][2] = l_cell_wire[58];							inform_L[61][2] = l_cell_wire[59];							inform_L[58][2] = l_cell_wire[60];							inform_L[62][2] = l_cell_wire[61];							inform_L[59][2] = l_cell_wire[62];							inform_L[63][2] = l_cell_wire[63];							inform_L[64][2] = l_cell_wire[64];							inform_L[68][2] = l_cell_wire[65];							inform_L[65][2] = l_cell_wire[66];							inform_L[69][2] = l_cell_wire[67];							inform_L[66][2] = l_cell_wire[68];							inform_L[70][2] = l_cell_wire[69];							inform_L[67][2] = l_cell_wire[70];							inform_L[71][2] = l_cell_wire[71];							inform_L[72][2] = l_cell_wire[72];							inform_L[76][2] = l_cell_wire[73];							inform_L[73][2] = l_cell_wire[74];							inform_L[77][2] = l_cell_wire[75];							inform_L[74][2] = l_cell_wire[76];							inform_L[78][2] = l_cell_wire[77];							inform_L[75][2] = l_cell_wire[78];							inform_L[79][2] = l_cell_wire[79];							inform_L[80][2] = l_cell_wire[80];							inform_L[84][2] = l_cell_wire[81];							inform_L[81][2] = l_cell_wire[82];							inform_L[85][2] = l_cell_wire[83];							inform_L[82][2] = l_cell_wire[84];							inform_L[86][2] = l_cell_wire[85];							inform_L[83][2] = l_cell_wire[86];							inform_L[87][2] = l_cell_wire[87];							inform_L[88][2] = l_cell_wire[88];							inform_L[92][2] = l_cell_wire[89];							inform_L[89][2] = l_cell_wire[90];							inform_L[93][2] = l_cell_wire[91];							inform_L[90][2] = l_cell_wire[92];							inform_L[94][2] = l_cell_wire[93];							inform_L[91][2] = l_cell_wire[94];							inform_L[95][2] = l_cell_wire[95];							inform_L[96][2] = l_cell_wire[96];							inform_L[100][2] = l_cell_wire[97];							inform_L[97][2] = l_cell_wire[98];							inform_L[101][2] = l_cell_wire[99];							inform_L[98][2] = l_cell_wire[100];							inform_L[102][2] = l_cell_wire[101];							inform_L[99][2] = l_cell_wire[102];							inform_L[103][2] = l_cell_wire[103];							inform_L[104][2] = l_cell_wire[104];							inform_L[108][2] = l_cell_wire[105];							inform_L[105][2] = l_cell_wire[106];							inform_L[109][2] = l_cell_wire[107];							inform_L[106][2] = l_cell_wire[108];							inform_L[110][2] = l_cell_wire[109];							inform_L[107][2] = l_cell_wire[110];							inform_L[111][2] = l_cell_wire[111];							inform_L[112][2] = l_cell_wire[112];							inform_L[116][2] = l_cell_wire[113];							inform_L[113][2] = l_cell_wire[114];							inform_L[117][2] = l_cell_wire[115];							inform_L[114][2] = l_cell_wire[116];							inform_L[118][2] = l_cell_wire[117];							inform_L[115][2] = l_cell_wire[118];							inform_L[119][2] = l_cell_wire[119];							inform_L[120][2] = l_cell_wire[120];							inform_L[124][2] = l_cell_wire[121];							inform_L[121][2] = l_cell_wire[122];							inform_L[125][2] = l_cell_wire[123];							inform_L[122][2] = l_cell_wire[124];							inform_L[126][2] = l_cell_wire[125];							inform_L[123][2] = l_cell_wire[126];							inform_L[127][2] = l_cell_wire[127];							inform_L[128][2] = l_cell_wire[128];							inform_L[132][2] = l_cell_wire[129];							inform_L[129][2] = l_cell_wire[130];							inform_L[133][2] = l_cell_wire[131];							inform_L[130][2] = l_cell_wire[132];							inform_L[134][2] = l_cell_wire[133];							inform_L[131][2] = l_cell_wire[134];							inform_L[135][2] = l_cell_wire[135];							inform_L[136][2] = l_cell_wire[136];							inform_L[140][2] = l_cell_wire[137];							inform_L[137][2] = l_cell_wire[138];							inform_L[141][2] = l_cell_wire[139];							inform_L[138][2] = l_cell_wire[140];							inform_L[142][2] = l_cell_wire[141];							inform_L[139][2] = l_cell_wire[142];							inform_L[143][2] = l_cell_wire[143];							inform_L[144][2] = l_cell_wire[144];							inform_L[148][2] = l_cell_wire[145];							inform_L[145][2] = l_cell_wire[146];							inform_L[149][2] = l_cell_wire[147];							inform_L[146][2] = l_cell_wire[148];							inform_L[150][2] = l_cell_wire[149];							inform_L[147][2] = l_cell_wire[150];							inform_L[151][2] = l_cell_wire[151];							inform_L[152][2] = l_cell_wire[152];							inform_L[156][2] = l_cell_wire[153];							inform_L[153][2] = l_cell_wire[154];							inform_L[157][2] = l_cell_wire[155];							inform_L[154][2] = l_cell_wire[156];							inform_L[158][2] = l_cell_wire[157];							inform_L[155][2] = l_cell_wire[158];							inform_L[159][2] = l_cell_wire[159];							inform_L[160][2] = l_cell_wire[160];							inform_L[164][2] = l_cell_wire[161];							inform_L[161][2] = l_cell_wire[162];							inform_L[165][2] = l_cell_wire[163];							inform_L[162][2] = l_cell_wire[164];							inform_L[166][2] = l_cell_wire[165];							inform_L[163][2] = l_cell_wire[166];							inform_L[167][2] = l_cell_wire[167];							inform_L[168][2] = l_cell_wire[168];							inform_L[172][2] = l_cell_wire[169];							inform_L[169][2] = l_cell_wire[170];							inform_L[173][2] = l_cell_wire[171];							inform_L[170][2] = l_cell_wire[172];							inform_L[174][2] = l_cell_wire[173];							inform_L[171][2] = l_cell_wire[174];							inform_L[175][2] = l_cell_wire[175];							inform_L[176][2] = l_cell_wire[176];							inform_L[180][2] = l_cell_wire[177];							inform_L[177][2] = l_cell_wire[178];							inform_L[181][2] = l_cell_wire[179];							inform_L[178][2] = l_cell_wire[180];							inform_L[182][2] = l_cell_wire[181];							inform_L[179][2] = l_cell_wire[182];							inform_L[183][2] = l_cell_wire[183];							inform_L[184][2] = l_cell_wire[184];							inform_L[188][2] = l_cell_wire[185];							inform_L[185][2] = l_cell_wire[186];							inform_L[189][2] = l_cell_wire[187];							inform_L[186][2] = l_cell_wire[188];							inform_L[190][2] = l_cell_wire[189];							inform_L[187][2] = l_cell_wire[190];							inform_L[191][2] = l_cell_wire[191];							inform_L[192][2] = l_cell_wire[192];							inform_L[196][2] = l_cell_wire[193];							inform_L[193][2] = l_cell_wire[194];							inform_L[197][2] = l_cell_wire[195];							inform_L[194][2] = l_cell_wire[196];							inform_L[198][2] = l_cell_wire[197];							inform_L[195][2] = l_cell_wire[198];							inform_L[199][2] = l_cell_wire[199];							inform_L[200][2] = l_cell_wire[200];							inform_L[204][2] = l_cell_wire[201];							inform_L[201][2] = l_cell_wire[202];							inform_L[205][2] = l_cell_wire[203];							inform_L[202][2] = l_cell_wire[204];							inform_L[206][2] = l_cell_wire[205];							inform_L[203][2] = l_cell_wire[206];							inform_L[207][2] = l_cell_wire[207];							inform_L[208][2] = l_cell_wire[208];							inform_L[212][2] = l_cell_wire[209];							inform_L[209][2] = l_cell_wire[210];							inform_L[213][2] = l_cell_wire[211];							inform_L[210][2] = l_cell_wire[212];							inform_L[214][2] = l_cell_wire[213];							inform_L[211][2] = l_cell_wire[214];							inform_L[215][2] = l_cell_wire[215];							inform_L[216][2] = l_cell_wire[216];							inform_L[220][2] = l_cell_wire[217];							inform_L[217][2] = l_cell_wire[218];							inform_L[221][2] = l_cell_wire[219];							inform_L[218][2] = l_cell_wire[220];							inform_L[222][2] = l_cell_wire[221];							inform_L[219][2] = l_cell_wire[222];							inform_L[223][2] = l_cell_wire[223];							inform_L[224][2] = l_cell_wire[224];							inform_L[228][2] = l_cell_wire[225];							inform_L[225][2] = l_cell_wire[226];							inform_L[229][2] = l_cell_wire[227];							inform_L[226][2] = l_cell_wire[228];							inform_L[230][2] = l_cell_wire[229];							inform_L[227][2] = l_cell_wire[230];							inform_L[231][2] = l_cell_wire[231];							inform_L[232][2] = l_cell_wire[232];							inform_L[236][2] = l_cell_wire[233];							inform_L[233][2] = l_cell_wire[234];							inform_L[237][2] = l_cell_wire[235];							inform_L[234][2] = l_cell_wire[236];							inform_L[238][2] = l_cell_wire[237];							inform_L[235][2] = l_cell_wire[238];							inform_L[239][2] = l_cell_wire[239];							inform_L[240][2] = l_cell_wire[240];							inform_L[244][2] = l_cell_wire[241];							inform_L[241][2] = l_cell_wire[242];							inform_L[245][2] = l_cell_wire[243];							inform_L[242][2] = l_cell_wire[244];							inform_L[246][2] = l_cell_wire[245];							inform_L[243][2] = l_cell_wire[246];							inform_L[247][2] = l_cell_wire[247];							inform_L[248][2] = l_cell_wire[248];							inform_L[252][2] = l_cell_wire[249];							inform_L[249][2] = l_cell_wire[250];							inform_L[253][2] = l_cell_wire[251];							inform_L[250][2] = l_cell_wire[252];							inform_L[254][2] = l_cell_wire[253];							inform_L[251][2] = l_cell_wire[254];							inform_L[255][2] = l_cell_wire[255];						end
						4:						begin							inform_R[0][4] = r_cell_wire[0];							inform_R[8][4] = r_cell_wire[1];							inform_R[1][4] = r_cell_wire[2];							inform_R[9][4] = r_cell_wire[3];							inform_R[2][4] = r_cell_wire[4];							inform_R[10][4] = r_cell_wire[5];							inform_R[3][4] = r_cell_wire[6];							inform_R[11][4] = r_cell_wire[7];							inform_R[4][4] = r_cell_wire[8];							inform_R[12][4] = r_cell_wire[9];							inform_R[5][4] = r_cell_wire[10];							inform_R[13][4] = r_cell_wire[11];							inform_R[6][4] = r_cell_wire[12];							inform_R[14][4] = r_cell_wire[13];							inform_R[7][4] = r_cell_wire[14];							inform_R[15][4] = r_cell_wire[15];							inform_R[16][4] = r_cell_wire[16];							inform_R[24][4] = r_cell_wire[17];							inform_R[17][4] = r_cell_wire[18];							inform_R[25][4] = r_cell_wire[19];							inform_R[18][4] = r_cell_wire[20];							inform_R[26][4] = r_cell_wire[21];							inform_R[19][4] = r_cell_wire[22];							inform_R[27][4] = r_cell_wire[23];							inform_R[20][4] = r_cell_wire[24];							inform_R[28][4] = r_cell_wire[25];							inform_R[21][4] = r_cell_wire[26];							inform_R[29][4] = r_cell_wire[27];							inform_R[22][4] = r_cell_wire[28];							inform_R[30][4] = r_cell_wire[29];							inform_R[23][4] = r_cell_wire[30];							inform_R[31][4] = r_cell_wire[31];							inform_R[32][4] = r_cell_wire[32];							inform_R[40][4] = r_cell_wire[33];							inform_R[33][4] = r_cell_wire[34];							inform_R[41][4] = r_cell_wire[35];							inform_R[34][4] = r_cell_wire[36];							inform_R[42][4] = r_cell_wire[37];							inform_R[35][4] = r_cell_wire[38];							inform_R[43][4] = r_cell_wire[39];							inform_R[36][4] = r_cell_wire[40];							inform_R[44][4] = r_cell_wire[41];							inform_R[37][4] = r_cell_wire[42];							inform_R[45][4] = r_cell_wire[43];							inform_R[38][4] = r_cell_wire[44];							inform_R[46][4] = r_cell_wire[45];							inform_R[39][4] = r_cell_wire[46];							inform_R[47][4] = r_cell_wire[47];							inform_R[48][4] = r_cell_wire[48];							inform_R[56][4] = r_cell_wire[49];							inform_R[49][4] = r_cell_wire[50];							inform_R[57][4] = r_cell_wire[51];							inform_R[50][4] = r_cell_wire[52];							inform_R[58][4] = r_cell_wire[53];							inform_R[51][4] = r_cell_wire[54];							inform_R[59][4] = r_cell_wire[55];							inform_R[52][4] = r_cell_wire[56];							inform_R[60][4] = r_cell_wire[57];							inform_R[53][4] = r_cell_wire[58];							inform_R[61][4] = r_cell_wire[59];							inform_R[54][4] = r_cell_wire[60];							inform_R[62][4] = r_cell_wire[61];							inform_R[55][4] = r_cell_wire[62];							inform_R[63][4] = r_cell_wire[63];							inform_R[64][4] = r_cell_wire[64];							inform_R[72][4] = r_cell_wire[65];							inform_R[65][4] = r_cell_wire[66];							inform_R[73][4] = r_cell_wire[67];							inform_R[66][4] = r_cell_wire[68];							inform_R[74][4] = r_cell_wire[69];							inform_R[67][4] = r_cell_wire[70];							inform_R[75][4] = r_cell_wire[71];							inform_R[68][4] = r_cell_wire[72];							inform_R[76][4] = r_cell_wire[73];							inform_R[69][4] = r_cell_wire[74];							inform_R[77][4] = r_cell_wire[75];							inform_R[70][4] = r_cell_wire[76];							inform_R[78][4] = r_cell_wire[77];							inform_R[71][4] = r_cell_wire[78];							inform_R[79][4] = r_cell_wire[79];							inform_R[80][4] = r_cell_wire[80];							inform_R[88][4] = r_cell_wire[81];							inform_R[81][4] = r_cell_wire[82];							inform_R[89][4] = r_cell_wire[83];							inform_R[82][4] = r_cell_wire[84];							inform_R[90][4] = r_cell_wire[85];							inform_R[83][4] = r_cell_wire[86];							inform_R[91][4] = r_cell_wire[87];							inform_R[84][4] = r_cell_wire[88];							inform_R[92][4] = r_cell_wire[89];							inform_R[85][4] = r_cell_wire[90];							inform_R[93][4] = r_cell_wire[91];							inform_R[86][4] = r_cell_wire[92];							inform_R[94][4] = r_cell_wire[93];							inform_R[87][4] = r_cell_wire[94];							inform_R[95][4] = r_cell_wire[95];							inform_R[96][4] = r_cell_wire[96];							inform_R[104][4] = r_cell_wire[97];							inform_R[97][4] = r_cell_wire[98];							inform_R[105][4] = r_cell_wire[99];							inform_R[98][4] = r_cell_wire[100];							inform_R[106][4] = r_cell_wire[101];							inform_R[99][4] = r_cell_wire[102];							inform_R[107][4] = r_cell_wire[103];							inform_R[100][4] = r_cell_wire[104];							inform_R[108][4] = r_cell_wire[105];							inform_R[101][4] = r_cell_wire[106];							inform_R[109][4] = r_cell_wire[107];							inform_R[102][4] = r_cell_wire[108];							inform_R[110][4] = r_cell_wire[109];							inform_R[103][4] = r_cell_wire[110];							inform_R[111][4] = r_cell_wire[111];							inform_R[112][4] = r_cell_wire[112];							inform_R[120][4] = r_cell_wire[113];							inform_R[113][4] = r_cell_wire[114];							inform_R[121][4] = r_cell_wire[115];							inform_R[114][4] = r_cell_wire[116];							inform_R[122][4] = r_cell_wire[117];							inform_R[115][4] = r_cell_wire[118];							inform_R[123][4] = r_cell_wire[119];							inform_R[116][4] = r_cell_wire[120];							inform_R[124][4] = r_cell_wire[121];							inform_R[117][4] = r_cell_wire[122];							inform_R[125][4] = r_cell_wire[123];							inform_R[118][4] = r_cell_wire[124];							inform_R[126][4] = r_cell_wire[125];							inform_R[119][4] = r_cell_wire[126];							inform_R[127][4] = r_cell_wire[127];							inform_R[128][4] = r_cell_wire[128];							inform_R[136][4] = r_cell_wire[129];							inform_R[129][4] = r_cell_wire[130];							inform_R[137][4] = r_cell_wire[131];							inform_R[130][4] = r_cell_wire[132];							inform_R[138][4] = r_cell_wire[133];							inform_R[131][4] = r_cell_wire[134];							inform_R[139][4] = r_cell_wire[135];							inform_R[132][4] = r_cell_wire[136];							inform_R[140][4] = r_cell_wire[137];							inform_R[133][4] = r_cell_wire[138];							inform_R[141][4] = r_cell_wire[139];							inform_R[134][4] = r_cell_wire[140];							inform_R[142][4] = r_cell_wire[141];							inform_R[135][4] = r_cell_wire[142];							inform_R[143][4] = r_cell_wire[143];							inform_R[144][4] = r_cell_wire[144];							inform_R[152][4] = r_cell_wire[145];							inform_R[145][4] = r_cell_wire[146];							inform_R[153][4] = r_cell_wire[147];							inform_R[146][4] = r_cell_wire[148];							inform_R[154][4] = r_cell_wire[149];							inform_R[147][4] = r_cell_wire[150];							inform_R[155][4] = r_cell_wire[151];							inform_R[148][4] = r_cell_wire[152];							inform_R[156][4] = r_cell_wire[153];							inform_R[149][4] = r_cell_wire[154];							inform_R[157][4] = r_cell_wire[155];							inform_R[150][4] = r_cell_wire[156];							inform_R[158][4] = r_cell_wire[157];							inform_R[151][4] = r_cell_wire[158];							inform_R[159][4] = r_cell_wire[159];							inform_R[160][4] = r_cell_wire[160];							inform_R[168][4] = r_cell_wire[161];							inform_R[161][4] = r_cell_wire[162];							inform_R[169][4] = r_cell_wire[163];							inform_R[162][4] = r_cell_wire[164];							inform_R[170][4] = r_cell_wire[165];							inform_R[163][4] = r_cell_wire[166];							inform_R[171][4] = r_cell_wire[167];							inform_R[164][4] = r_cell_wire[168];							inform_R[172][4] = r_cell_wire[169];							inform_R[165][4] = r_cell_wire[170];							inform_R[173][4] = r_cell_wire[171];							inform_R[166][4] = r_cell_wire[172];							inform_R[174][4] = r_cell_wire[173];							inform_R[167][4] = r_cell_wire[174];							inform_R[175][4] = r_cell_wire[175];							inform_R[176][4] = r_cell_wire[176];							inform_R[184][4] = r_cell_wire[177];							inform_R[177][4] = r_cell_wire[178];							inform_R[185][4] = r_cell_wire[179];							inform_R[178][4] = r_cell_wire[180];							inform_R[186][4] = r_cell_wire[181];							inform_R[179][4] = r_cell_wire[182];							inform_R[187][4] = r_cell_wire[183];							inform_R[180][4] = r_cell_wire[184];							inform_R[188][4] = r_cell_wire[185];							inform_R[181][4] = r_cell_wire[186];							inform_R[189][4] = r_cell_wire[187];							inform_R[182][4] = r_cell_wire[188];							inform_R[190][4] = r_cell_wire[189];							inform_R[183][4] = r_cell_wire[190];							inform_R[191][4] = r_cell_wire[191];							inform_R[192][4] = r_cell_wire[192];							inform_R[200][4] = r_cell_wire[193];							inform_R[193][4] = r_cell_wire[194];							inform_R[201][4] = r_cell_wire[195];							inform_R[194][4] = r_cell_wire[196];							inform_R[202][4] = r_cell_wire[197];							inform_R[195][4] = r_cell_wire[198];							inform_R[203][4] = r_cell_wire[199];							inform_R[196][4] = r_cell_wire[200];							inform_R[204][4] = r_cell_wire[201];							inform_R[197][4] = r_cell_wire[202];							inform_R[205][4] = r_cell_wire[203];							inform_R[198][4] = r_cell_wire[204];							inform_R[206][4] = r_cell_wire[205];							inform_R[199][4] = r_cell_wire[206];							inform_R[207][4] = r_cell_wire[207];							inform_R[208][4] = r_cell_wire[208];							inform_R[216][4] = r_cell_wire[209];							inform_R[209][4] = r_cell_wire[210];							inform_R[217][4] = r_cell_wire[211];							inform_R[210][4] = r_cell_wire[212];							inform_R[218][4] = r_cell_wire[213];							inform_R[211][4] = r_cell_wire[214];							inform_R[219][4] = r_cell_wire[215];							inform_R[212][4] = r_cell_wire[216];							inform_R[220][4] = r_cell_wire[217];							inform_R[213][4] = r_cell_wire[218];							inform_R[221][4] = r_cell_wire[219];							inform_R[214][4] = r_cell_wire[220];							inform_R[222][4] = r_cell_wire[221];							inform_R[215][4] = r_cell_wire[222];							inform_R[223][4] = r_cell_wire[223];							inform_R[224][4] = r_cell_wire[224];							inform_R[232][4] = r_cell_wire[225];							inform_R[225][4] = r_cell_wire[226];							inform_R[233][4] = r_cell_wire[227];							inform_R[226][4] = r_cell_wire[228];							inform_R[234][4] = r_cell_wire[229];							inform_R[227][4] = r_cell_wire[230];							inform_R[235][4] = r_cell_wire[231];							inform_R[228][4] = r_cell_wire[232];							inform_R[236][4] = r_cell_wire[233];							inform_R[229][4] = r_cell_wire[234];							inform_R[237][4] = r_cell_wire[235];							inform_R[230][4] = r_cell_wire[236];							inform_R[238][4] = r_cell_wire[237];							inform_R[231][4] = r_cell_wire[238];							inform_R[239][4] = r_cell_wire[239];							inform_R[240][4] = r_cell_wire[240];							inform_R[248][4] = r_cell_wire[241];							inform_R[241][4] = r_cell_wire[242];							inform_R[249][4] = r_cell_wire[243];							inform_R[242][4] = r_cell_wire[244];							inform_R[250][4] = r_cell_wire[245];							inform_R[243][4] = r_cell_wire[246];							inform_R[251][4] = r_cell_wire[247];							inform_R[244][4] = r_cell_wire[248];							inform_R[252][4] = r_cell_wire[249];							inform_R[245][4] = r_cell_wire[250];							inform_R[253][4] = r_cell_wire[251];							inform_R[246][4] = r_cell_wire[252];							inform_R[254][4] = r_cell_wire[253];							inform_R[247][4] = r_cell_wire[254];							inform_R[255][4] = r_cell_wire[255];							inform_L[0][3] = l_cell_wire[0];							inform_L[8][3] = l_cell_wire[1];							inform_L[1][3] = l_cell_wire[2];							inform_L[9][3] = l_cell_wire[3];							inform_L[2][3] = l_cell_wire[4];							inform_L[10][3] = l_cell_wire[5];							inform_L[3][3] = l_cell_wire[6];							inform_L[11][3] = l_cell_wire[7];							inform_L[4][3] = l_cell_wire[8];							inform_L[12][3] = l_cell_wire[9];							inform_L[5][3] = l_cell_wire[10];							inform_L[13][3] = l_cell_wire[11];							inform_L[6][3] = l_cell_wire[12];							inform_L[14][3] = l_cell_wire[13];							inform_L[7][3] = l_cell_wire[14];							inform_L[15][3] = l_cell_wire[15];							inform_L[16][3] = l_cell_wire[16];							inform_L[24][3] = l_cell_wire[17];							inform_L[17][3] = l_cell_wire[18];							inform_L[25][3] = l_cell_wire[19];							inform_L[18][3] = l_cell_wire[20];							inform_L[26][3] = l_cell_wire[21];							inform_L[19][3] = l_cell_wire[22];							inform_L[27][3] = l_cell_wire[23];							inform_L[20][3] = l_cell_wire[24];							inform_L[28][3] = l_cell_wire[25];							inform_L[21][3] = l_cell_wire[26];							inform_L[29][3] = l_cell_wire[27];							inform_L[22][3] = l_cell_wire[28];							inform_L[30][3] = l_cell_wire[29];							inform_L[23][3] = l_cell_wire[30];							inform_L[31][3] = l_cell_wire[31];							inform_L[32][3] = l_cell_wire[32];							inform_L[40][3] = l_cell_wire[33];							inform_L[33][3] = l_cell_wire[34];							inform_L[41][3] = l_cell_wire[35];							inform_L[34][3] = l_cell_wire[36];							inform_L[42][3] = l_cell_wire[37];							inform_L[35][3] = l_cell_wire[38];							inform_L[43][3] = l_cell_wire[39];							inform_L[36][3] = l_cell_wire[40];							inform_L[44][3] = l_cell_wire[41];							inform_L[37][3] = l_cell_wire[42];							inform_L[45][3] = l_cell_wire[43];							inform_L[38][3] = l_cell_wire[44];							inform_L[46][3] = l_cell_wire[45];							inform_L[39][3] = l_cell_wire[46];							inform_L[47][3] = l_cell_wire[47];							inform_L[48][3] = l_cell_wire[48];							inform_L[56][3] = l_cell_wire[49];							inform_L[49][3] = l_cell_wire[50];							inform_L[57][3] = l_cell_wire[51];							inform_L[50][3] = l_cell_wire[52];							inform_L[58][3] = l_cell_wire[53];							inform_L[51][3] = l_cell_wire[54];							inform_L[59][3] = l_cell_wire[55];							inform_L[52][3] = l_cell_wire[56];							inform_L[60][3] = l_cell_wire[57];							inform_L[53][3] = l_cell_wire[58];							inform_L[61][3] = l_cell_wire[59];							inform_L[54][3] = l_cell_wire[60];							inform_L[62][3] = l_cell_wire[61];							inform_L[55][3] = l_cell_wire[62];							inform_L[63][3] = l_cell_wire[63];							inform_L[64][3] = l_cell_wire[64];							inform_L[72][3] = l_cell_wire[65];							inform_L[65][3] = l_cell_wire[66];							inform_L[73][3] = l_cell_wire[67];							inform_L[66][3] = l_cell_wire[68];							inform_L[74][3] = l_cell_wire[69];							inform_L[67][3] = l_cell_wire[70];							inform_L[75][3] = l_cell_wire[71];							inform_L[68][3] = l_cell_wire[72];							inform_L[76][3] = l_cell_wire[73];							inform_L[69][3] = l_cell_wire[74];							inform_L[77][3] = l_cell_wire[75];							inform_L[70][3] = l_cell_wire[76];							inform_L[78][3] = l_cell_wire[77];							inform_L[71][3] = l_cell_wire[78];							inform_L[79][3] = l_cell_wire[79];							inform_L[80][3] = l_cell_wire[80];							inform_L[88][3] = l_cell_wire[81];							inform_L[81][3] = l_cell_wire[82];							inform_L[89][3] = l_cell_wire[83];							inform_L[82][3] = l_cell_wire[84];							inform_L[90][3] = l_cell_wire[85];							inform_L[83][3] = l_cell_wire[86];							inform_L[91][3] = l_cell_wire[87];							inform_L[84][3] = l_cell_wire[88];							inform_L[92][3] = l_cell_wire[89];							inform_L[85][3] = l_cell_wire[90];							inform_L[93][3] = l_cell_wire[91];							inform_L[86][3] = l_cell_wire[92];							inform_L[94][3] = l_cell_wire[93];							inform_L[87][3] = l_cell_wire[94];							inform_L[95][3] = l_cell_wire[95];							inform_L[96][3] = l_cell_wire[96];							inform_L[104][3] = l_cell_wire[97];							inform_L[97][3] = l_cell_wire[98];							inform_L[105][3] = l_cell_wire[99];							inform_L[98][3] = l_cell_wire[100];							inform_L[106][3] = l_cell_wire[101];							inform_L[99][3] = l_cell_wire[102];							inform_L[107][3] = l_cell_wire[103];							inform_L[100][3] = l_cell_wire[104];							inform_L[108][3] = l_cell_wire[105];							inform_L[101][3] = l_cell_wire[106];							inform_L[109][3] = l_cell_wire[107];							inform_L[102][3] = l_cell_wire[108];							inform_L[110][3] = l_cell_wire[109];							inform_L[103][3] = l_cell_wire[110];							inform_L[111][3] = l_cell_wire[111];							inform_L[112][3] = l_cell_wire[112];							inform_L[120][3] = l_cell_wire[113];							inform_L[113][3] = l_cell_wire[114];							inform_L[121][3] = l_cell_wire[115];							inform_L[114][3] = l_cell_wire[116];							inform_L[122][3] = l_cell_wire[117];							inform_L[115][3] = l_cell_wire[118];							inform_L[123][3] = l_cell_wire[119];							inform_L[116][3] = l_cell_wire[120];							inform_L[124][3] = l_cell_wire[121];							inform_L[117][3] = l_cell_wire[122];							inform_L[125][3] = l_cell_wire[123];							inform_L[118][3] = l_cell_wire[124];							inform_L[126][3] = l_cell_wire[125];							inform_L[119][3] = l_cell_wire[126];							inform_L[127][3] = l_cell_wire[127];							inform_L[128][3] = l_cell_wire[128];							inform_L[136][3] = l_cell_wire[129];							inform_L[129][3] = l_cell_wire[130];							inform_L[137][3] = l_cell_wire[131];							inform_L[130][3] = l_cell_wire[132];							inform_L[138][3] = l_cell_wire[133];							inform_L[131][3] = l_cell_wire[134];							inform_L[139][3] = l_cell_wire[135];							inform_L[132][3] = l_cell_wire[136];							inform_L[140][3] = l_cell_wire[137];							inform_L[133][3] = l_cell_wire[138];							inform_L[141][3] = l_cell_wire[139];							inform_L[134][3] = l_cell_wire[140];							inform_L[142][3] = l_cell_wire[141];							inform_L[135][3] = l_cell_wire[142];							inform_L[143][3] = l_cell_wire[143];							inform_L[144][3] = l_cell_wire[144];							inform_L[152][3] = l_cell_wire[145];							inform_L[145][3] = l_cell_wire[146];							inform_L[153][3] = l_cell_wire[147];							inform_L[146][3] = l_cell_wire[148];							inform_L[154][3] = l_cell_wire[149];							inform_L[147][3] = l_cell_wire[150];							inform_L[155][3] = l_cell_wire[151];							inform_L[148][3] = l_cell_wire[152];							inform_L[156][3] = l_cell_wire[153];							inform_L[149][3] = l_cell_wire[154];							inform_L[157][3] = l_cell_wire[155];							inform_L[150][3] = l_cell_wire[156];							inform_L[158][3] = l_cell_wire[157];							inform_L[151][3] = l_cell_wire[158];							inform_L[159][3] = l_cell_wire[159];							inform_L[160][3] = l_cell_wire[160];							inform_L[168][3] = l_cell_wire[161];							inform_L[161][3] = l_cell_wire[162];							inform_L[169][3] = l_cell_wire[163];							inform_L[162][3] = l_cell_wire[164];							inform_L[170][3] = l_cell_wire[165];							inform_L[163][3] = l_cell_wire[166];							inform_L[171][3] = l_cell_wire[167];							inform_L[164][3] = l_cell_wire[168];							inform_L[172][3] = l_cell_wire[169];							inform_L[165][3] = l_cell_wire[170];							inform_L[173][3] = l_cell_wire[171];							inform_L[166][3] = l_cell_wire[172];							inform_L[174][3] = l_cell_wire[173];							inform_L[167][3] = l_cell_wire[174];							inform_L[175][3] = l_cell_wire[175];							inform_L[176][3] = l_cell_wire[176];							inform_L[184][3] = l_cell_wire[177];							inform_L[177][3] = l_cell_wire[178];							inform_L[185][3] = l_cell_wire[179];							inform_L[178][3] = l_cell_wire[180];							inform_L[186][3] = l_cell_wire[181];							inform_L[179][3] = l_cell_wire[182];							inform_L[187][3] = l_cell_wire[183];							inform_L[180][3] = l_cell_wire[184];							inform_L[188][3] = l_cell_wire[185];							inform_L[181][3] = l_cell_wire[186];							inform_L[189][3] = l_cell_wire[187];							inform_L[182][3] = l_cell_wire[188];							inform_L[190][3] = l_cell_wire[189];							inform_L[183][3] = l_cell_wire[190];							inform_L[191][3] = l_cell_wire[191];							inform_L[192][3] = l_cell_wire[192];							inform_L[200][3] = l_cell_wire[193];							inform_L[193][3] = l_cell_wire[194];							inform_L[201][3] = l_cell_wire[195];							inform_L[194][3] = l_cell_wire[196];							inform_L[202][3] = l_cell_wire[197];							inform_L[195][3] = l_cell_wire[198];							inform_L[203][3] = l_cell_wire[199];							inform_L[196][3] = l_cell_wire[200];							inform_L[204][3] = l_cell_wire[201];							inform_L[197][3] = l_cell_wire[202];							inform_L[205][3] = l_cell_wire[203];							inform_L[198][3] = l_cell_wire[204];							inform_L[206][3] = l_cell_wire[205];							inform_L[199][3] = l_cell_wire[206];							inform_L[207][3] = l_cell_wire[207];							inform_L[208][3] = l_cell_wire[208];							inform_L[216][3] = l_cell_wire[209];							inform_L[209][3] = l_cell_wire[210];							inform_L[217][3] = l_cell_wire[211];							inform_L[210][3] = l_cell_wire[212];							inform_L[218][3] = l_cell_wire[213];							inform_L[211][3] = l_cell_wire[214];							inform_L[219][3] = l_cell_wire[215];							inform_L[212][3] = l_cell_wire[216];							inform_L[220][3] = l_cell_wire[217];							inform_L[213][3] = l_cell_wire[218];							inform_L[221][3] = l_cell_wire[219];							inform_L[214][3] = l_cell_wire[220];							inform_L[222][3] = l_cell_wire[221];							inform_L[215][3] = l_cell_wire[222];							inform_L[223][3] = l_cell_wire[223];							inform_L[224][3] = l_cell_wire[224];							inform_L[232][3] = l_cell_wire[225];							inform_L[225][3] = l_cell_wire[226];							inform_L[233][3] = l_cell_wire[227];							inform_L[226][3] = l_cell_wire[228];							inform_L[234][3] = l_cell_wire[229];							inform_L[227][3] = l_cell_wire[230];							inform_L[235][3] = l_cell_wire[231];							inform_L[228][3] = l_cell_wire[232];							inform_L[236][3] = l_cell_wire[233];							inform_L[229][3] = l_cell_wire[234];							inform_L[237][3] = l_cell_wire[235];							inform_L[230][3] = l_cell_wire[236];							inform_L[238][3] = l_cell_wire[237];							inform_L[231][3] = l_cell_wire[238];							inform_L[239][3] = l_cell_wire[239];							inform_L[240][3] = l_cell_wire[240];							inform_L[248][3] = l_cell_wire[241];							inform_L[241][3] = l_cell_wire[242];							inform_L[249][3] = l_cell_wire[243];							inform_L[242][3] = l_cell_wire[244];							inform_L[250][3] = l_cell_wire[245];							inform_L[243][3] = l_cell_wire[246];							inform_L[251][3] = l_cell_wire[247];							inform_L[244][3] = l_cell_wire[248];							inform_L[252][3] = l_cell_wire[249];							inform_L[245][3] = l_cell_wire[250];							inform_L[253][3] = l_cell_wire[251];							inform_L[246][3] = l_cell_wire[252];							inform_L[254][3] = l_cell_wire[253];							inform_L[247][3] = l_cell_wire[254];							inform_L[255][3] = l_cell_wire[255];						end
						5:						begin							inform_R[0][5] = r_cell_wire[0];							inform_R[16][5] = r_cell_wire[1];							inform_R[1][5] = r_cell_wire[2];							inform_R[17][5] = r_cell_wire[3];							inform_R[2][5] = r_cell_wire[4];							inform_R[18][5] = r_cell_wire[5];							inform_R[3][5] = r_cell_wire[6];							inform_R[19][5] = r_cell_wire[7];							inform_R[4][5] = r_cell_wire[8];							inform_R[20][5] = r_cell_wire[9];							inform_R[5][5] = r_cell_wire[10];							inform_R[21][5] = r_cell_wire[11];							inform_R[6][5] = r_cell_wire[12];							inform_R[22][5] = r_cell_wire[13];							inform_R[7][5] = r_cell_wire[14];							inform_R[23][5] = r_cell_wire[15];							inform_R[8][5] = r_cell_wire[16];							inform_R[24][5] = r_cell_wire[17];							inform_R[9][5] = r_cell_wire[18];							inform_R[25][5] = r_cell_wire[19];							inform_R[10][5] = r_cell_wire[20];							inform_R[26][5] = r_cell_wire[21];							inform_R[11][5] = r_cell_wire[22];							inform_R[27][5] = r_cell_wire[23];							inform_R[12][5] = r_cell_wire[24];							inform_R[28][5] = r_cell_wire[25];							inform_R[13][5] = r_cell_wire[26];							inform_R[29][5] = r_cell_wire[27];							inform_R[14][5] = r_cell_wire[28];							inform_R[30][5] = r_cell_wire[29];							inform_R[15][5] = r_cell_wire[30];							inform_R[31][5] = r_cell_wire[31];							inform_R[32][5] = r_cell_wire[32];							inform_R[48][5] = r_cell_wire[33];							inform_R[33][5] = r_cell_wire[34];							inform_R[49][5] = r_cell_wire[35];							inform_R[34][5] = r_cell_wire[36];							inform_R[50][5] = r_cell_wire[37];							inform_R[35][5] = r_cell_wire[38];							inform_R[51][5] = r_cell_wire[39];							inform_R[36][5] = r_cell_wire[40];							inform_R[52][5] = r_cell_wire[41];							inform_R[37][5] = r_cell_wire[42];							inform_R[53][5] = r_cell_wire[43];							inform_R[38][5] = r_cell_wire[44];							inform_R[54][5] = r_cell_wire[45];							inform_R[39][5] = r_cell_wire[46];							inform_R[55][5] = r_cell_wire[47];							inform_R[40][5] = r_cell_wire[48];							inform_R[56][5] = r_cell_wire[49];							inform_R[41][5] = r_cell_wire[50];							inform_R[57][5] = r_cell_wire[51];							inform_R[42][5] = r_cell_wire[52];							inform_R[58][5] = r_cell_wire[53];							inform_R[43][5] = r_cell_wire[54];							inform_R[59][5] = r_cell_wire[55];							inform_R[44][5] = r_cell_wire[56];							inform_R[60][5] = r_cell_wire[57];							inform_R[45][5] = r_cell_wire[58];							inform_R[61][5] = r_cell_wire[59];							inform_R[46][5] = r_cell_wire[60];							inform_R[62][5] = r_cell_wire[61];							inform_R[47][5] = r_cell_wire[62];							inform_R[63][5] = r_cell_wire[63];							inform_R[64][5] = r_cell_wire[64];							inform_R[80][5] = r_cell_wire[65];							inform_R[65][5] = r_cell_wire[66];							inform_R[81][5] = r_cell_wire[67];							inform_R[66][5] = r_cell_wire[68];							inform_R[82][5] = r_cell_wire[69];							inform_R[67][5] = r_cell_wire[70];							inform_R[83][5] = r_cell_wire[71];							inform_R[68][5] = r_cell_wire[72];							inform_R[84][5] = r_cell_wire[73];							inform_R[69][5] = r_cell_wire[74];							inform_R[85][5] = r_cell_wire[75];							inform_R[70][5] = r_cell_wire[76];							inform_R[86][5] = r_cell_wire[77];							inform_R[71][5] = r_cell_wire[78];							inform_R[87][5] = r_cell_wire[79];							inform_R[72][5] = r_cell_wire[80];							inform_R[88][5] = r_cell_wire[81];							inform_R[73][5] = r_cell_wire[82];							inform_R[89][5] = r_cell_wire[83];							inform_R[74][5] = r_cell_wire[84];							inform_R[90][5] = r_cell_wire[85];							inform_R[75][5] = r_cell_wire[86];							inform_R[91][5] = r_cell_wire[87];							inform_R[76][5] = r_cell_wire[88];							inform_R[92][5] = r_cell_wire[89];							inform_R[77][5] = r_cell_wire[90];							inform_R[93][5] = r_cell_wire[91];							inform_R[78][5] = r_cell_wire[92];							inform_R[94][5] = r_cell_wire[93];							inform_R[79][5] = r_cell_wire[94];							inform_R[95][5] = r_cell_wire[95];							inform_R[96][5] = r_cell_wire[96];							inform_R[112][5] = r_cell_wire[97];							inform_R[97][5] = r_cell_wire[98];							inform_R[113][5] = r_cell_wire[99];							inform_R[98][5] = r_cell_wire[100];							inform_R[114][5] = r_cell_wire[101];							inform_R[99][5] = r_cell_wire[102];							inform_R[115][5] = r_cell_wire[103];							inform_R[100][5] = r_cell_wire[104];							inform_R[116][5] = r_cell_wire[105];							inform_R[101][5] = r_cell_wire[106];							inform_R[117][5] = r_cell_wire[107];							inform_R[102][5] = r_cell_wire[108];							inform_R[118][5] = r_cell_wire[109];							inform_R[103][5] = r_cell_wire[110];							inform_R[119][5] = r_cell_wire[111];							inform_R[104][5] = r_cell_wire[112];							inform_R[120][5] = r_cell_wire[113];							inform_R[105][5] = r_cell_wire[114];							inform_R[121][5] = r_cell_wire[115];							inform_R[106][5] = r_cell_wire[116];							inform_R[122][5] = r_cell_wire[117];							inform_R[107][5] = r_cell_wire[118];							inform_R[123][5] = r_cell_wire[119];							inform_R[108][5] = r_cell_wire[120];							inform_R[124][5] = r_cell_wire[121];							inform_R[109][5] = r_cell_wire[122];							inform_R[125][5] = r_cell_wire[123];							inform_R[110][5] = r_cell_wire[124];							inform_R[126][5] = r_cell_wire[125];							inform_R[111][5] = r_cell_wire[126];							inform_R[127][5] = r_cell_wire[127];							inform_R[128][5] = r_cell_wire[128];							inform_R[144][5] = r_cell_wire[129];							inform_R[129][5] = r_cell_wire[130];							inform_R[145][5] = r_cell_wire[131];							inform_R[130][5] = r_cell_wire[132];							inform_R[146][5] = r_cell_wire[133];							inform_R[131][5] = r_cell_wire[134];							inform_R[147][5] = r_cell_wire[135];							inform_R[132][5] = r_cell_wire[136];							inform_R[148][5] = r_cell_wire[137];							inform_R[133][5] = r_cell_wire[138];							inform_R[149][5] = r_cell_wire[139];							inform_R[134][5] = r_cell_wire[140];							inform_R[150][5] = r_cell_wire[141];							inform_R[135][5] = r_cell_wire[142];							inform_R[151][5] = r_cell_wire[143];							inform_R[136][5] = r_cell_wire[144];							inform_R[152][5] = r_cell_wire[145];							inform_R[137][5] = r_cell_wire[146];							inform_R[153][5] = r_cell_wire[147];							inform_R[138][5] = r_cell_wire[148];							inform_R[154][5] = r_cell_wire[149];							inform_R[139][5] = r_cell_wire[150];							inform_R[155][5] = r_cell_wire[151];							inform_R[140][5] = r_cell_wire[152];							inform_R[156][5] = r_cell_wire[153];							inform_R[141][5] = r_cell_wire[154];							inform_R[157][5] = r_cell_wire[155];							inform_R[142][5] = r_cell_wire[156];							inform_R[158][5] = r_cell_wire[157];							inform_R[143][5] = r_cell_wire[158];							inform_R[159][5] = r_cell_wire[159];							inform_R[160][5] = r_cell_wire[160];							inform_R[176][5] = r_cell_wire[161];							inform_R[161][5] = r_cell_wire[162];							inform_R[177][5] = r_cell_wire[163];							inform_R[162][5] = r_cell_wire[164];							inform_R[178][5] = r_cell_wire[165];							inform_R[163][5] = r_cell_wire[166];							inform_R[179][5] = r_cell_wire[167];							inform_R[164][5] = r_cell_wire[168];							inform_R[180][5] = r_cell_wire[169];							inform_R[165][5] = r_cell_wire[170];							inform_R[181][5] = r_cell_wire[171];							inform_R[166][5] = r_cell_wire[172];							inform_R[182][5] = r_cell_wire[173];							inform_R[167][5] = r_cell_wire[174];							inform_R[183][5] = r_cell_wire[175];							inform_R[168][5] = r_cell_wire[176];							inform_R[184][5] = r_cell_wire[177];							inform_R[169][5] = r_cell_wire[178];							inform_R[185][5] = r_cell_wire[179];							inform_R[170][5] = r_cell_wire[180];							inform_R[186][5] = r_cell_wire[181];							inform_R[171][5] = r_cell_wire[182];							inform_R[187][5] = r_cell_wire[183];							inform_R[172][5] = r_cell_wire[184];							inform_R[188][5] = r_cell_wire[185];							inform_R[173][5] = r_cell_wire[186];							inform_R[189][5] = r_cell_wire[187];							inform_R[174][5] = r_cell_wire[188];							inform_R[190][5] = r_cell_wire[189];							inform_R[175][5] = r_cell_wire[190];							inform_R[191][5] = r_cell_wire[191];							inform_R[192][5] = r_cell_wire[192];							inform_R[208][5] = r_cell_wire[193];							inform_R[193][5] = r_cell_wire[194];							inform_R[209][5] = r_cell_wire[195];							inform_R[194][5] = r_cell_wire[196];							inform_R[210][5] = r_cell_wire[197];							inform_R[195][5] = r_cell_wire[198];							inform_R[211][5] = r_cell_wire[199];							inform_R[196][5] = r_cell_wire[200];							inform_R[212][5] = r_cell_wire[201];							inform_R[197][5] = r_cell_wire[202];							inform_R[213][5] = r_cell_wire[203];							inform_R[198][5] = r_cell_wire[204];							inform_R[214][5] = r_cell_wire[205];							inform_R[199][5] = r_cell_wire[206];							inform_R[215][5] = r_cell_wire[207];							inform_R[200][5] = r_cell_wire[208];							inform_R[216][5] = r_cell_wire[209];							inform_R[201][5] = r_cell_wire[210];							inform_R[217][5] = r_cell_wire[211];							inform_R[202][5] = r_cell_wire[212];							inform_R[218][5] = r_cell_wire[213];							inform_R[203][5] = r_cell_wire[214];							inform_R[219][5] = r_cell_wire[215];							inform_R[204][5] = r_cell_wire[216];							inform_R[220][5] = r_cell_wire[217];							inform_R[205][5] = r_cell_wire[218];							inform_R[221][5] = r_cell_wire[219];							inform_R[206][5] = r_cell_wire[220];							inform_R[222][5] = r_cell_wire[221];							inform_R[207][5] = r_cell_wire[222];							inform_R[223][5] = r_cell_wire[223];							inform_R[224][5] = r_cell_wire[224];							inform_R[240][5] = r_cell_wire[225];							inform_R[225][5] = r_cell_wire[226];							inform_R[241][5] = r_cell_wire[227];							inform_R[226][5] = r_cell_wire[228];							inform_R[242][5] = r_cell_wire[229];							inform_R[227][5] = r_cell_wire[230];							inform_R[243][5] = r_cell_wire[231];							inform_R[228][5] = r_cell_wire[232];							inform_R[244][5] = r_cell_wire[233];							inform_R[229][5] = r_cell_wire[234];							inform_R[245][5] = r_cell_wire[235];							inform_R[230][5] = r_cell_wire[236];							inform_R[246][5] = r_cell_wire[237];							inform_R[231][5] = r_cell_wire[238];							inform_R[247][5] = r_cell_wire[239];							inform_R[232][5] = r_cell_wire[240];							inform_R[248][5] = r_cell_wire[241];							inform_R[233][5] = r_cell_wire[242];							inform_R[249][5] = r_cell_wire[243];							inform_R[234][5] = r_cell_wire[244];							inform_R[250][5] = r_cell_wire[245];							inform_R[235][5] = r_cell_wire[246];							inform_R[251][5] = r_cell_wire[247];							inform_R[236][5] = r_cell_wire[248];							inform_R[252][5] = r_cell_wire[249];							inform_R[237][5] = r_cell_wire[250];							inform_R[253][5] = r_cell_wire[251];							inform_R[238][5] = r_cell_wire[252];							inform_R[254][5] = r_cell_wire[253];							inform_R[239][5] = r_cell_wire[254];							inform_R[255][5] = r_cell_wire[255];							inform_L[0][4] = l_cell_wire[0];							inform_L[16][4] = l_cell_wire[1];							inform_L[1][4] = l_cell_wire[2];							inform_L[17][4] = l_cell_wire[3];							inform_L[2][4] = l_cell_wire[4];							inform_L[18][4] = l_cell_wire[5];							inform_L[3][4] = l_cell_wire[6];							inform_L[19][4] = l_cell_wire[7];							inform_L[4][4] = l_cell_wire[8];							inform_L[20][4] = l_cell_wire[9];							inform_L[5][4] = l_cell_wire[10];							inform_L[21][4] = l_cell_wire[11];							inform_L[6][4] = l_cell_wire[12];							inform_L[22][4] = l_cell_wire[13];							inform_L[7][4] = l_cell_wire[14];							inform_L[23][4] = l_cell_wire[15];							inform_L[8][4] = l_cell_wire[16];							inform_L[24][4] = l_cell_wire[17];							inform_L[9][4] = l_cell_wire[18];							inform_L[25][4] = l_cell_wire[19];							inform_L[10][4] = l_cell_wire[20];							inform_L[26][4] = l_cell_wire[21];							inform_L[11][4] = l_cell_wire[22];							inform_L[27][4] = l_cell_wire[23];							inform_L[12][4] = l_cell_wire[24];							inform_L[28][4] = l_cell_wire[25];							inform_L[13][4] = l_cell_wire[26];							inform_L[29][4] = l_cell_wire[27];							inform_L[14][4] = l_cell_wire[28];							inform_L[30][4] = l_cell_wire[29];							inform_L[15][4] = l_cell_wire[30];							inform_L[31][4] = l_cell_wire[31];							inform_L[32][4] = l_cell_wire[32];							inform_L[48][4] = l_cell_wire[33];							inform_L[33][4] = l_cell_wire[34];							inform_L[49][4] = l_cell_wire[35];							inform_L[34][4] = l_cell_wire[36];							inform_L[50][4] = l_cell_wire[37];							inform_L[35][4] = l_cell_wire[38];							inform_L[51][4] = l_cell_wire[39];							inform_L[36][4] = l_cell_wire[40];							inform_L[52][4] = l_cell_wire[41];							inform_L[37][4] = l_cell_wire[42];							inform_L[53][4] = l_cell_wire[43];							inform_L[38][4] = l_cell_wire[44];							inform_L[54][4] = l_cell_wire[45];							inform_L[39][4] = l_cell_wire[46];							inform_L[55][4] = l_cell_wire[47];							inform_L[40][4] = l_cell_wire[48];							inform_L[56][4] = l_cell_wire[49];							inform_L[41][4] = l_cell_wire[50];							inform_L[57][4] = l_cell_wire[51];							inform_L[42][4] = l_cell_wire[52];							inform_L[58][4] = l_cell_wire[53];							inform_L[43][4] = l_cell_wire[54];							inform_L[59][4] = l_cell_wire[55];							inform_L[44][4] = l_cell_wire[56];							inform_L[60][4] = l_cell_wire[57];							inform_L[45][4] = l_cell_wire[58];							inform_L[61][4] = l_cell_wire[59];							inform_L[46][4] = l_cell_wire[60];							inform_L[62][4] = l_cell_wire[61];							inform_L[47][4] = l_cell_wire[62];							inform_L[63][4] = l_cell_wire[63];							inform_L[64][4] = l_cell_wire[64];							inform_L[80][4] = l_cell_wire[65];							inform_L[65][4] = l_cell_wire[66];							inform_L[81][4] = l_cell_wire[67];							inform_L[66][4] = l_cell_wire[68];							inform_L[82][4] = l_cell_wire[69];							inform_L[67][4] = l_cell_wire[70];							inform_L[83][4] = l_cell_wire[71];							inform_L[68][4] = l_cell_wire[72];							inform_L[84][4] = l_cell_wire[73];							inform_L[69][4] = l_cell_wire[74];							inform_L[85][4] = l_cell_wire[75];							inform_L[70][4] = l_cell_wire[76];							inform_L[86][4] = l_cell_wire[77];							inform_L[71][4] = l_cell_wire[78];							inform_L[87][4] = l_cell_wire[79];							inform_L[72][4] = l_cell_wire[80];							inform_L[88][4] = l_cell_wire[81];							inform_L[73][4] = l_cell_wire[82];							inform_L[89][4] = l_cell_wire[83];							inform_L[74][4] = l_cell_wire[84];							inform_L[90][4] = l_cell_wire[85];							inform_L[75][4] = l_cell_wire[86];							inform_L[91][4] = l_cell_wire[87];							inform_L[76][4] = l_cell_wire[88];							inform_L[92][4] = l_cell_wire[89];							inform_L[77][4] = l_cell_wire[90];							inform_L[93][4] = l_cell_wire[91];							inform_L[78][4] = l_cell_wire[92];							inform_L[94][4] = l_cell_wire[93];							inform_L[79][4] = l_cell_wire[94];							inform_L[95][4] = l_cell_wire[95];							inform_L[96][4] = l_cell_wire[96];							inform_L[112][4] = l_cell_wire[97];							inform_L[97][4] = l_cell_wire[98];							inform_L[113][4] = l_cell_wire[99];							inform_L[98][4] = l_cell_wire[100];							inform_L[114][4] = l_cell_wire[101];							inform_L[99][4] = l_cell_wire[102];							inform_L[115][4] = l_cell_wire[103];							inform_L[100][4] = l_cell_wire[104];							inform_L[116][4] = l_cell_wire[105];							inform_L[101][4] = l_cell_wire[106];							inform_L[117][4] = l_cell_wire[107];							inform_L[102][4] = l_cell_wire[108];							inform_L[118][4] = l_cell_wire[109];							inform_L[103][4] = l_cell_wire[110];							inform_L[119][4] = l_cell_wire[111];							inform_L[104][4] = l_cell_wire[112];							inform_L[120][4] = l_cell_wire[113];							inform_L[105][4] = l_cell_wire[114];							inform_L[121][4] = l_cell_wire[115];							inform_L[106][4] = l_cell_wire[116];							inform_L[122][4] = l_cell_wire[117];							inform_L[107][4] = l_cell_wire[118];							inform_L[123][4] = l_cell_wire[119];							inform_L[108][4] = l_cell_wire[120];							inform_L[124][4] = l_cell_wire[121];							inform_L[109][4] = l_cell_wire[122];							inform_L[125][4] = l_cell_wire[123];							inform_L[110][4] = l_cell_wire[124];							inform_L[126][4] = l_cell_wire[125];							inform_L[111][4] = l_cell_wire[126];							inform_L[127][4] = l_cell_wire[127];							inform_L[128][4] = l_cell_wire[128];							inform_L[144][4] = l_cell_wire[129];							inform_L[129][4] = l_cell_wire[130];							inform_L[145][4] = l_cell_wire[131];							inform_L[130][4] = l_cell_wire[132];							inform_L[146][4] = l_cell_wire[133];							inform_L[131][4] = l_cell_wire[134];							inform_L[147][4] = l_cell_wire[135];							inform_L[132][4] = l_cell_wire[136];							inform_L[148][4] = l_cell_wire[137];							inform_L[133][4] = l_cell_wire[138];							inform_L[149][4] = l_cell_wire[139];							inform_L[134][4] = l_cell_wire[140];							inform_L[150][4] = l_cell_wire[141];							inform_L[135][4] = l_cell_wire[142];							inform_L[151][4] = l_cell_wire[143];							inform_L[136][4] = l_cell_wire[144];							inform_L[152][4] = l_cell_wire[145];							inform_L[137][4] = l_cell_wire[146];							inform_L[153][4] = l_cell_wire[147];							inform_L[138][4] = l_cell_wire[148];							inform_L[154][4] = l_cell_wire[149];							inform_L[139][4] = l_cell_wire[150];							inform_L[155][4] = l_cell_wire[151];							inform_L[140][4] = l_cell_wire[152];							inform_L[156][4] = l_cell_wire[153];							inform_L[141][4] = l_cell_wire[154];							inform_L[157][4] = l_cell_wire[155];							inform_L[142][4] = l_cell_wire[156];							inform_L[158][4] = l_cell_wire[157];							inform_L[143][4] = l_cell_wire[158];							inform_L[159][4] = l_cell_wire[159];							inform_L[160][4] = l_cell_wire[160];							inform_L[176][4] = l_cell_wire[161];							inform_L[161][4] = l_cell_wire[162];							inform_L[177][4] = l_cell_wire[163];							inform_L[162][4] = l_cell_wire[164];							inform_L[178][4] = l_cell_wire[165];							inform_L[163][4] = l_cell_wire[166];							inform_L[179][4] = l_cell_wire[167];							inform_L[164][4] = l_cell_wire[168];							inform_L[180][4] = l_cell_wire[169];							inform_L[165][4] = l_cell_wire[170];							inform_L[181][4] = l_cell_wire[171];							inform_L[166][4] = l_cell_wire[172];							inform_L[182][4] = l_cell_wire[173];							inform_L[167][4] = l_cell_wire[174];							inform_L[183][4] = l_cell_wire[175];							inform_L[168][4] = l_cell_wire[176];							inform_L[184][4] = l_cell_wire[177];							inform_L[169][4] = l_cell_wire[178];							inform_L[185][4] = l_cell_wire[179];							inform_L[170][4] = l_cell_wire[180];							inform_L[186][4] = l_cell_wire[181];							inform_L[171][4] = l_cell_wire[182];							inform_L[187][4] = l_cell_wire[183];							inform_L[172][4] = l_cell_wire[184];							inform_L[188][4] = l_cell_wire[185];							inform_L[173][4] = l_cell_wire[186];							inform_L[189][4] = l_cell_wire[187];							inform_L[174][4] = l_cell_wire[188];							inform_L[190][4] = l_cell_wire[189];							inform_L[175][4] = l_cell_wire[190];							inform_L[191][4] = l_cell_wire[191];							inform_L[192][4] = l_cell_wire[192];							inform_L[208][4] = l_cell_wire[193];							inform_L[193][4] = l_cell_wire[194];							inform_L[209][4] = l_cell_wire[195];							inform_L[194][4] = l_cell_wire[196];							inform_L[210][4] = l_cell_wire[197];							inform_L[195][4] = l_cell_wire[198];							inform_L[211][4] = l_cell_wire[199];							inform_L[196][4] = l_cell_wire[200];							inform_L[212][4] = l_cell_wire[201];							inform_L[197][4] = l_cell_wire[202];							inform_L[213][4] = l_cell_wire[203];							inform_L[198][4] = l_cell_wire[204];							inform_L[214][4] = l_cell_wire[205];							inform_L[199][4] = l_cell_wire[206];							inform_L[215][4] = l_cell_wire[207];							inform_L[200][4] = l_cell_wire[208];							inform_L[216][4] = l_cell_wire[209];							inform_L[201][4] = l_cell_wire[210];							inform_L[217][4] = l_cell_wire[211];							inform_L[202][4] = l_cell_wire[212];							inform_L[218][4] = l_cell_wire[213];							inform_L[203][4] = l_cell_wire[214];							inform_L[219][4] = l_cell_wire[215];							inform_L[204][4] = l_cell_wire[216];							inform_L[220][4] = l_cell_wire[217];							inform_L[205][4] = l_cell_wire[218];							inform_L[221][4] = l_cell_wire[219];							inform_L[206][4] = l_cell_wire[220];							inform_L[222][4] = l_cell_wire[221];							inform_L[207][4] = l_cell_wire[222];							inform_L[223][4] = l_cell_wire[223];							inform_L[224][4] = l_cell_wire[224];							inform_L[240][4] = l_cell_wire[225];							inform_L[225][4] = l_cell_wire[226];							inform_L[241][4] = l_cell_wire[227];							inform_L[226][4] = l_cell_wire[228];							inform_L[242][4] = l_cell_wire[229];							inform_L[227][4] = l_cell_wire[230];							inform_L[243][4] = l_cell_wire[231];							inform_L[228][4] = l_cell_wire[232];							inform_L[244][4] = l_cell_wire[233];							inform_L[229][4] = l_cell_wire[234];							inform_L[245][4] = l_cell_wire[235];							inform_L[230][4] = l_cell_wire[236];							inform_L[246][4] = l_cell_wire[237];							inform_L[231][4] = l_cell_wire[238];							inform_L[247][4] = l_cell_wire[239];							inform_L[232][4] = l_cell_wire[240];							inform_L[248][4] = l_cell_wire[241];							inform_L[233][4] = l_cell_wire[242];							inform_L[249][4] = l_cell_wire[243];							inform_L[234][4] = l_cell_wire[244];							inform_L[250][4] = l_cell_wire[245];							inform_L[235][4] = l_cell_wire[246];							inform_L[251][4] = l_cell_wire[247];							inform_L[236][4] = l_cell_wire[248];							inform_L[252][4] = l_cell_wire[249];							inform_L[237][4] = l_cell_wire[250];							inform_L[253][4] = l_cell_wire[251];							inform_L[238][4] = l_cell_wire[252];							inform_L[254][4] = l_cell_wire[253];							inform_L[239][4] = l_cell_wire[254];							inform_L[255][4] = l_cell_wire[255];						end
						6:						begin							inform_R[0][6] = r_cell_wire[0];							inform_R[32][6] = r_cell_wire[1];							inform_R[1][6] = r_cell_wire[2];							inform_R[33][6] = r_cell_wire[3];							inform_R[2][6] = r_cell_wire[4];							inform_R[34][6] = r_cell_wire[5];							inform_R[3][6] = r_cell_wire[6];							inform_R[35][6] = r_cell_wire[7];							inform_R[4][6] = r_cell_wire[8];							inform_R[36][6] = r_cell_wire[9];							inform_R[5][6] = r_cell_wire[10];							inform_R[37][6] = r_cell_wire[11];							inform_R[6][6] = r_cell_wire[12];							inform_R[38][6] = r_cell_wire[13];							inform_R[7][6] = r_cell_wire[14];							inform_R[39][6] = r_cell_wire[15];							inform_R[8][6] = r_cell_wire[16];							inform_R[40][6] = r_cell_wire[17];							inform_R[9][6] = r_cell_wire[18];							inform_R[41][6] = r_cell_wire[19];							inform_R[10][6] = r_cell_wire[20];							inform_R[42][6] = r_cell_wire[21];							inform_R[11][6] = r_cell_wire[22];							inform_R[43][6] = r_cell_wire[23];							inform_R[12][6] = r_cell_wire[24];							inform_R[44][6] = r_cell_wire[25];							inform_R[13][6] = r_cell_wire[26];							inform_R[45][6] = r_cell_wire[27];							inform_R[14][6] = r_cell_wire[28];							inform_R[46][6] = r_cell_wire[29];							inform_R[15][6] = r_cell_wire[30];							inform_R[47][6] = r_cell_wire[31];							inform_R[16][6] = r_cell_wire[32];							inform_R[48][6] = r_cell_wire[33];							inform_R[17][6] = r_cell_wire[34];							inform_R[49][6] = r_cell_wire[35];							inform_R[18][6] = r_cell_wire[36];							inform_R[50][6] = r_cell_wire[37];							inform_R[19][6] = r_cell_wire[38];							inform_R[51][6] = r_cell_wire[39];							inform_R[20][6] = r_cell_wire[40];							inform_R[52][6] = r_cell_wire[41];							inform_R[21][6] = r_cell_wire[42];							inform_R[53][6] = r_cell_wire[43];							inform_R[22][6] = r_cell_wire[44];							inform_R[54][6] = r_cell_wire[45];							inform_R[23][6] = r_cell_wire[46];							inform_R[55][6] = r_cell_wire[47];							inform_R[24][6] = r_cell_wire[48];							inform_R[56][6] = r_cell_wire[49];							inform_R[25][6] = r_cell_wire[50];							inform_R[57][6] = r_cell_wire[51];							inform_R[26][6] = r_cell_wire[52];							inform_R[58][6] = r_cell_wire[53];							inform_R[27][6] = r_cell_wire[54];							inform_R[59][6] = r_cell_wire[55];							inform_R[28][6] = r_cell_wire[56];							inform_R[60][6] = r_cell_wire[57];							inform_R[29][6] = r_cell_wire[58];							inform_R[61][6] = r_cell_wire[59];							inform_R[30][6] = r_cell_wire[60];							inform_R[62][6] = r_cell_wire[61];							inform_R[31][6] = r_cell_wire[62];							inform_R[63][6] = r_cell_wire[63];							inform_R[64][6] = r_cell_wire[64];							inform_R[96][6] = r_cell_wire[65];							inform_R[65][6] = r_cell_wire[66];							inform_R[97][6] = r_cell_wire[67];							inform_R[66][6] = r_cell_wire[68];							inform_R[98][6] = r_cell_wire[69];							inform_R[67][6] = r_cell_wire[70];							inform_R[99][6] = r_cell_wire[71];							inform_R[68][6] = r_cell_wire[72];							inform_R[100][6] = r_cell_wire[73];							inform_R[69][6] = r_cell_wire[74];							inform_R[101][6] = r_cell_wire[75];							inform_R[70][6] = r_cell_wire[76];							inform_R[102][6] = r_cell_wire[77];							inform_R[71][6] = r_cell_wire[78];							inform_R[103][6] = r_cell_wire[79];							inform_R[72][6] = r_cell_wire[80];							inform_R[104][6] = r_cell_wire[81];							inform_R[73][6] = r_cell_wire[82];							inform_R[105][6] = r_cell_wire[83];							inform_R[74][6] = r_cell_wire[84];							inform_R[106][6] = r_cell_wire[85];							inform_R[75][6] = r_cell_wire[86];							inform_R[107][6] = r_cell_wire[87];							inform_R[76][6] = r_cell_wire[88];							inform_R[108][6] = r_cell_wire[89];							inform_R[77][6] = r_cell_wire[90];							inform_R[109][6] = r_cell_wire[91];							inform_R[78][6] = r_cell_wire[92];							inform_R[110][6] = r_cell_wire[93];							inform_R[79][6] = r_cell_wire[94];							inform_R[111][6] = r_cell_wire[95];							inform_R[80][6] = r_cell_wire[96];							inform_R[112][6] = r_cell_wire[97];							inform_R[81][6] = r_cell_wire[98];							inform_R[113][6] = r_cell_wire[99];							inform_R[82][6] = r_cell_wire[100];							inform_R[114][6] = r_cell_wire[101];							inform_R[83][6] = r_cell_wire[102];							inform_R[115][6] = r_cell_wire[103];							inform_R[84][6] = r_cell_wire[104];							inform_R[116][6] = r_cell_wire[105];							inform_R[85][6] = r_cell_wire[106];							inform_R[117][6] = r_cell_wire[107];							inform_R[86][6] = r_cell_wire[108];							inform_R[118][6] = r_cell_wire[109];							inform_R[87][6] = r_cell_wire[110];							inform_R[119][6] = r_cell_wire[111];							inform_R[88][6] = r_cell_wire[112];							inform_R[120][6] = r_cell_wire[113];							inform_R[89][6] = r_cell_wire[114];							inform_R[121][6] = r_cell_wire[115];							inform_R[90][6] = r_cell_wire[116];							inform_R[122][6] = r_cell_wire[117];							inform_R[91][6] = r_cell_wire[118];							inform_R[123][6] = r_cell_wire[119];							inform_R[92][6] = r_cell_wire[120];							inform_R[124][6] = r_cell_wire[121];							inform_R[93][6] = r_cell_wire[122];							inform_R[125][6] = r_cell_wire[123];							inform_R[94][6] = r_cell_wire[124];							inform_R[126][6] = r_cell_wire[125];							inform_R[95][6] = r_cell_wire[126];							inform_R[127][6] = r_cell_wire[127];							inform_R[128][6] = r_cell_wire[128];							inform_R[160][6] = r_cell_wire[129];							inform_R[129][6] = r_cell_wire[130];							inform_R[161][6] = r_cell_wire[131];							inform_R[130][6] = r_cell_wire[132];							inform_R[162][6] = r_cell_wire[133];							inform_R[131][6] = r_cell_wire[134];							inform_R[163][6] = r_cell_wire[135];							inform_R[132][6] = r_cell_wire[136];							inform_R[164][6] = r_cell_wire[137];							inform_R[133][6] = r_cell_wire[138];							inform_R[165][6] = r_cell_wire[139];							inform_R[134][6] = r_cell_wire[140];							inform_R[166][6] = r_cell_wire[141];							inform_R[135][6] = r_cell_wire[142];							inform_R[167][6] = r_cell_wire[143];							inform_R[136][6] = r_cell_wire[144];							inform_R[168][6] = r_cell_wire[145];							inform_R[137][6] = r_cell_wire[146];							inform_R[169][6] = r_cell_wire[147];							inform_R[138][6] = r_cell_wire[148];							inform_R[170][6] = r_cell_wire[149];							inform_R[139][6] = r_cell_wire[150];							inform_R[171][6] = r_cell_wire[151];							inform_R[140][6] = r_cell_wire[152];							inform_R[172][6] = r_cell_wire[153];							inform_R[141][6] = r_cell_wire[154];							inform_R[173][6] = r_cell_wire[155];							inform_R[142][6] = r_cell_wire[156];							inform_R[174][6] = r_cell_wire[157];							inform_R[143][6] = r_cell_wire[158];							inform_R[175][6] = r_cell_wire[159];							inform_R[144][6] = r_cell_wire[160];							inform_R[176][6] = r_cell_wire[161];							inform_R[145][6] = r_cell_wire[162];							inform_R[177][6] = r_cell_wire[163];							inform_R[146][6] = r_cell_wire[164];							inform_R[178][6] = r_cell_wire[165];							inform_R[147][6] = r_cell_wire[166];							inform_R[179][6] = r_cell_wire[167];							inform_R[148][6] = r_cell_wire[168];							inform_R[180][6] = r_cell_wire[169];							inform_R[149][6] = r_cell_wire[170];							inform_R[181][6] = r_cell_wire[171];							inform_R[150][6] = r_cell_wire[172];							inform_R[182][6] = r_cell_wire[173];							inform_R[151][6] = r_cell_wire[174];							inform_R[183][6] = r_cell_wire[175];							inform_R[152][6] = r_cell_wire[176];							inform_R[184][6] = r_cell_wire[177];							inform_R[153][6] = r_cell_wire[178];							inform_R[185][6] = r_cell_wire[179];							inform_R[154][6] = r_cell_wire[180];							inform_R[186][6] = r_cell_wire[181];							inform_R[155][6] = r_cell_wire[182];							inform_R[187][6] = r_cell_wire[183];							inform_R[156][6] = r_cell_wire[184];							inform_R[188][6] = r_cell_wire[185];							inform_R[157][6] = r_cell_wire[186];							inform_R[189][6] = r_cell_wire[187];							inform_R[158][6] = r_cell_wire[188];							inform_R[190][6] = r_cell_wire[189];							inform_R[159][6] = r_cell_wire[190];							inform_R[191][6] = r_cell_wire[191];							inform_R[192][6] = r_cell_wire[192];							inform_R[224][6] = r_cell_wire[193];							inform_R[193][6] = r_cell_wire[194];							inform_R[225][6] = r_cell_wire[195];							inform_R[194][6] = r_cell_wire[196];							inform_R[226][6] = r_cell_wire[197];							inform_R[195][6] = r_cell_wire[198];							inform_R[227][6] = r_cell_wire[199];							inform_R[196][6] = r_cell_wire[200];							inform_R[228][6] = r_cell_wire[201];							inform_R[197][6] = r_cell_wire[202];							inform_R[229][6] = r_cell_wire[203];							inform_R[198][6] = r_cell_wire[204];							inform_R[230][6] = r_cell_wire[205];							inform_R[199][6] = r_cell_wire[206];							inform_R[231][6] = r_cell_wire[207];							inform_R[200][6] = r_cell_wire[208];							inform_R[232][6] = r_cell_wire[209];							inform_R[201][6] = r_cell_wire[210];							inform_R[233][6] = r_cell_wire[211];							inform_R[202][6] = r_cell_wire[212];							inform_R[234][6] = r_cell_wire[213];							inform_R[203][6] = r_cell_wire[214];							inform_R[235][6] = r_cell_wire[215];							inform_R[204][6] = r_cell_wire[216];							inform_R[236][6] = r_cell_wire[217];							inform_R[205][6] = r_cell_wire[218];							inform_R[237][6] = r_cell_wire[219];							inform_R[206][6] = r_cell_wire[220];							inform_R[238][6] = r_cell_wire[221];							inform_R[207][6] = r_cell_wire[222];							inform_R[239][6] = r_cell_wire[223];							inform_R[208][6] = r_cell_wire[224];							inform_R[240][6] = r_cell_wire[225];							inform_R[209][6] = r_cell_wire[226];							inform_R[241][6] = r_cell_wire[227];							inform_R[210][6] = r_cell_wire[228];							inform_R[242][6] = r_cell_wire[229];							inform_R[211][6] = r_cell_wire[230];							inform_R[243][6] = r_cell_wire[231];							inform_R[212][6] = r_cell_wire[232];							inform_R[244][6] = r_cell_wire[233];							inform_R[213][6] = r_cell_wire[234];							inform_R[245][6] = r_cell_wire[235];							inform_R[214][6] = r_cell_wire[236];							inform_R[246][6] = r_cell_wire[237];							inform_R[215][6] = r_cell_wire[238];							inform_R[247][6] = r_cell_wire[239];							inform_R[216][6] = r_cell_wire[240];							inform_R[248][6] = r_cell_wire[241];							inform_R[217][6] = r_cell_wire[242];							inform_R[249][6] = r_cell_wire[243];							inform_R[218][6] = r_cell_wire[244];							inform_R[250][6] = r_cell_wire[245];							inform_R[219][6] = r_cell_wire[246];							inform_R[251][6] = r_cell_wire[247];							inform_R[220][6] = r_cell_wire[248];							inform_R[252][6] = r_cell_wire[249];							inform_R[221][6] = r_cell_wire[250];							inform_R[253][6] = r_cell_wire[251];							inform_R[222][6] = r_cell_wire[252];							inform_R[254][6] = r_cell_wire[253];							inform_R[223][6] = r_cell_wire[254];							inform_R[255][6] = r_cell_wire[255];							inform_L[0][5] = l_cell_wire[0];							inform_L[32][5] = l_cell_wire[1];							inform_L[1][5] = l_cell_wire[2];							inform_L[33][5] = l_cell_wire[3];							inform_L[2][5] = l_cell_wire[4];							inform_L[34][5] = l_cell_wire[5];							inform_L[3][5] = l_cell_wire[6];							inform_L[35][5] = l_cell_wire[7];							inform_L[4][5] = l_cell_wire[8];							inform_L[36][5] = l_cell_wire[9];							inform_L[5][5] = l_cell_wire[10];							inform_L[37][5] = l_cell_wire[11];							inform_L[6][5] = l_cell_wire[12];							inform_L[38][5] = l_cell_wire[13];							inform_L[7][5] = l_cell_wire[14];							inform_L[39][5] = l_cell_wire[15];							inform_L[8][5] = l_cell_wire[16];							inform_L[40][5] = l_cell_wire[17];							inform_L[9][5] = l_cell_wire[18];							inform_L[41][5] = l_cell_wire[19];							inform_L[10][5] = l_cell_wire[20];							inform_L[42][5] = l_cell_wire[21];							inform_L[11][5] = l_cell_wire[22];							inform_L[43][5] = l_cell_wire[23];							inform_L[12][5] = l_cell_wire[24];							inform_L[44][5] = l_cell_wire[25];							inform_L[13][5] = l_cell_wire[26];							inform_L[45][5] = l_cell_wire[27];							inform_L[14][5] = l_cell_wire[28];							inform_L[46][5] = l_cell_wire[29];							inform_L[15][5] = l_cell_wire[30];							inform_L[47][5] = l_cell_wire[31];							inform_L[16][5] = l_cell_wire[32];							inform_L[48][5] = l_cell_wire[33];							inform_L[17][5] = l_cell_wire[34];							inform_L[49][5] = l_cell_wire[35];							inform_L[18][5] = l_cell_wire[36];							inform_L[50][5] = l_cell_wire[37];							inform_L[19][5] = l_cell_wire[38];							inform_L[51][5] = l_cell_wire[39];							inform_L[20][5] = l_cell_wire[40];							inform_L[52][5] = l_cell_wire[41];							inform_L[21][5] = l_cell_wire[42];							inform_L[53][5] = l_cell_wire[43];							inform_L[22][5] = l_cell_wire[44];							inform_L[54][5] = l_cell_wire[45];							inform_L[23][5] = l_cell_wire[46];							inform_L[55][5] = l_cell_wire[47];							inform_L[24][5] = l_cell_wire[48];							inform_L[56][5] = l_cell_wire[49];							inform_L[25][5] = l_cell_wire[50];							inform_L[57][5] = l_cell_wire[51];							inform_L[26][5] = l_cell_wire[52];							inform_L[58][5] = l_cell_wire[53];							inform_L[27][5] = l_cell_wire[54];							inform_L[59][5] = l_cell_wire[55];							inform_L[28][5] = l_cell_wire[56];							inform_L[60][5] = l_cell_wire[57];							inform_L[29][5] = l_cell_wire[58];							inform_L[61][5] = l_cell_wire[59];							inform_L[30][5] = l_cell_wire[60];							inform_L[62][5] = l_cell_wire[61];							inform_L[31][5] = l_cell_wire[62];							inform_L[63][5] = l_cell_wire[63];							inform_L[64][5] = l_cell_wire[64];							inform_L[96][5] = l_cell_wire[65];							inform_L[65][5] = l_cell_wire[66];							inform_L[97][5] = l_cell_wire[67];							inform_L[66][5] = l_cell_wire[68];							inform_L[98][5] = l_cell_wire[69];							inform_L[67][5] = l_cell_wire[70];							inform_L[99][5] = l_cell_wire[71];							inform_L[68][5] = l_cell_wire[72];							inform_L[100][5] = l_cell_wire[73];							inform_L[69][5] = l_cell_wire[74];							inform_L[101][5] = l_cell_wire[75];							inform_L[70][5] = l_cell_wire[76];							inform_L[102][5] = l_cell_wire[77];							inform_L[71][5] = l_cell_wire[78];							inform_L[103][5] = l_cell_wire[79];							inform_L[72][5] = l_cell_wire[80];							inform_L[104][5] = l_cell_wire[81];							inform_L[73][5] = l_cell_wire[82];							inform_L[105][5] = l_cell_wire[83];							inform_L[74][5] = l_cell_wire[84];							inform_L[106][5] = l_cell_wire[85];							inform_L[75][5] = l_cell_wire[86];							inform_L[107][5] = l_cell_wire[87];							inform_L[76][5] = l_cell_wire[88];							inform_L[108][5] = l_cell_wire[89];							inform_L[77][5] = l_cell_wire[90];							inform_L[109][5] = l_cell_wire[91];							inform_L[78][5] = l_cell_wire[92];							inform_L[110][5] = l_cell_wire[93];							inform_L[79][5] = l_cell_wire[94];							inform_L[111][5] = l_cell_wire[95];							inform_L[80][5] = l_cell_wire[96];							inform_L[112][5] = l_cell_wire[97];							inform_L[81][5] = l_cell_wire[98];							inform_L[113][5] = l_cell_wire[99];							inform_L[82][5] = l_cell_wire[100];							inform_L[114][5] = l_cell_wire[101];							inform_L[83][5] = l_cell_wire[102];							inform_L[115][5] = l_cell_wire[103];							inform_L[84][5] = l_cell_wire[104];							inform_L[116][5] = l_cell_wire[105];							inform_L[85][5] = l_cell_wire[106];							inform_L[117][5] = l_cell_wire[107];							inform_L[86][5] = l_cell_wire[108];							inform_L[118][5] = l_cell_wire[109];							inform_L[87][5] = l_cell_wire[110];							inform_L[119][5] = l_cell_wire[111];							inform_L[88][5] = l_cell_wire[112];							inform_L[120][5] = l_cell_wire[113];							inform_L[89][5] = l_cell_wire[114];							inform_L[121][5] = l_cell_wire[115];							inform_L[90][5] = l_cell_wire[116];							inform_L[122][5] = l_cell_wire[117];							inform_L[91][5] = l_cell_wire[118];							inform_L[123][5] = l_cell_wire[119];							inform_L[92][5] = l_cell_wire[120];							inform_L[124][5] = l_cell_wire[121];							inform_L[93][5] = l_cell_wire[122];							inform_L[125][5] = l_cell_wire[123];							inform_L[94][5] = l_cell_wire[124];							inform_L[126][5] = l_cell_wire[125];							inform_L[95][5] = l_cell_wire[126];							inform_L[127][5] = l_cell_wire[127];							inform_L[128][5] = l_cell_wire[128];							inform_L[160][5] = l_cell_wire[129];							inform_L[129][5] = l_cell_wire[130];							inform_L[161][5] = l_cell_wire[131];							inform_L[130][5] = l_cell_wire[132];							inform_L[162][5] = l_cell_wire[133];							inform_L[131][5] = l_cell_wire[134];							inform_L[163][5] = l_cell_wire[135];							inform_L[132][5] = l_cell_wire[136];							inform_L[164][5] = l_cell_wire[137];							inform_L[133][5] = l_cell_wire[138];							inform_L[165][5] = l_cell_wire[139];							inform_L[134][5] = l_cell_wire[140];							inform_L[166][5] = l_cell_wire[141];							inform_L[135][5] = l_cell_wire[142];							inform_L[167][5] = l_cell_wire[143];							inform_L[136][5] = l_cell_wire[144];							inform_L[168][5] = l_cell_wire[145];							inform_L[137][5] = l_cell_wire[146];							inform_L[169][5] = l_cell_wire[147];							inform_L[138][5] = l_cell_wire[148];							inform_L[170][5] = l_cell_wire[149];							inform_L[139][5] = l_cell_wire[150];							inform_L[171][5] = l_cell_wire[151];							inform_L[140][5] = l_cell_wire[152];							inform_L[172][5] = l_cell_wire[153];							inform_L[141][5] = l_cell_wire[154];							inform_L[173][5] = l_cell_wire[155];							inform_L[142][5] = l_cell_wire[156];							inform_L[174][5] = l_cell_wire[157];							inform_L[143][5] = l_cell_wire[158];							inform_L[175][5] = l_cell_wire[159];							inform_L[144][5] = l_cell_wire[160];							inform_L[176][5] = l_cell_wire[161];							inform_L[145][5] = l_cell_wire[162];							inform_L[177][5] = l_cell_wire[163];							inform_L[146][5] = l_cell_wire[164];							inform_L[178][5] = l_cell_wire[165];							inform_L[147][5] = l_cell_wire[166];							inform_L[179][5] = l_cell_wire[167];							inform_L[148][5] = l_cell_wire[168];							inform_L[180][5] = l_cell_wire[169];							inform_L[149][5] = l_cell_wire[170];							inform_L[181][5] = l_cell_wire[171];							inform_L[150][5] = l_cell_wire[172];							inform_L[182][5] = l_cell_wire[173];							inform_L[151][5] = l_cell_wire[174];							inform_L[183][5] = l_cell_wire[175];							inform_L[152][5] = l_cell_wire[176];							inform_L[184][5] = l_cell_wire[177];							inform_L[153][5] = l_cell_wire[178];							inform_L[185][5] = l_cell_wire[179];							inform_L[154][5] = l_cell_wire[180];							inform_L[186][5] = l_cell_wire[181];							inform_L[155][5] = l_cell_wire[182];							inform_L[187][5] = l_cell_wire[183];							inform_L[156][5] = l_cell_wire[184];							inform_L[188][5] = l_cell_wire[185];							inform_L[157][5] = l_cell_wire[186];							inform_L[189][5] = l_cell_wire[187];							inform_L[158][5] = l_cell_wire[188];							inform_L[190][5] = l_cell_wire[189];							inform_L[159][5] = l_cell_wire[190];							inform_L[191][5] = l_cell_wire[191];							inform_L[192][5] = l_cell_wire[192];							inform_L[224][5] = l_cell_wire[193];							inform_L[193][5] = l_cell_wire[194];							inform_L[225][5] = l_cell_wire[195];							inform_L[194][5] = l_cell_wire[196];							inform_L[226][5] = l_cell_wire[197];							inform_L[195][5] = l_cell_wire[198];							inform_L[227][5] = l_cell_wire[199];							inform_L[196][5] = l_cell_wire[200];							inform_L[228][5] = l_cell_wire[201];							inform_L[197][5] = l_cell_wire[202];							inform_L[229][5] = l_cell_wire[203];							inform_L[198][5] = l_cell_wire[204];							inform_L[230][5] = l_cell_wire[205];							inform_L[199][5] = l_cell_wire[206];							inform_L[231][5] = l_cell_wire[207];							inform_L[200][5] = l_cell_wire[208];							inform_L[232][5] = l_cell_wire[209];							inform_L[201][5] = l_cell_wire[210];							inform_L[233][5] = l_cell_wire[211];							inform_L[202][5] = l_cell_wire[212];							inform_L[234][5] = l_cell_wire[213];							inform_L[203][5] = l_cell_wire[214];							inform_L[235][5] = l_cell_wire[215];							inform_L[204][5] = l_cell_wire[216];							inform_L[236][5] = l_cell_wire[217];							inform_L[205][5] = l_cell_wire[218];							inform_L[237][5] = l_cell_wire[219];							inform_L[206][5] = l_cell_wire[220];							inform_L[238][5] = l_cell_wire[221];							inform_L[207][5] = l_cell_wire[222];							inform_L[239][5] = l_cell_wire[223];							inform_L[208][5] = l_cell_wire[224];							inform_L[240][5] = l_cell_wire[225];							inform_L[209][5] = l_cell_wire[226];							inform_L[241][5] = l_cell_wire[227];							inform_L[210][5] = l_cell_wire[228];							inform_L[242][5] = l_cell_wire[229];							inform_L[211][5] = l_cell_wire[230];							inform_L[243][5] = l_cell_wire[231];							inform_L[212][5] = l_cell_wire[232];							inform_L[244][5] = l_cell_wire[233];							inform_L[213][5] = l_cell_wire[234];							inform_L[245][5] = l_cell_wire[235];							inform_L[214][5] = l_cell_wire[236];							inform_L[246][5] = l_cell_wire[237];							inform_L[215][5] = l_cell_wire[238];							inform_L[247][5] = l_cell_wire[239];							inform_L[216][5] = l_cell_wire[240];							inform_L[248][5] = l_cell_wire[241];							inform_L[217][5] = l_cell_wire[242];							inform_L[249][5] = l_cell_wire[243];							inform_L[218][5] = l_cell_wire[244];							inform_L[250][5] = l_cell_wire[245];							inform_L[219][5] = l_cell_wire[246];							inform_L[251][5] = l_cell_wire[247];							inform_L[220][5] = l_cell_wire[248];							inform_L[252][5] = l_cell_wire[249];							inform_L[221][5] = l_cell_wire[250];							inform_L[253][5] = l_cell_wire[251];							inform_L[222][5] = l_cell_wire[252];							inform_L[254][5] = l_cell_wire[253];							inform_L[223][5] = l_cell_wire[254];							inform_L[255][5] = l_cell_wire[255];						end
						7:						begin							inform_R[0][7] = r_cell_wire[0];							inform_R[64][7] = r_cell_wire[1];							inform_R[1][7] = r_cell_wire[2];							inform_R[65][7] = r_cell_wire[3];							inform_R[2][7] = r_cell_wire[4];							inform_R[66][7] = r_cell_wire[5];							inform_R[3][7] = r_cell_wire[6];							inform_R[67][7] = r_cell_wire[7];							inform_R[4][7] = r_cell_wire[8];							inform_R[68][7] = r_cell_wire[9];							inform_R[5][7] = r_cell_wire[10];							inform_R[69][7] = r_cell_wire[11];							inform_R[6][7] = r_cell_wire[12];							inform_R[70][7] = r_cell_wire[13];							inform_R[7][7] = r_cell_wire[14];							inform_R[71][7] = r_cell_wire[15];							inform_R[8][7] = r_cell_wire[16];							inform_R[72][7] = r_cell_wire[17];							inform_R[9][7] = r_cell_wire[18];							inform_R[73][7] = r_cell_wire[19];							inform_R[10][7] = r_cell_wire[20];							inform_R[74][7] = r_cell_wire[21];							inform_R[11][7] = r_cell_wire[22];							inform_R[75][7] = r_cell_wire[23];							inform_R[12][7] = r_cell_wire[24];							inform_R[76][7] = r_cell_wire[25];							inform_R[13][7] = r_cell_wire[26];							inform_R[77][7] = r_cell_wire[27];							inform_R[14][7] = r_cell_wire[28];							inform_R[78][7] = r_cell_wire[29];							inform_R[15][7] = r_cell_wire[30];							inform_R[79][7] = r_cell_wire[31];							inform_R[16][7] = r_cell_wire[32];							inform_R[80][7] = r_cell_wire[33];							inform_R[17][7] = r_cell_wire[34];							inform_R[81][7] = r_cell_wire[35];							inform_R[18][7] = r_cell_wire[36];							inform_R[82][7] = r_cell_wire[37];							inform_R[19][7] = r_cell_wire[38];							inform_R[83][7] = r_cell_wire[39];							inform_R[20][7] = r_cell_wire[40];							inform_R[84][7] = r_cell_wire[41];							inform_R[21][7] = r_cell_wire[42];							inform_R[85][7] = r_cell_wire[43];							inform_R[22][7] = r_cell_wire[44];							inform_R[86][7] = r_cell_wire[45];							inform_R[23][7] = r_cell_wire[46];							inform_R[87][7] = r_cell_wire[47];							inform_R[24][7] = r_cell_wire[48];							inform_R[88][7] = r_cell_wire[49];							inform_R[25][7] = r_cell_wire[50];							inform_R[89][7] = r_cell_wire[51];							inform_R[26][7] = r_cell_wire[52];							inform_R[90][7] = r_cell_wire[53];							inform_R[27][7] = r_cell_wire[54];							inform_R[91][7] = r_cell_wire[55];							inform_R[28][7] = r_cell_wire[56];							inform_R[92][7] = r_cell_wire[57];							inform_R[29][7] = r_cell_wire[58];							inform_R[93][7] = r_cell_wire[59];							inform_R[30][7] = r_cell_wire[60];							inform_R[94][7] = r_cell_wire[61];							inform_R[31][7] = r_cell_wire[62];							inform_R[95][7] = r_cell_wire[63];							inform_R[32][7] = r_cell_wire[64];							inform_R[96][7] = r_cell_wire[65];							inform_R[33][7] = r_cell_wire[66];							inform_R[97][7] = r_cell_wire[67];							inform_R[34][7] = r_cell_wire[68];							inform_R[98][7] = r_cell_wire[69];							inform_R[35][7] = r_cell_wire[70];							inform_R[99][7] = r_cell_wire[71];							inform_R[36][7] = r_cell_wire[72];							inform_R[100][7] = r_cell_wire[73];							inform_R[37][7] = r_cell_wire[74];							inform_R[101][7] = r_cell_wire[75];							inform_R[38][7] = r_cell_wire[76];							inform_R[102][7] = r_cell_wire[77];							inform_R[39][7] = r_cell_wire[78];							inform_R[103][7] = r_cell_wire[79];							inform_R[40][7] = r_cell_wire[80];							inform_R[104][7] = r_cell_wire[81];							inform_R[41][7] = r_cell_wire[82];							inform_R[105][7] = r_cell_wire[83];							inform_R[42][7] = r_cell_wire[84];							inform_R[106][7] = r_cell_wire[85];							inform_R[43][7] = r_cell_wire[86];							inform_R[107][7] = r_cell_wire[87];							inform_R[44][7] = r_cell_wire[88];							inform_R[108][7] = r_cell_wire[89];							inform_R[45][7] = r_cell_wire[90];							inform_R[109][7] = r_cell_wire[91];							inform_R[46][7] = r_cell_wire[92];							inform_R[110][7] = r_cell_wire[93];							inform_R[47][7] = r_cell_wire[94];							inform_R[111][7] = r_cell_wire[95];							inform_R[48][7] = r_cell_wire[96];							inform_R[112][7] = r_cell_wire[97];							inform_R[49][7] = r_cell_wire[98];							inform_R[113][7] = r_cell_wire[99];							inform_R[50][7] = r_cell_wire[100];							inform_R[114][7] = r_cell_wire[101];							inform_R[51][7] = r_cell_wire[102];							inform_R[115][7] = r_cell_wire[103];							inform_R[52][7] = r_cell_wire[104];							inform_R[116][7] = r_cell_wire[105];							inform_R[53][7] = r_cell_wire[106];							inform_R[117][7] = r_cell_wire[107];							inform_R[54][7] = r_cell_wire[108];							inform_R[118][7] = r_cell_wire[109];							inform_R[55][7] = r_cell_wire[110];							inform_R[119][7] = r_cell_wire[111];							inform_R[56][7] = r_cell_wire[112];							inform_R[120][7] = r_cell_wire[113];							inform_R[57][7] = r_cell_wire[114];							inform_R[121][7] = r_cell_wire[115];							inform_R[58][7] = r_cell_wire[116];							inform_R[122][7] = r_cell_wire[117];							inform_R[59][7] = r_cell_wire[118];							inform_R[123][7] = r_cell_wire[119];							inform_R[60][7] = r_cell_wire[120];							inform_R[124][7] = r_cell_wire[121];							inform_R[61][7] = r_cell_wire[122];							inform_R[125][7] = r_cell_wire[123];							inform_R[62][7] = r_cell_wire[124];							inform_R[126][7] = r_cell_wire[125];							inform_R[63][7] = r_cell_wire[126];							inform_R[127][7] = r_cell_wire[127];							inform_R[128][7] = r_cell_wire[128];							inform_R[192][7] = r_cell_wire[129];							inform_R[129][7] = r_cell_wire[130];							inform_R[193][7] = r_cell_wire[131];							inform_R[130][7] = r_cell_wire[132];							inform_R[194][7] = r_cell_wire[133];							inform_R[131][7] = r_cell_wire[134];							inform_R[195][7] = r_cell_wire[135];							inform_R[132][7] = r_cell_wire[136];							inform_R[196][7] = r_cell_wire[137];							inform_R[133][7] = r_cell_wire[138];							inform_R[197][7] = r_cell_wire[139];							inform_R[134][7] = r_cell_wire[140];							inform_R[198][7] = r_cell_wire[141];							inform_R[135][7] = r_cell_wire[142];							inform_R[199][7] = r_cell_wire[143];							inform_R[136][7] = r_cell_wire[144];							inform_R[200][7] = r_cell_wire[145];							inform_R[137][7] = r_cell_wire[146];							inform_R[201][7] = r_cell_wire[147];							inform_R[138][7] = r_cell_wire[148];							inform_R[202][7] = r_cell_wire[149];							inform_R[139][7] = r_cell_wire[150];							inform_R[203][7] = r_cell_wire[151];							inform_R[140][7] = r_cell_wire[152];							inform_R[204][7] = r_cell_wire[153];							inform_R[141][7] = r_cell_wire[154];							inform_R[205][7] = r_cell_wire[155];							inform_R[142][7] = r_cell_wire[156];							inform_R[206][7] = r_cell_wire[157];							inform_R[143][7] = r_cell_wire[158];							inform_R[207][7] = r_cell_wire[159];							inform_R[144][7] = r_cell_wire[160];							inform_R[208][7] = r_cell_wire[161];							inform_R[145][7] = r_cell_wire[162];							inform_R[209][7] = r_cell_wire[163];							inform_R[146][7] = r_cell_wire[164];							inform_R[210][7] = r_cell_wire[165];							inform_R[147][7] = r_cell_wire[166];							inform_R[211][7] = r_cell_wire[167];							inform_R[148][7] = r_cell_wire[168];							inform_R[212][7] = r_cell_wire[169];							inform_R[149][7] = r_cell_wire[170];							inform_R[213][7] = r_cell_wire[171];							inform_R[150][7] = r_cell_wire[172];							inform_R[214][7] = r_cell_wire[173];							inform_R[151][7] = r_cell_wire[174];							inform_R[215][7] = r_cell_wire[175];							inform_R[152][7] = r_cell_wire[176];							inform_R[216][7] = r_cell_wire[177];							inform_R[153][7] = r_cell_wire[178];							inform_R[217][7] = r_cell_wire[179];							inform_R[154][7] = r_cell_wire[180];							inform_R[218][7] = r_cell_wire[181];							inform_R[155][7] = r_cell_wire[182];							inform_R[219][7] = r_cell_wire[183];							inform_R[156][7] = r_cell_wire[184];							inform_R[220][7] = r_cell_wire[185];							inform_R[157][7] = r_cell_wire[186];							inform_R[221][7] = r_cell_wire[187];							inform_R[158][7] = r_cell_wire[188];							inform_R[222][7] = r_cell_wire[189];							inform_R[159][7] = r_cell_wire[190];							inform_R[223][7] = r_cell_wire[191];							inform_R[160][7] = r_cell_wire[192];							inform_R[224][7] = r_cell_wire[193];							inform_R[161][7] = r_cell_wire[194];							inform_R[225][7] = r_cell_wire[195];							inform_R[162][7] = r_cell_wire[196];							inform_R[226][7] = r_cell_wire[197];							inform_R[163][7] = r_cell_wire[198];							inform_R[227][7] = r_cell_wire[199];							inform_R[164][7] = r_cell_wire[200];							inform_R[228][7] = r_cell_wire[201];							inform_R[165][7] = r_cell_wire[202];							inform_R[229][7] = r_cell_wire[203];							inform_R[166][7] = r_cell_wire[204];							inform_R[230][7] = r_cell_wire[205];							inform_R[167][7] = r_cell_wire[206];							inform_R[231][7] = r_cell_wire[207];							inform_R[168][7] = r_cell_wire[208];							inform_R[232][7] = r_cell_wire[209];							inform_R[169][7] = r_cell_wire[210];							inform_R[233][7] = r_cell_wire[211];							inform_R[170][7] = r_cell_wire[212];							inform_R[234][7] = r_cell_wire[213];							inform_R[171][7] = r_cell_wire[214];							inform_R[235][7] = r_cell_wire[215];							inform_R[172][7] = r_cell_wire[216];							inform_R[236][7] = r_cell_wire[217];							inform_R[173][7] = r_cell_wire[218];							inform_R[237][7] = r_cell_wire[219];							inform_R[174][7] = r_cell_wire[220];							inform_R[238][7] = r_cell_wire[221];							inform_R[175][7] = r_cell_wire[222];							inform_R[239][7] = r_cell_wire[223];							inform_R[176][7] = r_cell_wire[224];							inform_R[240][7] = r_cell_wire[225];							inform_R[177][7] = r_cell_wire[226];							inform_R[241][7] = r_cell_wire[227];							inform_R[178][7] = r_cell_wire[228];							inform_R[242][7] = r_cell_wire[229];							inform_R[179][7] = r_cell_wire[230];							inform_R[243][7] = r_cell_wire[231];							inform_R[180][7] = r_cell_wire[232];							inform_R[244][7] = r_cell_wire[233];							inform_R[181][7] = r_cell_wire[234];							inform_R[245][7] = r_cell_wire[235];							inform_R[182][7] = r_cell_wire[236];							inform_R[246][7] = r_cell_wire[237];							inform_R[183][7] = r_cell_wire[238];							inform_R[247][7] = r_cell_wire[239];							inform_R[184][7] = r_cell_wire[240];							inform_R[248][7] = r_cell_wire[241];							inform_R[185][7] = r_cell_wire[242];							inform_R[249][7] = r_cell_wire[243];							inform_R[186][7] = r_cell_wire[244];							inform_R[250][7] = r_cell_wire[245];							inform_R[187][7] = r_cell_wire[246];							inform_R[251][7] = r_cell_wire[247];							inform_R[188][7] = r_cell_wire[248];							inform_R[252][7] = r_cell_wire[249];							inform_R[189][7] = r_cell_wire[250];							inform_R[253][7] = r_cell_wire[251];							inform_R[190][7] = r_cell_wire[252];							inform_R[254][7] = r_cell_wire[253];							inform_R[191][7] = r_cell_wire[254];							inform_R[255][7] = r_cell_wire[255];							inform_L[0][6] = l_cell_wire[0];							inform_L[64][6] = l_cell_wire[1];							inform_L[1][6] = l_cell_wire[2];							inform_L[65][6] = l_cell_wire[3];							inform_L[2][6] = l_cell_wire[4];							inform_L[66][6] = l_cell_wire[5];							inform_L[3][6] = l_cell_wire[6];							inform_L[67][6] = l_cell_wire[7];							inform_L[4][6] = l_cell_wire[8];							inform_L[68][6] = l_cell_wire[9];							inform_L[5][6] = l_cell_wire[10];							inform_L[69][6] = l_cell_wire[11];							inform_L[6][6] = l_cell_wire[12];							inform_L[70][6] = l_cell_wire[13];							inform_L[7][6] = l_cell_wire[14];							inform_L[71][6] = l_cell_wire[15];							inform_L[8][6] = l_cell_wire[16];							inform_L[72][6] = l_cell_wire[17];							inform_L[9][6] = l_cell_wire[18];							inform_L[73][6] = l_cell_wire[19];							inform_L[10][6] = l_cell_wire[20];							inform_L[74][6] = l_cell_wire[21];							inform_L[11][6] = l_cell_wire[22];							inform_L[75][6] = l_cell_wire[23];							inform_L[12][6] = l_cell_wire[24];							inform_L[76][6] = l_cell_wire[25];							inform_L[13][6] = l_cell_wire[26];							inform_L[77][6] = l_cell_wire[27];							inform_L[14][6] = l_cell_wire[28];							inform_L[78][6] = l_cell_wire[29];							inform_L[15][6] = l_cell_wire[30];							inform_L[79][6] = l_cell_wire[31];							inform_L[16][6] = l_cell_wire[32];							inform_L[80][6] = l_cell_wire[33];							inform_L[17][6] = l_cell_wire[34];							inform_L[81][6] = l_cell_wire[35];							inform_L[18][6] = l_cell_wire[36];							inform_L[82][6] = l_cell_wire[37];							inform_L[19][6] = l_cell_wire[38];							inform_L[83][6] = l_cell_wire[39];							inform_L[20][6] = l_cell_wire[40];							inform_L[84][6] = l_cell_wire[41];							inform_L[21][6] = l_cell_wire[42];							inform_L[85][6] = l_cell_wire[43];							inform_L[22][6] = l_cell_wire[44];							inform_L[86][6] = l_cell_wire[45];							inform_L[23][6] = l_cell_wire[46];							inform_L[87][6] = l_cell_wire[47];							inform_L[24][6] = l_cell_wire[48];							inform_L[88][6] = l_cell_wire[49];							inform_L[25][6] = l_cell_wire[50];							inform_L[89][6] = l_cell_wire[51];							inform_L[26][6] = l_cell_wire[52];							inform_L[90][6] = l_cell_wire[53];							inform_L[27][6] = l_cell_wire[54];							inform_L[91][6] = l_cell_wire[55];							inform_L[28][6] = l_cell_wire[56];							inform_L[92][6] = l_cell_wire[57];							inform_L[29][6] = l_cell_wire[58];							inform_L[93][6] = l_cell_wire[59];							inform_L[30][6] = l_cell_wire[60];							inform_L[94][6] = l_cell_wire[61];							inform_L[31][6] = l_cell_wire[62];							inform_L[95][6] = l_cell_wire[63];							inform_L[32][6] = l_cell_wire[64];							inform_L[96][6] = l_cell_wire[65];							inform_L[33][6] = l_cell_wire[66];							inform_L[97][6] = l_cell_wire[67];							inform_L[34][6] = l_cell_wire[68];							inform_L[98][6] = l_cell_wire[69];							inform_L[35][6] = l_cell_wire[70];							inform_L[99][6] = l_cell_wire[71];							inform_L[36][6] = l_cell_wire[72];							inform_L[100][6] = l_cell_wire[73];							inform_L[37][6] = l_cell_wire[74];							inform_L[101][6] = l_cell_wire[75];							inform_L[38][6] = l_cell_wire[76];							inform_L[102][6] = l_cell_wire[77];							inform_L[39][6] = l_cell_wire[78];							inform_L[103][6] = l_cell_wire[79];							inform_L[40][6] = l_cell_wire[80];							inform_L[104][6] = l_cell_wire[81];							inform_L[41][6] = l_cell_wire[82];							inform_L[105][6] = l_cell_wire[83];							inform_L[42][6] = l_cell_wire[84];							inform_L[106][6] = l_cell_wire[85];							inform_L[43][6] = l_cell_wire[86];							inform_L[107][6] = l_cell_wire[87];							inform_L[44][6] = l_cell_wire[88];							inform_L[108][6] = l_cell_wire[89];							inform_L[45][6] = l_cell_wire[90];							inform_L[109][6] = l_cell_wire[91];							inform_L[46][6] = l_cell_wire[92];							inform_L[110][6] = l_cell_wire[93];							inform_L[47][6] = l_cell_wire[94];							inform_L[111][6] = l_cell_wire[95];							inform_L[48][6] = l_cell_wire[96];							inform_L[112][6] = l_cell_wire[97];							inform_L[49][6] = l_cell_wire[98];							inform_L[113][6] = l_cell_wire[99];							inform_L[50][6] = l_cell_wire[100];							inform_L[114][6] = l_cell_wire[101];							inform_L[51][6] = l_cell_wire[102];							inform_L[115][6] = l_cell_wire[103];							inform_L[52][6] = l_cell_wire[104];							inform_L[116][6] = l_cell_wire[105];							inform_L[53][6] = l_cell_wire[106];							inform_L[117][6] = l_cell_wire[107];							inform_L[54][6] = l_cell_wire[108];							inform_L[118][6] = l_cell_wire[109];							inform_L[55][6] = l_cell_wire[110];							inform_L[119][6] = l_cell_wire[111];							inform_L[56][6] = l_cell_wire[112];							inform_L[120][6] = l_cell_wire[113];							inform_L[57][6] = l_cell_wire[114];							inform_L[121][6] = l_cell_wire[115];							inform_L[58][6] = l_cell_wire[116];							inform_L[122][6] = l_cell_wire[117];							inform_L[59][6] = l_cell_wire[118];							inform_L[123][6] = l_cell_wire[119];							inform_L[60][6] = l_cell_wire[120];							inform_L[124][6] = l_cell_wire[121];							inform_L[61][6] = l_cell_wire[122];							inform_L[125][6] = l_cell_wire[123];							inform_L[62][6] = l_cell_wire[124];							inform_L[126][6] = l_cell_wire[125];							inform_L[63][6] = l_cell_wire[126];							inform_L[127][6] = l_cell_wire[127];							inform_L[128][6] = l_cell_wire[128];							inform_L[192][6] = l_cell_wire[129];							inform_L[129][6] = l_cell_wire[130];							inform_L[193][6] = l_cell_wire[131];							inform_L[130][6] = l_cell_wire[132];							inform_L[194][6] = l_cell_wire[133];							inform_L[131][6] = l_cell_wire[134];							inform_L[195][6] = l_cell_wire[135];							inform_L[132][6] = l_cell_wire[136];							inform_L[196][6] = l_cell_wire[137];							inform_L[133][6] = l_cell_wire[138];							inform_L[197][6] = l_cell_wire[139];							inform_L[134][6] = l_cell_wire[140];							inform_L[198][6] = l_cell_wire[141];							inform_L[135][6] = l_cell_wire[142];							inform_L[199][6] = l_cell_wire[143];							inform_L[136][6] = l_cell_wire[144];							inform_L[200][6] = l_cell_wire[145];							inform_L[137][6] = l_cell_wire[146];							inform_L[201][6] = l_cell_wire[147];							inform_L[138][6] = l_cell_wire[148];							inform_L[202][6] = l_cell_wire[149];							inform_L[139][6] = l_cell_wire[150];							inform_L[203][6] = l_cell_wire[151];							inform_L[140][6] = l_cell_wire[152];							inform_L[204][6] = l_cell_wire[153];							inform_L[141][6] = l_cell_wire[154];							inform_L[205][6] = l_cell_wire[155];							inform_L[142][6] = l_cell_wire[156];							inform_L[206][6] = l_cell_wire[157];							inform_L[143][6] = l_cell_wire[158];							inform_L[207][6] = l_cell_wire[159];							inform_L[144][6] = l_cell_wire[160];							inform_L[208][6] = l_cell_wire[161];							inform_L[145][6] = l_cell_wire[162];							inform_L[209][6] = l_cell_wire[163];							inform_L[146][6] = l_cell_wire[164];							inform_L[210][6] = l_cell_wire[165];							inform_L[147][6] = l_cell_wire[166];							inform_L[211][6] = l_cell_wire[167];							inform_L[148][6] = l_cell_wire[168];							inform_L[212][6] = l_cell_wire[169];							inform_L[149][6] = l_cell_wire[170];							inform_L[213][6] = l_cell_wire[171];							inform_L[150][6] = l_cell_wire[172];							inform_L[214][6] = l_cell_wire[173];							inform_L[151][6] = l_cell_wire[174];							inform_L[215][6] = l_cell_wire[175];							inform_L[152][6] = l_cell_wire[176];							inform_L[216][6] = l_cell_wire[177];							inform_L[153][6] = l_cell_wire[178];							inform_L[217][6] = l_cell_wire[179];							inform_L[154][6] = l_cell_wire[180];							inform_L[218][6] = l_cell_wire[181];							inform_L[155][6] = l_cell_wire[182];							inform_L[219][6] = l_cell_wire[183];							inform_L[156][6] = l_cell_wire[184];							inform_L[220][6] = l_cell_wire[185];							inform_L[157][6] = l_cell_wire[186];							inform_L[221][6] = l_cell_wire[187];							inform_L[158][6] = l_cell_wire[188];							inform_L[222][6] = l_cell_wire[189];							inform_L[159][6] = l_cell_wire[190];							inform_L[223][6] = l_cell_wire[191];							inform_L[160][6] = l_cell_wire[192];							inform_L[224][6] = l_cell_wire[193];							inform_L[161][6] = l_cell_wire[194];							inform_L[225][6] = l_cell_wire[195];							inform_L[162][6] = l_cell_wire[196];							inform_L[226][6] = l_cell_wire[197];							inform_L[163][6] = l_cell_wire[198];							inform_L[227][6] = l_cell_wire[199];							inform_L[164][6] = l_cell_wire[200];							inform_L[228][6] = l_cell_wire[201];							inform_L[165][6] = l_cell_wire[202];							inform_L[229][6] = l_cell_wire[203];							inform_L[166][6] = l_cell_wire[204];							inform_L[230][6] = l_cell_wire[205];							inform_L[167][6] = l_cell_wire[206];							inform_L[231][6] = l_cell_wire[207];							inform_L[168][6] = l_cell_wire[208];							inform_L[232][6] = l_cell_wire[209];							inform_L[169][6] = l_cell_wire[210];							inform_L[233][6] = l_cell_wire[211];							inform_L[170][6] = l_cell_wire[212];							inform_L[234][6] = l_cell_wire[213];							inform_L[171][6] = l_cell_wire[214];							inform_L[235][6] = l_cell_wire[215];							inform_L[172][6] = l_cell_wire[216];							inform_L[236][6] = l_cell_wire[217];							inform_L[173][6] = l_cell_wire[218];							inform_L[237][6] = l_cell_wire[219];							inform_L[174][6] = l_cell_wire[220];							inform_L[238][6] = l_cell_wire[221];							inform_L[175][6] = l_cell_wire[222];							inform_L[239][6] = l_cell_wire[223];							inform_L[176][6] = l_cell_wire[224];							inform_L[240][6] = l_cell_wire[225];							inform_L[177][6] = l_cell_wire[226];							inform_L[241][6] = l_cell_wire[227];							inform_L[178][6] = l_cell_wire[228];							inform_L[242][6] = l_cell_wire[229];							inform_L[179][6] = l_cell_wire[230];							inform_L[243][6] = l_cell_wire[231];							inform_L[180][6] = l_cell_wire[232];							inform_L[244][6] = l_cell_wire[233];							inform_L[181][6] = l_cell_wire[234];							inform_L[245][6] = l_cell_wire[235];							inform_L[182][6] = l_cell_wire[236];							inform_L[246][6] = l_cell_wire[237];							inform_L[183][6] = l_cell_wire[238];							inform_L[247][6] = l_cell_wire[239];							inform_L[184][6] = l_cell_wire[240];							inform_L[248][6] = l_cell_wire[241];							inform_L[185][6] = l_cell_wire[242];							inform_L[249][6] = l_cell_wire[243];							inform_L[186][6] = l_cell_wire[244];							inform_L[250][6] = l_cell_wire[245];							inform_L[187][6] = l_cell_wire[246];							inform_L[251][6] = l_cell_wire[247];							inform_L[188][6] = l_cell_wire[248];							inform_L[252][6] = l_cell_wire[249];							inform_L[189][6] = l_cell_wire[250];							inform_L[253][6] = l_cell_wire[251];							inform_L[190][6] = l_cell_wire[252];							inform_L[254][6] = l_cell_wire[253];							inform_L[191][6] = l_cell_wire[254];							inform_L[255][6] = l_cell_wire[255];						end
						8:						begin							inform_R[0][8] = r_cell_wire[0];							inform_R[128][8] = r_cell_wire[1];							inform_R[1][8] = r_cell_wire[2];							inform_R[129][8] = r_cell_wire[3];							inform_R[2][8] = r_cell_wire[4];							inform_R[130][8] = r_cell_wire[5];							inform_R[3][8] = r_cell_wire[6];							inform_R[131][8] = r_cell_wire[7];							inform_R[4][8] = r_cell_wire[8];							inform_R[132][8] = r_cell_wire[9];							inform_R[5][8] = r_cell_wire[10];							inform_R[133][8] = r_cell_wire[11];							inform_R[6][8] = r_cell_wire[12];							inform_R[134][8] = r_cell_wire[13];							inform_R[7][8] = r_cell_wire[14];							inform_R[135][8] = r_cell_wire[15];							inform_R[8][8] = r_cell_wire[16];							inform_R[136][8] = r_cell_wire[17];							inform_R[9][8] = r_cell_wire[18];							inform_R[137][8] = r_cell_wire[19];							inform_R[10][8] = r_cell_wire[20];							inform_R[138][8] = r_cell_wire[21];							inform_R[11][8] = r_cell_wire[22];							inform_R[139][8] = r_cell_wire[23];							inform_R[12][8] = r_cell_wire[24];							inform_R[140][8] = r_cell_wire[25];							inform_R[13][8] = r_cell_wire[26];							inform_R[141][8] = r_cell_wire[27];							inform_R[14][8] = r_cell_wire[28];							inform_R[142][8] = r_cell_wire[29];							inform_R[15][8] = r_cell_wire[30];							inform_R[143][8] = r_cell_wire[31];							inform_R[16][8] = r_cell_wire[32];							inform_R[144][8] = r_cell_wire[33];							inform_R[17][8] = r_cell_wire[34];							inform_R[145][8] = r_cell_wire[35];							inform_R[18][8] = r_cell_wire[36];							inform_R[146][8] = r_cell_wire[37];							inform_R[19][8] = r_cell_wire[38];							inform_R[147][8] = r_cell_wire[39];							inform_R[20][8] = r_cell_wire[40];							inform_R[148][8] = r_cell_wire[41];							inform_R[21][8] = r_cell_wire[42];							inform_R[149][8] = r_cell_wire[43];							inform_R[22][8] = r_cell_wire[44];							inform_R[150][8] = r_cell_wire[45];							inform_R[23][8] = r_cell_wire[46];							inform_R[151][8] = r_cell_wire[47];							inform_R[24][8] = r_cell_wire[48];							inform_R[152][8] = r_cell_wire[49];							inform_R[25][8] = r_cell_wire[50];							inform_R[153][8] = r_cell_wire[51];							inform_R[26][8] = r_cell_wire[52];							inform_R[154][8] = r_cell_wire[53];							inform_R[27][8] = r_cell_wire[54];							inform_R[155][8] = r_cell_wire[55];							inform_R[28][8] = r_cell_wire[56];							inform_R[156][8] = r_cell_wire[57];							inform_R[29][8] = r_cell_wire[58];							inform_R[157][8] = r_cell_wire[59];							inform_R[30][8] = r_cell_wire[60];							inform_R[158][8] = r_cell_wire[61];							inform_R[31][8] = r_cell_wire[62];							inform_R[159][8] = r_cell_wire[63];							inform_R[32][8] = r_cell_wire[64];							inform_R[160][8] = r_cell_wire[65];							inform_R[33][8] = r_cell_wire[66];							inform_R[161][8] = r_cell_wire[67];							inform_R[34][8] = r_cell_wire[68];							inform_R[162][8] = r_cell_wire[69];							inform_R[35][8] = r_cell_wire[70];							inform_R[163][8] = r_cell_wire[71];							inform_R[36][8] = r_cell_wire[72];							inform_R[164][8] = r_cell_wire[73];							inform_R[37][8] = r_cell_wire[74];							inform_R[165][8] = r_cell_wire[75];							inform_R[38][8] = r_cell_wire[76];							inform_R[166][8] = r_cell_wire[77];							inform_R[39][8] = r_cell_wire[78];							inform_R[167][8] = r_cell_wire[79];							inform_R[40][8] = r_cell_wire[80];							inform_R[168][8] = r_cell_wire[81];							inform_R[41][8] = r_cell_wire[82];							inform_R[169][8] = r_cell_wire[83];							inform_R[42][8] = r_cell_wire[84];							inform_R[170][8] = r_cell_wire[85];							inform_R[43][8] = r_cell_wire[86];							inform_R[171][8] = r_cell_wire[87];							inform_R[44][8] = r_cell_wire[88];							inform_R[172][8] = r_cell_wire[89];							inform_R[45][8] = r_cell_wire[90];							inform_R[173][8] = r_cell_wire[91];							inform_R[46][8] = r_cell_wire[92];							inform_R[174][8] = r_cell_wire[93];							inform_R[47][8] = r_cell_wire[94];							inform_R[175][8] = r_cell_wire[95];							inform_R[48][8] = r_cell_wire[96];							inform_R[176][8] = r_cell_wire[97];							inform_R[49][8] = r_cell_wire[98];							inform_R[177][8] = r_cell_wire[99];							inform_R[50][8] = r_cell_wire[100];							inform_R[178][8] = r_cell_wire[101];							inform_R[51][8] = r_cell_wire[102];							inform_R[179][8] = r_cell_wire[103];							inform_R[52][8] = r_cell_wire[104];							inform_R[180][8] = r_cell_wire[105];							inform_R[53][8] = r_cell_wire[106];							inform_R[181][8] = r_cell_wire[107];							inform_R[54][8] = r_cell_wire[108];							inform_R[182][8] = r_cell_wire[109];							inform_R[55][8] = r_cell_wire[110];							inform_R[183][8] = r_cell_wire[111];							inform_R[56][8] = r_cell_wire[112];							inform_R[184][8] = r_cell_wire[113];							inform_R[57][8] = r_cell_wire[114];							inform_R[185][8] = r_cell_wire[115];							inform_R[58][8] = r_cell_wire[116];							inform_R[186][8] = r_cell_wire[117];							inform_R[59][8] = r_cell_wire[118];							inform_R[187][8] = r_cell_wire[119];							inform_R[60][8] = r_cell_wire[120];							inform_R[188][8] = r_cell_wire[121];							inform_R[61][8] = r_cell_wire[122];							inform_R[189][8] = r_cell_wire[123];							inform_R[62][8] = r_cell_wire[124];							inform_R[190][8] = r_cell_wire[125];							inform_R[63][8] = r_cell_wire[126];							inform_R[191][8] = r_cell_wire[127];							inform_R[64][8] = r_cell_wire[128];							inform_R[192][8] = r_cell_wire[129];							inform_R[65][8] = r_cell_wire[130];							inform_R[193][8] = r_cell_wire[131];							inform_R[66][8] = r_cell_wire[132];							inform_R[194][8] = r_cell_wire[133];							inform_R[67][8] = r_cell_wire[134];							inform_R[195][8] = r_cell_wire[135];							inform_R[68][8] = r_cell_wire[136];							inform_R[196][8] = r_cell_wire[137];							inform_R[69][8] = r_cell_wire[138];							inform_R[197][8] = r_cell_wire[139];							inform_R[70][8] = r_cell_wire[140];							inform_R[198][8] = r_cell_wire[141];							inform_R[71][8] = r_cell_wire[142];							inform_R[199][8] = r_cell_wire[143];							inform_R[72][8] = r_cell_wire[144];							inform_R[200][8] = r_cell_wire[145];							inform_R[73][8] = r_cell_wire[146];							inform_R[201][8] = r_cell_wire[147];							inform_R[74][8] = r_cell_wire[148];							inform_R[202][8] = r_cell_wire[149];							inform_R[75][8] = r_cell_wire[150];							inform_R[203][8] = r_cell_wire[151];							inform_R[76][8] = r_cell_wire[152];							inform_R[204][8] = r_cell_wire[153];							inform_R[77][8] = r_cell_wire[154];							inform_R[205][8] = r_cell_wire[155];							inform_R[78][8] = r_cell_wire[156];							inform_R[206][8] = r_cell_wire[157];							inform_R[79][8] = r_cell_wire[158];							inform_R[207][8] = r_cell_wire[159];							inform_R[80][8] = r_cell_wire[160];							inform_R[208][8] = r_cell_wire[161];							inform_R[81][8] = r_cell_wire[162];							inform_R[209][8] = r_cell_wire[163];							inform_R[82][8] = r_cell_wire[164];							inform_R[210][8] = r_cell_wire[165];							inform_R[83][8] = r_cell_wire[166];							inform_R[211][8] = r_cell_wire[167];							inform_R[84][8] = r_cell_wire[168];							inform_R[212][8] = r_cell_wire[169];							inform_R[85][8] = r_cell_wire[170];							inform_R[213][8] = r_cell_wire[171];							inform_R[86][8] = r_cell_wire[172];							inform_R[214][8] = r_cell_wire[173];							inform_R[87][8] = r_cell_wire[174];							inform_R[215][8] = r_cell_wire[175];							inform_R[88][8] = r_cell_wire[176];							inform_R[216][8] = r_cell_wire[177];							inform_R[89][8] = r_cell_wire[178];							inform_R[217][8] = r_cell_wire[179];							inform_R[90][8] = r_cell_wire[180];							inform_R[218][8] = r_cell_wire[181];							inform_R[91][8] = r_cell_wire[182];							inform_R[219][8] = r_cell_wire[183];							inform_R[92][8] = r_cell_wire[184];							inform_R[220][8] = r_cell_wire[185];							inform_R[93][8] = r_cell_wire[186];							inform_R[221][8] = r_cell_wire[187];							inform_R[94][8] = r_cell_wire[188];							inform_R[222][8] = r_cell_wire[189];							inform_R[95][8] = r_cell_wire[190];							inform_R[223][8] = r_cell_wire[191];							inform_R[96][8] = r_cell_wire[192];							inform_R[224][8] = r_cell_wire[193];							inform_R[97][8] = r_cell_wire[194];							inform_R[225][8] = r_cell_wire[195];							inform_R[98][8] = r_cell_wire[196];							inform_R[226][8] = r_cell_wire[197];							inform_R[99][8] = r_cell_wire[198];							inform_R[227][8] = r_cell_wire[199];							inform_R[100][8] = r_cell_wire[200];							inform_R[228][8] = r_cell_wire[201];							inform_R[101][8] = r_cell_wire[202];							inform_R[229][8] = r_cell_wire[203];							inform_R[102][8] = r_cell_wire[204];							inform_R[230][8] = r_cell_wire[205];							inform_R[103][8] = r_cell_wire[206];							inform_R[231][8] = r_cell_wire[207];							inform_R[104][8] = r_cell_wire[208];							inform_R[232][8] = r_cell_wire[209];							inform_R[105][8] = r_cell_wire[210];							inform_R[233][8] = r_cell_wire[211];							inform_R[106][8] = r_cell_wire[212];							inform_R[234][8] = r_cell_wire[213];							inform_R[107][8] = r_cell_wire[214];							inform_R[235][8] = r_cell_wire[215];							inform_R[108][8] = r_cell_wire[216];							inform_R[236][8] = r_cell_wire[217];							inform_R[109][8] = r_cell_wire[218];							inform_R[237][8] = r_cell_wire[219];							inform_R[110][8] = r_cell_wire[220];							inform_R[238][8] = r_cell_wire[221];							inform_R[111][8] = r_cell_wire[222];							inform_R[239][8] = r_cell_wire[223];							inform_R[112][8] = r_cell_wire[224];							inform_R[240][8] = r_cell_wire[225];							inform_R[113][8] = r_cell_wire[226];							inform_R[241][8] = r_cell_wire[227];							inform_R[114][8] = r_cell_wire[228];							inform_R[242][8] = r_cell_wire[229];							inform_R[115][8] = r_cell_wire[230];							inform_R[243][8] = r_cell_wire[231];							inform_R[116][8] = r_cell_wire[232];							inform_R[244][8] = r_cell_wire[233];							inform_R[117][8] = r_cell_wire[234];							inform_R[245][8] = r_cell_wire[235];							inform_R[118][8] = r_cell_wire[236];							inform_R[246][8] = r_cell_wire[237];							inform_R[119][8] = r_cell_wire[238];							inform_R[247][8] = r_cell_wire[239];							inform_R[120][8] = r_cell_wire[240];							inform_R[248][8] = r_cell_wire[241];							inform_R[121][8] = r_cell_wire[242];							inform_R[249][8] = r_cell_wire[243];							inform_R[122][8] = r_cell_wire[244];							inform_R[250][8] = r_cell_wire[245];							inform_R[123][8] = r_cell_wire[246];							inform_R[251][8] = r_cell_wire[247];							inform_R[124][8] = r_cell_wire[248];							inform_R[252][8] = r_cell_wire[249];							inform_R[125][8] = r_cell_wire[250];							inform_R[253][8] = r_cell_wire[251];							inform_R[126][8] = r_cell_wire[252];							inform_R[254][8] = r_cell_wire[253];							inform_R[127][8] = r_cell_wire[254];							inform_R[255][8] = r_cell_wire[255];							inform_L[0][7] = l_cell_wire[0];							inform_L[128][7] = l_cell_wire[1];							inform_L[1][7] = l_cell_wire[2];							inform_L[129][7] = l_cell_wire[3];							inform_L[2][7] = l_cell_wire[4];							inform_L[130][7] = l_cell_wire[5];							inform_L[3][7] = l_cell_wire[6];							inform_L[131][7] = l_cell_wire[7];							inform_L[4][7] = l_cell_wire[8];							inform_L[132][7] = l_cell_wire[9];							inform_L[5][7] = l_cell_wire[10];							inform_L[133][7] = l_cell_wire[11];							inform_L[6][7] = l_cell_wire[12];							inform_L[134][7] = l_cell_wire[13];							inform_L[7][7] = l_cell_wire[14];							inform_L[135][7] = l_cell_wire[15];							inform_L[8][7] = l_cell_wire[16];							inform_L[136][7] = l_cell_wire[17];							inform_L[9][7] = l_cell_wire[18];							inform_L[137][7] = l_cell_wire[19];							inform_L[10][7] = l_cell_wire[20];							inform_L[138][7] = l_cell_wire[21];							inform_L[11][7] = l_cell_wire[22];							inform_L[139][7] = l_cell_wire[23];							inform_L[12][7] = l_cell_wire[24];							inform_L[140][7] = l_cell_wire[25];							inform_L[13][7] = l_cell_wire[26];							inform_L[141][7] = l_cell_wire[27];							inform_L[14][7] = l_cell_wire[28];							inform_L[142][7] = l_cell_wire[29];							inform_L[15][7] = l_cell_wire[30];							inform_L[143][7] = l_cell_wire[31];							inform_L[16][7] = l_cell_wire[32];							inform_L[144][7] = l_cell_wire[33];							inform_L[17][7] = l_cell_wire[34];							inform_L[145][7] = l_cell_wire[35];							inform_L[18][7] = l_cell_wire[36];							inform_L[146][7] = l_cell_wire[37];							inform_L[19][7] = l_cell_wire[38];							inform_L[147][7] = l_cell_wire[39];							inform_L[20][7] = l_cell_wire[40];							inform_L[148][7] = l_cell_wire[41];							inform_L[21][7] = l_cell_wire[42];							inform_L[149][7] = l_cell_wire[43];							inform_L[22][7] = l_cell_wire[44];							inform_L[150][7] = l_cell_wire[45];							inform_L[23][7] = l_cell_wire[46];							inform_L[151][7] = l_cell_wire[47];							inform_L[24][7] = l_cell_wire[48];							inform_L[152][7] = l_cell_wire[49];							inform_L[25][7] = l_cell_wire[50];							inform_L[153][7] = l_cell_wire[51];							inform_L[26][7] = l_cell_wire[52];							inform_L[154][7] = l_cell_wire[53];							inform_L[27][7] = l_cell_wire[54];							inform_L[155][7] = l_cell_wire[55];							inform_L[28][7] = l_cell_wire[56];							inform_L[156][7] = l_cell_wire[57];							inform_L[29][7] = l_cell_wire[58];							inform_L[157][7] = l_cell_wire[59];							inform_L[30][7] = l_cell_wire[60];							inform_L[158][7] = l_cell_wire[61];							inform_L[31][7] = l_cell_wire[62];							inform_L[159][7] = l_cell_wire[63];							inform_L[32][7] = l_cell_wire[64];							inform_L[160][7] = l_cell_wire[65];							inform_L[33][7] = l_cell_wire[66];							inform_L[161][7] = l_cell_wire[67];							inform_L[34][7] = l_cell_wire[68];							inform_L[162][7] = l_cell_wire[69];							inform_L[35][7] = l_cell_wire[70];							inform_L[163][7] = l_cell_wire[71];							inform_L[36][7] = l_cell_wire[72];							inform_L[164][7] = l_cell_wire[73];							inform_L[37][7] = l_cell_wire[74];							inform_L[165][7] = l_cell_wire[75];							inform_L[38][7] = l_cell_wire[76];							inform_L[166][7] = l_cell_wire[77];							inform_L[39][7] = l_cell_wire[78];							inform_L[167][7] = l_cell_wire[79];							inform_L[40][7] = l_cell_wire[80];							inform_L[168][7] = l_cell_wire[81];							inform_L[41][7] = l_cell_wire[82];							inform_L[169][7] = l_cell_wire[83];							inform_L[42][7] = l_cell_wire[84];							inform_L[170][7] = l_cell_wire[85];							inform_L[43][7] = l_cell_wire[86];							inform_L[171][7] = l_cell_wire[87];							inform_L[44][7] = l_cell_wire[88];							inform_L[172][7] = l_cell_wire[89];							inform_L[45][7] = l_cell_wire[90];							inform_L[173][7] = l_cell_wire[91];							inform_L[46][7] = l_cell_wire[92];							inform_L[174][7] = l_cell_wire[93];							inform_L[47][7] = l_cell_wire[94];							inform_L[175][7] = l_cell_wire[95];							inform_L[48][7] = l_cell_wire[96];							inform_L[176][7] = l_cell_wire[97];							inform_L[49][7] = l_cell_wire[98];							inform_L[177][7] = l_cell_wire[99];							inform_L[50][7] = l_cell_wire[100];							inform_L[178][7] = l_cell_wire[101];							inform_L[51][7] = l_cell_wire[102];							inform_L[179][7] = l_cell_wire[103];							inform_L[52][7] = l_cell_wire[104];							inform_L[180][7] = l_cell_wire[105];							inform_L[53][7] = l_cell_wire[106];							inform_L[181][7] = l_cell_wire[107];							inform_L[54][7] = l_cell_wire[108];							inform_L[182][7] = l_cell_wire[109];							inform_L[55][7] = l_cell_wire[110];							inform_L[183][7] = l_cell_wire[111];							inform_L[56][7] = l_cell_wire[112];							inform_L[184][7] = l_cell_wire[113];							inform_L[57][7] = l_cell_wire[114];							inform_L[185][7] = l_cell_wire[115];							inform_L[58][7] = l_cell_wire[116];							inform_L[186][7] = l_cell_wire[117];							inform_L[59][7] = l_cell_wire[118];							inform_L[187][7] = l_cell_wire[119];							inform_L[60][7] = l_cell_wire[120];							inform_L[188][7] = l_cell_wire[121];							inform_L[61][7] = l_cell_wire[122];							inform_L[189][7] = l_cell_wire[123];							inform_L[62][7] = l_cell_wire[124];							inform_L[190][7] = l_cell_wire[125];							inform_L[63][7] = l_cell_wire[126];							inform_L[191][7] = l_cell_wire[127];							inform_L[64][7] = l_cell_wire[128];							inform_L[192][7] = l_cell_wire[129];							inform_L[65][7] = l_cell_wire[130];							inform_L[193][7] = l_cell_wire[131];							inform_L[66][7] = l_cell_wire[132];							inform_L[194][7] = l_cell_wire[133];							inform_L[67][7] = l_cell_wire[134];							inform_L[195][7] = l_cell_wire[135];							inform_L[68][7] = l_cell_wire[136];							inform_L[196][7] = l_cell_wire[137];							inform_L[69][7] = l_cell_wire[138];							inform_L[197][7] = l_cell_wire[139];							inform_L[70][7] = l_cell_wire[140];							inform_L[198][7] = l_cell_wire[141];							inform_L[71][7] = l_cell_wire[142];							inform_L[199][7] = l_cell_wire[143];							inform_L[72][7] = l_cell_wire[144];							inform_L[200][7] = l_cell_wire[145];							inform_L[73][7] = l_cell_wire[146];							inform_L[201][7] = l_cell_wire[147];							inform_L[74][7] = l_cell_wire[148];							inform_L[202][7] = l_cell_wire[149];							inform_L[75][7] = l_cell_wire[150];							inform_L[203][7] = l_cell_wire[151];							inform_L[76][7] = l_cell_wire[152];							inform_L[204][7] = l_cell_wire[153];							inform_L[77][7] = l_cell_wire[154];							inform_L[205][7] = l_cell_wire[155];							inform_L[78][7] = l_cell_wire[156];							inform_L[206][7] = l_cell_wire[157];							inform_L[79][7] = l_cell_wire[158];							inform_L[207][7] = l_cell_wire[159];							inform_L[80][7] = l_cell_wire[160];							inform_L[208][7] = l_cell_wire[161];							inform_L[81][7] = l_cell_wire[162];							inform_L[209][7] = l_cell_wire[163];							inform_L[82][7] = l_cell_wire[164];							inform_L[210][7] = l_cell_wire[165];							inform_L[83][7] = l_cell_wire[166];							inform_L[211][7] = l_cell_wire[167];							inform_L[84][7] = l_cell_wire[168];							inform_L[212][7] = l_cell_wire[169];							inform_L[85][7] = l_cell_wire[170];							inform_L[213][7] = l_cell_wire[171];							inform_L[86][7] = l_cell_wire[172];							inform_L[214][7] = l_cell_wire[173];							inform_L[87][7] = l_cell_wire[174];							inform_L[215][7] = l_cell_wire[175];							inform_L[88][7] = l_cell_wire[176];							inform_L[216][7] = l_cell_wire[177];							inform_L[89][7] = l_cell_wire[178];							inform_L[217][7] = l_cell_wire[179];							inform_L[90][7] = l_cell_wire[180];							inform_L[218][7] = l_cell_wire[181];							inform_L[91][7] = l_cell_wire[182];							inform_L[219][7] = l_cell_wire[183];							inform_L[92][7] = l_cell_wire[184];							inform_L[220][7] = l_cell_wire[185];							inform_L[93][7] = l_cell_wire[186];							inform_L[221][7] = l_cell_wire[187];							inform_L[94][7] = l_cell_wire[188];							inform_L[222][7] = l_cell_wire[189];							inform_L[95][7] = l_cell_wire[190];							inform_L[223][7] = l_cell_wire[191];							inform_L[96][7] = l_cell_wire[192];							inform_L[224][7] = l_cell_wire[193];							inform_L[97][7] = l_cell_wire[194];							inform_L[225][7] = l_cell_wire[195];							inform_L[98][7] = l_cell_wire[196];							inform_L[226][7] = l_cell_wire[197];							inform_L[99][7] = l_cell_wire[198];							inform_L[227][7] = l_cell_wire[199];							inform_L[100][7] = l_cell_wire[200];							inform_L[228][7] = l_cell_wire[201];							inform_L[101][7] = l_cell_wire[202];							inform_L[229][7] = l_cell_wire[203];							inform_L[102][7] = l_cell_wire[204];							inform_L[230][7] = l_cell_wire[205];							inform_L[103][7] = l_cell_wire[206];							inform_L[231][7] = l_cell_wire[207];							inform_L[104][7] = l_cell_wire[208];							inform_L[232][7] = l_cell_wire[209];							inform_L[105][7] = l_cell_wire[210];							inform_L[233][7] = l_cell_wire[211];							inform_L[106][7] = l_cell_wire[212];							inform_L[234][7] = l_cell_wire[213];							inform_L[107][7] = l_cell_wire[214];							inform_L[235][7] = l_cell_wire[215];							inform_L[108][7] = l_cell_wire[216];							inform_L[236][7] = l_cell_wire[217];							inform_L[109][7] = l_cell_wire[218];							inform_L[237][7] = l_cell_wire[219];							inform_L[110][7] = l_cell_wire[220];							inform_L[238][7] = l_cell_wire[221];							inform_L[111][7] = l_cell_wire[222];							inform_L[239][7] = l_cell_wire[223];							inform_L[112][7] = l_cell_wire[224];							inform_L[240][7] = l_cell_wire[225];							inform_L[113][7] = l_cell_wire[226];							inform_L[241][7] = l_cell_wire[227];							inform_L[114][7] = l_cell_wire[228];							inform_L[242][7] = l_cell_wire[229];							inform_L[115][7] = l_cell_wire[230];							inform_L[243][7] = l_cell_wire[231];							inform_L[116][7] = l_cell_wire[232];							inform_L[244][7] = l_cell_wire[233];							inform_L[117][7] = l_cell_wire[234];							inform_L[245][7] = l_cell_wire[235];							inform_L[118][7] = l_cell_wire[236];							inform_L[246][7] = l_cell_wire[237];							inform_L[119][7] = l_cell_wire[238];							inform_L[247][7] = l_cell_wire[239];							inform_L[120][7] = l_cell_wire[240];							inform_L[248][7] = l_cell_wire[241];							inform_L[121][7] = l_cell_wire[242];							inform_L[249][7] = l_cell_wire[243];							inform_L[122][7] = l_cell_wire[244];							inform_L[250][7] = l_cell_wire[245];							inform_L[123][7] = l_cell_wire[246];							inform_L[251][7] = l_cell_wire[247];							inform_L[124][7] = l_cell_wire[248];							inform_L[252][7] = l_cell_wire[249];							inform_L[125][7] = l_cell_wire[250];							inform_L[253][7] = l_cell_wire[251];							inform_L[126][7] = l_cell_wire[252];							inform_L[254][7] = l_cell_wire[253];							inform_L[127][7] = l_cell_wire[254];							inform_L[255][7] = l_cell_wire[255];						end
						default:							for (x = 0; x < 256; x = x + 1)								for (y = 0; y < 8; y = y + 1)								begin									inform_R[x][y+1] <= 8'd0;									inform_L[x][y] <= 8'd0;								end					endcase				end			end
			BUSY_RIGHT:			begin				if(clk_counter == 2'b11)begin					case (w2r)						1:						begin							inform_R[0][1] = r_cell_wire[0];							inform_R[1][1] = r_cell_wire[1];							inform_R[2][1] = r_cell_wire[2];							inform_R[3][1] = r_cell_wire[3];							inform_R[4][1] = r_cell_wire[4];							inform_R[5][1] = r_cell_wire[5];							inform_R[6][1] = r_cell_wire[6];							inform_R[7][1] = r_cell_wire[7];							inform_R[8][1] = r_cell_wire[8];							inform_R[9][1] = r_cell_wire[9];							inform_R[10][1] = r_cell_wire[10];							inform_R[11][1] = r_cell_wire[11];							inform_R[12][1] = r_cell_wire[12];							inform_R[13][1] = r_cell_wire[13];							inform_R[14][1] = r_cell_wire[14];							inform_R[15][1] = r_cell_wire[15];							inform_R[16][1] = r_cell_wire[16];							inform_R[17][1] = r_cell_wire[17];							inform_R[18][1] = r_cell_wire[18];							inform_R[19][1] = r_cell_wire[19];							inform_R[20][1] = r_cell_wire[20];							inform_R[21][1] = r_cell_wire[21];							inform_R[22][1] = r_cell_wire[22];							inform_R[23][1] = r_cell_wire[23];							inform_R[24][1] = r_cell_wire[24];							inform_R[25][1] = r_cell_wire[25];							inform_R[26][1] = r_cell_wire[26];							inform_R[27][1] = r_cell_wire[27];							inform_R[28][1] = r_cell_wire[28];							inform_R[29][1] = r_cell_wire[29];							inform_R[30][1] = r_cell_wire[30];							inform_R[31][1] = r_cell_wire[31];							inform_R[32][1] = r_cell_wire[32];							inform_R[33][1] = r_cell_wire[33];							inform_R[34][1] = r_cell_wire[34];							inform_R[35][1] = r_cell_wire[35];							inform_R[36][1] = r_cell_wire[36];							inform_R[37][1] = r_cell_wire[37];							inform_R[38][1] = r_cell_wire[38];							inform_R[39][1] = r_cell_wire[39];							inform_R[40][1] = r_cell_wire[40];							inform_R[41][1] = r_cell_wire[41];							inform_R[42][1] = r_cell_wire[42];							inform_R[43][1] = r_cell_wire[43];							inform_R[44][1] = r_cell_wire[44];							inform_R[45][1] = r_cell_wire[45];							inform_R[46][1] = r_cell_wire[46];							inform_R[47][1] = r_cell_wire[47];							inform_R[48][1] = r_cell_wire[48];							inform_R[49][1] = r_cell_wire[49];							inform_R[50][1] = r_cell_wire[50];							inform_R[51][1] = r_cell_wire[51];							inform_R[52][1] = r_cell_wire[52];							inform_R[53][1] = r_cell_wire[53];							inform_R[54][1] = r_cell_wire[54];							inform_R[55][1] = r_cell_wire[55];							inform_R[56][1] = r_cell_wire[56];							inform_R[57][1] = r_cell_wire[57];							inform_R[58][1] = r_cell_wire[58];							inform_R[59][1] = r_cell_wire[59];							inform_R[60][1] = r_cell_wire[60];							inform_R[61][1] = r_cell_wire[61];							inform_R[62][1] = r_cell_wire[62];							inform_R[63][1] = r_cell_wire[63];							inform_R[64][1] = r_cell_wire[64];							inform_R[65][1] = r_cell_wire[65];							inform_R[66][1] = r_cell_wire[66];							inform_R[67][1] = r_cell_wire[67];							inform_R[68][1] = r_cell_wire[68];							inform_R[69][1] = r_cell_wire[69];							inform_R[70][1] = r_cell_wire[70];							inform_R[71][1] = r_cell_wire[71];							inform_R[72][1] = r_cell_wire[72];							inform_R[73][1] = r_cell_wire[73];							inform_R[74][1] = r_cell_wire[74];							inform_R[75][1] = r_cell_wire[75];							inform_R[76][1] = r_cell_wire[76];							inform_R[77][1] = r_cell_wire[77];							inform_R[78][1] = r_cell_wire[78];							inform_R[79][1] = r_cell_wire[79];							inform_R[80][1] = r_cell_wire[80];							inform_R[81][1] = r_cell_wire[81];							inform_R[82][1] = r_cell_wire[82];							inform_R[83][1] = r_cell_wire[83];							inform_R[84][1] = r_cell_wire[84];							inform_R[85][1] = r_cell_wire[85];							inform_R[86][1] = r_cell_wire[86];							inform_R[87][1] = r_cell_wire[87];							inform_R[88][1] = r_cell_wire[88];							inform_R[89][1] = r_cell_wire[89];							inform_R[90][1] = r_cell_wire[90];							inform_R[91][1] = r_cell_wire[91];							inform_R[92][1] = r_cell_wire[92];							inform_R[93][1] = r_cell_wire[93];							inform_R[94][1] = r_cell_wire[94];							inform_R[95][1] = r_cell_wire[95];							inform_R[96][1] = r_cell_wire[96];							inform_R[97][1] = r_cell_wire[97];							inform_R[98][1] = r_cell_wire[98];							inform_R[99][1] = r_cell_wire[99];							inform_R[100][1] = r_cell_wire[100];							inform_R[101][1] = r_cell_wire[101];							inform_R[102][1] = r_cell_wire[102];							inform_R[103][1] = r_cell_wire[103];							inform_R[104][1] = r_cell_wire[104];							inform_R[105][1] = r_cell_wire[105];							inform_R[106][1] = r_cell_wire[106];							inform_R[107][1] = r_cell_wire[107];							inform_R[108][1] = r_cell_wire[108];							inform_R[109][1] = r_cell_wire[109];							inform_R[110][1] = r_cell_wire[110];							inform_R[111][1] = r_cell_wire[111];							inform_R[112][1] = r_cell_wire[112];							inform_R[113][1] = r_cell_wire[113];							inform_R[114][1] = r_cell_wire[114];							inform_R[115][1] = r_cell_wire[115];							inform_R[116][1] = r_cell_wire[116];							inform_R[117][1] = r_cell_wire[117];							inform_R[118][1] = r_cell_wire[118];							inform_R[119][1] = r_cell_wire[119];							inform_R[120][1] = r_cell_wire[120];							inform_R[121][1] = r_cell_wire[121];							inform_R[122][1] = r_cell_wire[122];							inform_R[123][1] = r_cell_wire[123];							inform_R[124][1] = r_cell_wire[124];							inform_R[125][1] = r_cell_wire[125];							inform_R[126][1] = r_cell_wire[126];							inform_R[127][1] = r_cell_wire[127];							inform_R[128][1] = r_cell_wire[128];							inform_R[129][1] = r_cell_wire[129];							inform_R[130][1] = r_cell_wire[130];							inform_R[131][1] = r_cell_wire[131];							inform_R[132][1] = r_cell_wire[132];							inform_R[133][1] = r_cell_wire[133];							inform_R[134][1] = r_cell_wire[134];							inform_R[135][1] = r_cell_wire[135];							inform_R[136][1] = r_cell_wire[136];							inform_R[137][1] = r_cell_wire[137];							inform_R[138][1] = r_cell_wire[138];							inform_R[139][1] = r_cell_wire[139];							inform_R[140][1] = r_cell_wire[140];							inform_R[141][1] = r_cell_wire[141];							inform_R[142][1] = r_cell_wire[142];							inform_R[143][1] = r_cell_wire[143];							inform_R[144][1] = r_cell_wire[144];							inform_R[145][1] = r_cell_wire[145];							inform_R[146][1] = r_cell_wire[146];							inform_R[147][1] = r_cell_wire[147];							inform_R[148][1] = r_cell_wire[148];							inform_R[149][1] = r_cell_wire[149];							inform_R[150][1] = r_cell_wire[150];							inform_R[151][1] = r_cell_wire[151];							inform_R[152][1] = r_cell_wire[152];							inform_R[153][1] = r_cell_wire[153];							inform_R[154][1] = r_cell_wire[154];							inform_R[155][1] = r_cell_wire[155];							inform_R[156][1] = r_cell_wire[156];							inform_R[157][1] = r_cell_wire[157];							inform_R[158][1] = r_cell_wire[158];							inform_R[159][1] = r_cell_wire[159];							inform_R[160][1] = r_cell_wire[160];							inform_R[161][1] = r_cell_wire[161];							inform_R[162][1] = r_cell_wire[162];							inform_R[163][1] = r_cell_wire[163];							inform_R[164][1] = r_cell_wire[164];							inform_R[165][1] = r_cell_wire[165];							inform_R[166][1] = r_cell_wire[166];							inform_R[167][1] = r_cell_wire[167];							inform_R[168][1] = r_cell_wire[168];							inform_R[169][1] = r_cell_wire[169];							inform_R[170][1] = r_cell_wire[170];							inform_R[171][1] = r_cell_wire[171];							inform_R[172][1] = r_cell_wire[172];							inform_R[173][1] = r_cell_wire[173];							inform_R[174][1] = r_cell_wire[174];							inform_R[175][1] = r_cell_wire[175];							inform_R[176][1] = r_cell_wire[176];							inform_R[177][1] = r_cell_wire[177];							inform_R[178][1] = r_cell_wire[178];							inform_R[179][1] = r_cell_wire[179];							inform_R[180][1] = r_cell_wire[180];							inform_R[181][1] = r_cell_wire[181];							inform_R[182][1] = r_cell_wire[182];							inform_R[183][1] = r_cell_wire[183];							inform_R[184][1] = r_cell_wire[184];							inform_R[185][1] = r_cell_wire[185];							inform_R[186][1] = r_cell_wire[186];							inform_R[187][1] = r_cell_wire[187];							inform_R[188][1] = r_cell_wire[188];							inform_R[189][1] = r_cell_wire[189];							inform_R[190][1] = r_cell_wire[190];							inform_R[191][1] = r_cell_wire[191];							inform_R[192][1] = r_cell_wire[192];							inform_R[193][1] = r_cell_wire[193];							inform_R[194][1] = r_cell_wire[194];							inform_R[195][1] = r_cell_wire[195];							inform_R[196][1] = r_cell_wire[196];							inform_R[197][1] = r_cell_wire[197];							inform_R[198][1] = r_cell_wire[198];							inform_R[199][1] = r_cell_wire[199];							inform_R[200][1] = r_cell_wire[200];							inform_R[201][1] = r_cell_wire[201];							inform_R[202][1] = r_cell_wire[202];							inform_R[203][1] = r_cell_wire[203];							inform_R[204][1] = r_cell_wire[204];							inform_R[205][1] = r_cell_wire[205];							inform_R[206][1] = r_cell_wire[206];							inform_R[207][1] = r_cell_wire[207];							inform_R[208][1] = r_cell_wire[208];							inform_R[209][1] = r_cell_wire[209];							inform_R[210][1] = r_cell_wire[210];							inform_R[211][1] = r_cell_wire[211];							inform_R[212][1] = r_cell_wire[212];							inform_R[213][1] = r_cell_wire[213];							inform_R[214][1] = r_cell_wire[214];							inform_R[215][1] = r_cell_wire[215];							inform_R[216][1] = r_cell_wire[216];							inform_R[217][1] = r_cell_wire[217];							inform_R[218][1] = r_cell_wire[218];							inform_R[219][1] = r_cell_wire[219];							inform_R[220][1] = r_cell_wire[220];							inform_R[221][1] = r_cell_wire[221];							inform_R[222][1] = r_cell_wire[222];							inform_R[223][1] = r_cell_wire[223];							inform_R[224][1] = r_cell_wire[224];							inform_R[225][1] = r_cell_wire[225];							inform_R[226][1] = r_cell_wire[226];							inform_R[227][1] = r_cell_wire[227];							inform_R[228][1] = r_cell_wire[228];							inform_R[229][1] = r_cell_wire[229];							inform_R[230][1] = r_cell_wire[230];							inform_R[231][1] = r_cell_wire[231];							inform_R[232][1] = r_cell_wire[232];							inform_R[233][1] = r_cell_wire[233];							inform_R[234][1] = r_cell_wire[234];							inform_R[235][1] = r_cell_wire[235];							inform_R[236][1] = r_cell_wire[236];							inform_R[237][1] = r_cell_wire[237];							inform_R[238][1] = r_cell_wire[238];							inform_R[239][1] = r_cell_wire[239];							inform_R[240][1] = r_cell_wire[240];							inform_R[241][1] = r_cell_wire[241];							inform_R[242][1] = r_cell_wire[242];							inform_R[243][1] = r_cell_wire[243];							inform_R[244][1] = r_cell_wire[244];							inform_R[245][1] = r_cell_wire[245];							inform_R[246][1] = r_cell_wire[246];							inform_R[247][1] = r_cell_wire[247];							inform_R[248][1] = r_cell_wire[248];							inform_R[249][1] = r_cell_wire[249];							inform_R[250][1] = r_cell_wire[250];							inform_R[251][1] = r_cell_wire[251];							inform_R[252][1] = r_cell_wire[252];							inform_R[253][1] = r_cell_wire[253];							inform_R[254][1] = r_cell_wire[254];							inform_R[255][1] = r_cell_wire[255];							inform_L[0][0] = l_cell_wire[0];							inform_L[1][0] = l_cell_wire[1];							inform_L[2][0] = l_cell_wire[2];							inform_L[3][0] = l_cell_wire[3];							inform_L[4][0] = l_cell_wire[4];							inform_L[5][0] = l_cell_wire[5];							inform_L[6][0] = l_cell_wire[6];							inform_L[7][0] = l_cell_wire[7];							inform_L[8][0] = l_cell_wire[8];							inform_L[9][0] = l_cell_wire[9];							inform_L[10][0] = l_cell_wire[10];							inform_L[11][0] = l_cell_wire[11];							inform_L[12][0] = l_cell_wire[12];							inform_L[13][0] = l_cell_wire[13];							inform_L[14][0] = l_cell_wire[14];							inform_L[15][0] = l_cell_wire[15];							inform_L[16][0] = l_cell_wire[16];							inform_L[17][0] = l_cell_wire[17];							inform_L[18][0] = l_cell_wire[18];							inform_L[19][0] = l_cell_wire[19];							inform_L[20][0] = l_cell_wire[20];							inform_L[21][0] = l_cell_wire[21];							inform_L[22][0] = l_cell_wire[22];							inform_L[23][0] = l_cell_wire[23];							inform_L[24][0] = l_cell_wire[24];							inform_L[25][0] = l_cell_wire[25];							inform_L[26][0] = l_cell_wire[26];							inform_L[27][0] = l_cell_wire[27];							inform_L[28][0] = l_cell_wire[28];							inform_L[29][0] = l_cell_wire[29];							inform_L[30][0] = l_cell_wire[30];							inform_L[31][0] = l_cell_wire[31];							inform_L[32][0] = l_cell_wire[32];							inform_L[33][0] = l_cell_wire[33];							inform_L[34][0] = l_cell_wire[34];							inform_L[35][0] = l_cell_wire[35];							inform_L[36][0] = l_cell_wire[36];							inform_L[37][0] = l_cell_wire[37];							inform_L[38][0] = l_cell_wire[38];							inform_L[39][0] = l_cell_wire[39];							inform_L[40][0] = l_cell_wire[40];							inform_L[41][0] = l_cell_wire[41];							inform_L[42][0] = l_cell_wire[42];							inform_L[43][0] = l_cell_wire[43];							inform_L[44][0] = l_cell_wire[44];							inform_L[45][0] = l_cell_wire[45];							inform_L[46][0] = l_cell_wire[46];							inform_L[47][0] = l_cell_wire[47];							inform_L[48][0] = l_cell_wire[48];							inform_L[49][0] = l_cell_wire[49];							inform_L[50][0] = l_cell_wire[50];							inform_L[51][0] = l_cell_wire[51];							inform_L[52][0] = l_cell_wire[52];							inform_L[53][0] = l_cell_wire[53];							inform_L[54][0] = l_cell_wire[54];							inform_L[55][0] = l_cell_wire[55];							inform_L[56][0] = l_cell_wire[56];							inform_L[57][0] = l_cell_wire[57];							inform_L[58][0] = l_cell_wire[58];							inform_L[59][0] = l_cell_wire[59];							inform_L[60][0] = l_cell_wire[60];							inform_L[61][0] = l_cell_wire[61];							inform_L[62][0] = l_cell_wire[62];							inform_L[63][0] = l_cell_wire[63];							inform_L[64][0] = l_cell_wire[64];							inform_L[65][0] = l_cell_wire[65];							inform_L[66][0] = l_cell_wire[66];							inform_L[67][0] = l_cell_wire[67];							inform_L[68][0] = l_cell_wire[68];							inform_L[69][0] = l_cell_wire[69];							inform_L[70][0] = l_cell_wire[70];							inform_L[71][0] = l_cell_wire[71];							inform_L[72][0] = l_cell_wire[72];							inform_L[73][0] = l_cell_wire[73];							inform_L[74][0] = l_cell_wire[74];							inform_L[75][0] = l_cell_wire[75];							inform_L[76][0] = l_cell_wire[76];							inform_L[77][0] = l_cell_wire[77];							inform_L[78][0] = l_cell_wire[78];							inform_L[79][0] = l_cell_wire[79];							inform_L[80][0] = l_cell_wire[80];							inform_L[81][0] = l_cell_wire[81];							inform_L[82][0] = l_cell_wire[82];							inform_L[83][0] = l_cell_wire[83];							inform_L[84][0] = l_cell_wire[84];							inform_L[85][0] = l_cell_wire[85];							inform_L[86][0] = l_cell_wire[86];							inform_L[87][0] = l_cell_wire[87];							inform_L[88][0] = l_cell_wire[88];							inform_L[89][0] = l_cell_wire[89];							inform_L[90][0] = l_cell_wire[90];							inform_L[91][0] = l_cell_wire[91];							inform_L[92][0] = l_cell_wire[92];							inform_L[93][0] = l_cell_wire[93];							inform_L[94][0] = l_cell_wire[94];							inform_L[95][0] = l_cell_wire[95];							inform_L[96][0] = l_cell_wire[96];							inform_L[97][0] = l_cell_wire[97];							inform_L[98][0] = l_cell_wire[98];							inform_L[99][0] = l_cell_wire[99];							inform_L[100][0] = l_cell_wire[100];							inform_L[101][0] = l_cell_wire[101];							inform_L[102][0] = l_cell_wire[102];							inform_L[103][0] = l_cell_wire[103];							inform_L[104][0] = l_cell_wire[104];							inform_L[105][0] = l_cell_wire[105];							inform_L[106][0] = l_cell_wire[106];							inform_L[107][0] = l_cell_wire[107];							inform_L[108][0] = l_cell_wire[108];							inform_L[109][0] = l_cell_wire[109];							inform_L[110][0] = l_cell_wire[110];							inform_L[111][0] = l_cell_wire[111];							inform_L[112][0] = l_cell_wire[112];							inform_L[113][0] = l_cell_wire[113];							inform_L[114][0] = l_cell_wire[114];							inform_L[115][0] = l_cell_wire[115];							inform_L[116][0] = l_cell_wire[116];							inform_L[117][0] = l_cell_wire[117];							inform_L[118][0] = l_cell_wire[118];							inform_L[119][0] = l_cell_wire[119];							inform_L[120][0] = l_cell_wire[120];							inform_L[121][0] = l_cell_wire[121];							inform_L[122][0] = l_cell_wire[122];							inform_L[123][0] = l_cell_wire[123];							inform_L[124][0] = l_cell_wire[124];							inform_L[125][0] = l_cell_wire[125];							inform_L[126][0] = l_cell_wire[126];							inform_L[127][0] = l_cell_wire[127];							inform_L[128][0] = l_cell_wire[128];							inform_L[129][0] = l_cell_wire[129];							inform_L[130][0] = l_cell_wire[130];							inform_L[131][0] = l_cell_wire[131];							inform_L[132][0] = l_cell_wire[132];							inform_L[133][0] = l_cell_wire[133];							inform_L[134][0] = l_cell_wire[134];							inform_L[135][0] = l_cell_wire[135];							inform_L[136][0] = l_cell_wire[136];							inform_L[137][0] = l_cell_wire[137];							inform_L[138][0] = l_cell_wire[138];							inform_L[139][0] = l_cell_wire[139];							inform_L[140][0] = l_cell_wire[140];							inform_L[141][0] = l_cell_wire[141];							inform_L[142][0] = l_cell_wire[142];							inform_L[143][0] = l_cell_wire[143];							inform_L[144][0] = l_cell_wire[144];							inform_L[145][0] = l_cell_wire[145];							inform_L[146][0] = l_cell_wire[146];							inform_L[147][0] = l_cell_wire[147];							inform_L[148][0] = l_cell_wire[148];							inform_L[149][0] = l_cell_wire[149];							inform_L[150][0] = l_cell_wire[150];							inform_L[151][0] = l_cell_wire[151];							inform_L[152][0] = l_cell_wire[152];							inform_L[153][0] = l_cell_wire[153];							inform_L[154][0] = l_cell_wire[154];							inform_L[155][0] = l_cell_wire[155];							inform_L[156][0] = l_cell_wire[156];							inform_L[157][0] = l_cell_wire[157];							inform_L[158][0] = l_cell_wire[158];							inform_L[159][0] = l_cell_wire[159];							inform_L[160][0] = l_cell_wire[160];							inform_L[161][0] = l_cell_wire[161];							inform_L[162][0] = l_cell_wire[162];							inform_L[163][0] = l_cell_wire[163];							inform_L[164][0] = l_cell_wire[164];							inform_L[165][0] = l_cell_wire[165];							inform_L[166][0] = l_cell_wire[166];							inform_L[167][0] = l_cell_wire[167];							inform_L[168][0] = l_cell_wire[168];							inform_L[169][0] = l_cell_wire[169];							inform_L[170][0] = l_cell_wire[170];							inform_L[171][0] = l_cell_wire[171];							inform_L[172][0] = l_cell_wire[172];							inform_L[173][0] = l_cell_wire[173];							inform_L[174][0] = l_cell_wire[174];							inform_L[175][0] = l_cell_wire[175];							inform_L[176][0] = l_cell_wire[176];							inform_L[177][0] = l_cell_wire[177];							inform_L[178][0] = l_cell_wire[178];							inform_L[179][0] = l_cell_wire[179];							inform_L[180][0] = l_cell_wire[180];							inform_L[181][0] = l_cell_wire[181];							inform_L[182][0] = l_cell_wire[182];							inform_L[183][0] = l_cell_wire[183];							inform_L[184][0] = l_cell_wire[184];							inform_L[185][0] = l_cell_wire[185];							inform_L[186][0] = l_cell_wire[186];							inform_L[187][0] = l_cell_wire[187];							inform_L[188][0] = l_cell_wire[188];							inform_L[189][0] = l_cell_wire[189];							inform_L[190][0] = l_cell_wire[190];							inform_L[191][0] = l_cell_wire[191];							inform_L[192][0] = l_cell_wire[192];							inform_L[193][0] = l_cell_wire[193];							inform_L[194][0] = l_cell_wire[194];							inform_L[195][0] = l_cell_wire[195];							inform_L[196][0] = l_cell_wire[196];							inform_L[197][0] = l_cell_wire[197];							inform_L[198][0] = l_cell_wire[198];							inform_L[199][0] = l_cell_wire[199];							inform_L[200][0] = l_cell_wire[200];							inform_L[201][0] = l_cell_wire[201];							inform_L[202][0] = l_cell_wire[202];							inform_L[203][0] = l_cell_wire[203];							inform_L[204][0] = l_cell_wire[204];							inform_L[205][0] = l_cell_wire[205];							inform_L[206][0] = l_cell_wire[206];							inform_L[207][0] = l_cell_wire[207];							inform_L[208][0] = l_cell_wire[208];							inform_L[209][0] = l_cell_wire[209];							inform_L[210][0] = l_cell_wire[210];							inform_L[211][0] = l_cell_wire[211];							inform_L[212][0] = l_cell_wire[212];							inform_L[213][0] = l_cell_wire[213];							inform_L[214][0] = l_cell_wire[214];							inform_L[215][0] = l_cell_wire[215];							inform_L[216][0] = l_cell_wire[216];							inform_L[217][0] = l_cell_wire[217];							inform_L[218][0] = l_cell_wire[218];							inform_L[219][0] = l_cell_wire[219];							inform_L[220][0] = l_cell_wire[220];							inform_L[221][0] = l_cell_wire[221];							inform_L[222][0] = l_cell_wire[222];							inform_L[223][0] = l_cell_wire[223];							inform_L[224][0] = l_cell_wire[224];							inform_L[225][0] = l_cell_wire[225];							inform_L[226][0] = l_cell_wire[226];							inform_L[227][0] = l_cell_wire[227];							inform_L[228][0] = l_cell_wire[228];							inform_L[229][0] = l_cell_wire[229];							inform_L[230][0] = l_cell_wire[230];							inform_L[231][0] = l_cell_wire[231];							inform_L[232][0] = l_cell_wire[232];							inform_L[233][0] = l_cell_wire[233];							inform_L[234][0] = l_cell_wire[234];							inform_L[235][0] = l_cell_wire[235];							inform_L[236][0] = l_cell_wire[236];							inform_L[237][0] = l_cell_wire[237];							inform_L[238][0] = l_cell_wire[238];							inform_L[239][0] = l_cell_wire[239];							inform_L[240][0] = l_cell_wire[240];							inform_L[241][0] = l_cell_wire[241];							inform_L[242][0] = l_cell_wire[242];							inform_L[243][0] = l_cell_wire[243];							inform_L[244][0] = l_cell_wire[244];							inform_L[245][0] = l_cell_wire[245];							inform_L[246][0] = l_cell_wire[246];							inform_L[247][0] = l_cell_wire[247];							inform_L[248][0] = l_cell_wire[248];							inform_L[249][0] = l_cell_wire[249];							inform_L[250][0] = l_cell_wire[250];							inform_L[251][0] = l_cell_wire[251];							inform_L[252][0] = l_cell_wire[252];							inform_L[253][0] = l_cell_wire[253];							inform_L[254][0] = l_cell_wire[254];							inform_L[255][0] = l_cell_wire[255];						end
						2:						begin							inform_R[0][2] = r_cell_wire[0];							inform_R[2][2] = r_cell_wire[1];							inform_R[1][2] = r_cell_wire[2];							inform_R[3][2] = r_cell_wire[3];							inform_R[4][2] = r_cell_wire[4];							inform_R[6][2] = r_cell_wire[5];							inform_R[5][2] = r_cell_wire[6];							inform_R[7][2] = r_cell_wire[7];							inform_R[8][2] = r_cell_wire[8];							inform_R[10][2] = r_cell_wire[9];							inform_R[9][2] = r_cell_wire[10];							inform_R[11][2] = r_cell_wire[11];							inform_R[12][2] = r_cell_wire[12];							inform_R[14][2] = r_cell_wire[13];							inform_R[13][2] = r_cell_wire[14];							inform_R[15][2] = r_cell_wire[15];							inform_R[16][2] = r_cell_wire[16];							inform_R[18][2] = r_cell_wire[17];							inform_R[17][2] = r_cell_wire[18];							inform_R[19][2] = r_cell_wire[19];							inform_R[20][2] = r_cell_wire[20];							inform_R[22][2] = r_cell_wire[21];							inform_R[21][2] = r_cell_wire[22];							inform_R[23][2] = r_cell_wire[23];							inform_R[24][2] = r_cell_wire[24];							inform_R[26][2] = r_cell_wire[25];							inform_R[25][2] = r_cell_wire[26];							inform_R[27][2] = r_cell_wire[27];							inform_R[28][2] = r_cell_wire[28];							inform_R[30][2] = r_cell_wire[29];							inform_R[29][2] = r_cell_wire[30];							inform_R[31][2] = r_cell_wire[31];							inform_R[32][2] = r_cell_wire[32];							inform_R[34][2] = r_cell_wire[33];							inform_R[33][2] = r_cell_wire[34];							inform_R[35][2] = r_cell_wire[35];							inform_R[36][2] = r_cell_wire[36];							inform_R[38][2] = r_cell_wire[37];							inform_R[37][2] = r_cell_wire[38];							inform_R[39][2] = r_cell_wire[39];							inform_R[40][2] = r_cell_wire[40];							inform_R[42][2] = r_cell_wire[41];							inform_R[41][2] = r_cell_wire[42];							inform_R[43][2] = r_cell_wire[43];							inform_R[44][2] = r_cell_wire[44];							inform_R[46][2] = r_cell_wire[45];							inform_R[45][2] = r_cell_wire[46];							inform_R[47][2] = r_cell_wire[47];							inform_R[48][2] = r_cell_wire[48];							inform_R[50][2] = r_cell_wire[49];							inform_R[49][2] = r_cell_wire[50];							inform_R[51][2] = r_cell_wire[51];							inform_R[52][2] = r_cell_wire[52];							inform_R[54][2] = r_cell_wire[53];							inform_R[53][2] = r_cell_wire[54];							inform_R[55][2] = r_cell_wire[55];							inform_R[56][2] = r_cell_wire[56];							inform_R[58][2] = r_cell_wire[57];							inform_R[57][2] = r_cell_wire[58];							inform_R[59][2] = r_cell_wire[59];							inform_R[60][2] = r_cell_wire[60];							inform_R[62][2] = r_cell_wire[61];							inform_R[61][2] = r_cell_wire[62];							inform_R[63][2] = r_cell_wire[63];							inform_R[64][2] = r_cell_wire[64];							inform_R[66][2] = r_cell_wire[65];							inform_R[65][2] = r_cell_wire[66];							inform_R[67][2] = r_cell_wire[67];							inform_R[68][2] = r_cell_wire[68];							inform_R[70][2] = r_cell_wire[69];							inform_R[69][2] = r_cell_wire[70];							inform_R[71][2] = r_cell_wire[71];							inform_R[72][2] = r_cell_wire[72];							inform_R[74][2] = r_cell_wire[73];							inform_R[73][2] = r_cell_wire[74];							inform_R[75][2] = r_cell_wire[75];							inform_R[76][2] = r_cell_wire[76];							inform_R[78][2] = r_cell_wire[77];							inform_R[77][2] = r_cell_wire[78];							inform_R[79][2] = r_cell_wire[79];							inform_R[80][2] = r_cell_wire[80];							inform_R[82][2] = r_cell_wire[81];							inform_R[81][2] = r_cell_wire[82];							inform_R[83][2] = r_cell_wire[83];							inform_R[84][2] = r_cell_wire[84];							inform_R[86][2] = r_cell_wire[85];							inform_R[85][2] = r_cell_wire[86];							inform_R[87][2] = r_cell_wire[87];							inform_R[88][2] = r_cell_wire[88];							inform_R[90][2] = r_cell_wire[89];							inform_R[89][2] = r_cell_wire[90];							inform_R[91][2] = r_cell_wire[91];							inform_R[92][2] = r_cell_wire[92];							inform_R[94][2] = r_cell_wire[93];							inform_R[93][2] = r_cell_wire[94];							inform_R[95][2] = r_cell_wire[95];							inform_R[96][2] = r_cell_wire[96];							inform_R[98][2] = r_cell_wire[97];							inform_R[97][2] = r_cell_wire[98];							inform_R[99][2] = r_cell_wire[99];							inform_R[100][2] = r_cell_wire[100];							inform_R[102][2] = r_cell_wire[101];							inform_R[101][2] = r_cell_wire[102];							inform_R[103][2] = r_cell_wire[103];							inform_R[104][2] = r_cell_wire[104];							inform_R[106][2] = r_cell_wire[105];							inform_R[105][2] = r_cell_wire[106];							inform_R[107][2] = r_cell_wire[107];							inform_R[108][2] = r_cell_wire[108];							inform_R[110][2] = r_cell_wire[109];							inform_R[109][2] = r_cell_wire[110];							inform_R[111][2] = r_cell_wire[111];							inform_R[112][2] = r_cell_wire[112];							inform_R[114][2] = r_cell_wire[113];							inform_R[113][2] = r_cell_wire[114];							inform_R[115][2] = r_cell_wire[115];							inform_R[116][2] = r_cell_wire[116];							inform_R[118][2] = r_cell_wire[117];							inform_R[117][2] = r_cell_wire[118];							inform_R[119][2] = r_cell_wire[119];							inform_R[120][2] = r_cell_wire[120];							inform_R[122][2] = r_cell_wire[121];							inform_R[121][2] = r_cell_wire[122];							inform_R[123][2] = r_cell_wire[123];							inform_R[124][2] = r_cell_wire[124];							inform_R[126][2] = r_cell_wire[125];							inform_R[125][2] = r_cell_wire[126];							inform_R[127][2] = r_cell_wire[127];							inform_R[128][2] = r_cell_wire[128];							inform_R[130][2] = r_cell_wire[129];							inform_R[129][2] = r_cell_wire[130];							inform_R[131][2] = r_cell_wire[131];							inform_R[132][2] = r_cell_wire[132];							inform_R[134][2] = r_cell_wire[133];							inform_R[133][2] = r_cell_wire[134];							inform_R[135][2] = r_cell_wire[135];							inform_R[136][2] = r_cell_wire[136];							inform_R[138][2] = r_cell_wire[137];							inform_R[137][2] = r_cell_wire[138];							inform_R[139][2] = r_cell_wire[139];							inform_R[140][2] = r_cell_wire[140];							inform_R[142][2] = r_cell_wire[141];							inform_R[141][2] = r_cell_wire[142];							inform_R[143][2] = r_cell_wire[143];							inform_R[144][2] = r_cell_wire[144];							inform_R[146][2] = r_cell_wire[145];							inform_R[145][2] = r_cell_wire[146];							inform_R[147][2] = r_cell_wire[147];							inform_R[148][2] = r_cell_wire[148];							inform_R[150][2] = r_cell_wire[149];							inform_R[149][2] = r_cell_wire[150];							inform_R[151][2] = r_cell_wire[151];							inform_R[152][2] = r_cell_wire[152];							inform_R[154][2] = r_cell_wire[153];							inform_R[153][2] = r_cell_wire[154];							inform_R[155][2] = r_cell_wire[155];							inform_R[156][2] = r_cell_wire[156];							inform_R[158][2] = r_cell_wire[157];							inform_R[157][2] = r_cell_wire[158];							inform_R[159][2] = r_cell_wire[159];							inform_R[160][2] = r_cell_wire[160];							inform_R[162][2] = r_cell_wire[161];							inform_R[161][2] = r_cell_wire[162];							inform_R[163][2] = r_cell_wire[163];							inform_R[164][2] = r_cell_wire[164];							inform_R[166][2] = r_cell_wire[165];							inform_R[165][2] = r_cell_wire[166];							inform_R[167][2] = r_cell_wire[167];							inform_R[168][2] = r_cell_wire[168];							inform_R[170][2] = r_cell_wire[169];							inform_R[169][2] = r_cell_wire[170];							inform_R[171][2] = r_cell_wire[171];							inform_R[172][2] = r_cell_wire[172];							inform_R[174][2] = r_cell_wire[173];							inform_R[173][2] = r_cell_wire[174];							inform_R[175][2] = r_cell_wire[175];							inform_R[176][2] = r_cell_wire[176];							inform_R[178][2] = r_cell_wire[177];							inform_R[177][2] = r_cell_wire[178];							inform_R[179][2] = r_cell_wire[179];							inform_R[180][2] = r_cell_wire[180];							inform_R[182][2] = r_cell_wire[181];							inform_R[181][2] = r_cell_wire[182];							inform_R[183][2] = r_cell_wire[183];							inform_R[184][2] = r_cell_wire[184];							inform_R[186][2] = r_cell_wire[185];							inform_R[185][2] = r_cell_wire[186];							inform_R[187][2] = r_cell_wire[187];							inform_R[188][2] = r_cell_wire[188];							inform_R[190][2] = r_cell_wire[189];							inform_R[189][2] = r_cell_wire[190];							inform_R[191][2] = r_cell_wire[191];							inform_R[192][2] = r_cell_wire[192];							inform_R[194][2] = r_cell_wire[193];							inform_R[193][2] = r_cell_wire[194];							inform_R[195][2] = r_cell_wire[195];							inform_R[196][2] = r_cell_wire[196];							inform_R[198][2] = r_cell_wire[197];							inform_R[197][2] = r_cell_wire[198];							inform_R[199][2] = r_cell_wire[199];							inform_R[200][2] = r_cell_wire[200];							inform_R[202][2] = r_cell_wire[201];							inform_R[201][2] = r_cell_wire[202];							inform_R[203][2] = r_cell_wire[203];							inform_R[204][2] = r_cell_wire[204];							inform_R[206][2] = r_cell_wire[205];							inform_R[205][2] = r_cell_wire[206];							inform_R[207][2] = r_cell_wire[207];							inform_R[208][2] = r_cell_wire[208];							inform_R[210][2] = r_cell_wire[209];							inform_R[209][2] = r_cell_wire[210];							inform_R[211][2] = r_cell_wire[211];							inform_R[212][2] = r_cell_wire[212];							inform_R[214][2] = r_cell_wire[213];							inform_R[213][2] = r_cell_wire[214];							inform_R[215][2] = r_cell_wire[215];							inform_R[216][2] = r_cell_wire[216];							inform_R[218][2] = r_cell_wire[217];							inform_R[217][2] = r_cell_wire[218];							inform_R[219][2] = r_cell_wire[219];							inform_R[220][2] = r_cell_wire[220];							inform_R[222][2] = r_cell_wire[221];							inform_R[221][2] = r_cell_wire[222];							inform_R[223][2] = r_cell_wire[223];							inform_R[224][2] = r_cell_wire[224];							inform_R[226][2] = r_cell_wire[225];							inform_R[225][2] = r_cell_wire[226];							inform_R[227][2] = r_cell_wire[227];							inform_R[228][2] = r_cell_wire[228];							inform_R[230][2] = r_cell_wire[229];							inform_R[229][2] = r_cell_wire[230];							inform_R[231][2] = r_cell_wire[231];							inform_R[232][2] = r_cell_wire[232];							inform_R[234][2] = r_cell_wire[233];							inform_R[233][2] = r_cell_wire[234];							inform_R[235][2] = r_cell_wire[235];							inform_R[236][2] = r_cell_wire[236];							inform_R[238][2] = r_cell_wire[237];							inform_R[237][2] = r_cell_wire[238];							inform_R[239][2] = r_cell_wire[239];							inform_R[240][2] = r_cell_wire[240];							inform_R[242][2] = r_cell_wire[241];							inform_R[241][2] = r_cell_wire[242];							inform_R[243][2] = r_cell_wire[243];							inform_R[244][2] = r_cell_wire[244];							inform_R[246][2] = r_cell_wire[245];							inform_R[245][2] = r_cell_wire[246];							inform_R[247][2] = r_cell_wire[247];							inform_R[248][2] = r_cell_wire[248];							inform_R[250][2] = r_cell_wire[249];							inform_R[249][2] = r_cell_wire[250];							inform_R[251][2] = r_cell_wire[251];							inform_R[252][2] = r_cell_wire[252];							inform_R[254][2] = r_cell_wire[253];							inform_R[253][2] = r_cell_wire[254];							inform_R[255][2] = r_cell_wire[255];							inform_L[0][1] = l_cell_wire[0];							inform_L[2][1] = l_cell_wire[1];							inform_L[1][1] = l_cell_wire[2];							inform_L[3][1] = l_cell_wire[3];							inform_L[4][1] = l_cell_wire[4];							inform_L[6][1] = l_cell_wire[5];							inform_L[5][1] = l_cell_wire[6];							inform_L[7][1] = l_cell_wire[7];							inform_L[8][1] = l_cell_wire[8];							inform_L[10][1] = l_cell_wire[9];							inform_L[9][1] = l_cell_wire[10];							inform_L[11][1] = l_cell_wire[11];							inform_L[12][1] = l_cell_wire[12];							inform_L[14][1] = l_cell_wire[13];							inform_L[13][1] = l_cell_wire[14];							inform_L[15][1] = l_cell_wire[15];							inform_L[16][1] = l_cell_wire[16];							inform_L[18][1] = l_cell_wire[17];							inform_L[17][1] = l_cell_wire[18];							inform_L[19][1] = l_cell_wire[19];							inform_L[20][1] = l_cell_wire[20];							inform_L[22][1] = l_cell_wire[21];							inform_L[21][1] = l_cell_wire[22];							inform_L[23][1] = l_cell_wire[23];							inform_L[24][1] = l_cell_wire[24];							inform_L[26][1] = l_cell_wire[25];							inform_L[25][1] = l_cell_wire[26];							inform_L[27][1] = l_cell_wire[27];							inform_L[28][1] = l_cell_wire[28];							inform_L[30][1] = l_cell_wire[29];							inform_L[29][1] = l_cell_wire[30];							inform_L[31][1] = l_cell_wire[31];							inform_L[32][1] = l_cell_wire[32];							inform_L[34][1] = l_cell_wire[33];							inform_L[33][1] = l_cell_wire[34];							inform_L[35][1] = l_cell_wire[35];							inform_L[36][1] = l_cell_wire[36];							inform_L[38][1] = l_cell_wire[37];							inform_L[37][1] = l_cell_wire[38];							inform_L[39][1] = l_cell_wire[39];							inform_L[40][1] = l_cell_wire[40];							inform_L[42][1] = l_cell_wire[41];							inform_L[41][1] = l_cell_wire[42];							inform_L[43][1] = l_cell_wire[43];							inform_L[44][1] = l_cell_wire[44];							inform_L[46][1] = l_cell_wire[45];							inform_L[45][1] = l_cell_wire[46];							inform_L[47][1] = l_cell_wire[47];							inform_L[48][1] = l_cell_wire[48];							inform_L[50][1] = l_cell_wire[49];							inform_L[49][1] = l_cell_wire[50];							inform_L[51][1] = l_cell_wire[51];							inform_L[52][1] = l_cell_wire[52];							inform_L[54][1] = l_cell_wire[53];							inform_L[53][1] = l_cell_wire[54];							inform_L[55][1] = l_cell_wire[55];							inform_L[56][1] = l_cell_wire[56];							inform_L[58][1] = l_cell_wire[57];							inform_L[57][1] = l_cell_wire[58];							inform_L[59][1] = l_cell_wire[59];							inform_L[60][1] = l_cell_wire[60];							inform_L[62][1] = l_cell_wire[61];							inform_L[61][1] = l_cell_wire[62];							inform_L[63][1] = l_cell_wire[63];							inform_L[64][1] = l_cell_wire[64];							inform_L[66][1] = l_cell_wire[65];							inform_L[65][1] = l_cell_wire[66];							inform_L[67][1] = l_cell_wire[67];							inform_L[68][1] = l_cell_wire[68];							inform_L[70][1] = l_cell_wire[69];							inform_L[69][1] = l_cell_wire[70];							inform_L[71][1] = l_cell_wire[71];							inform_L[72][1] = l_cell_wire[72];							inform_L[74][1] = l_cell_wire[73];							inform_L[73][1] = l_cell_wire[74];							inform_L[75][1] = l_cell_wire[75];							inform_L[76][1] = l_cell_wire[76];							inform_L[78][1] = l_cell_wire[77];							inform_L[77][1] = l_cell_wire[78];							inform_L[79][1] = l_cell_wire[79];							inform_L[80][1] = l_cell_wire[80];							inform_L[82][1] = l_cell_wire[81];							inform_L[81][1] = l_cell_wire[82];							inform_L[83][1] = l_cell_wire[83];							inform_L[84][1] = l_cell_wire[84];							inform_L[86][1] = l_cell_wire[85];							inform_L[85][1] = l_cell_wire[86];							inform_L[87][1] = l_cell_wire[87];							inform_L[88][1] = l_cell_wire[88];							inform_L[90][1] = l_cell_wire[89];							inform_L[89][1] = l_cell_wire[90];							inform_L[91][1] = l_cell_wire[91];							inform_L[92][1] = l_cell_wire[92];							inform_L[94][1] = l_cell_wire[93];							inform_L[93][1] = l_cell_wire[94];							inform_L[95][1] = l_cell_wire[95];							inform_L[96][1] = l_cell_wire[96];							inform_L[98][1] = l_cell_wire[97];							inform_L[97][1] = l_cell_wire[98];							inform_L[99][1] = l_cell_wire[99];							inform_L[100][1] = l_cell_wire[100];							inform_L[102][1] = l_cell_wire[101];							inform_L[101][1] = l_cell_wire[102];							inform_L[103][1] = l_cell_wire[103];							inform_L[104][1] = l_cell_wire[104];							inform_L[106][1] = l_cell_wire[105];							inform_L[105][1] = l_cell_wire[106];							inform_L[107][1] = l_cell_wire[107];							inform_L[108][1] = l_cell_wire[108];							inform_L[110][1] = l_cell_wire[109];							inform_L[109][1] = l_cell_wire[110];							inform_L[111][1] = l_cell_wire[111];							inform_L[112][1] = l_cell_wire[112];							inform_L[114][1] = l_cell_wire[113];							inform_L[113][1] = l_cell_wire[114];							inform_L[115][1] = l_cell_wire[115];							inform_L[116][1] = l_cell_wire[116];							inform_L[118][1] = l_cell_wire[117];							inform_L[117][1] = l_cell_wire[118];							inform_L[119][1] = l_cell_wire[119];							inform_L[120][1] = l_cell_wire[120];							inform_L[122][1] = l_cell_wire[121];							inform_L[121][1] = l_cell_wire[122];							inform_L[123][1] = l_cell_wire[123];							inform_L[124][1] = l_cell_wire[124];							inform_L[126][1] = l_cell_wire[125];							inform_L[125][1] = l_cell_wire[126];							inform_L[127][1] = l_cell_wire[127];							inform_L[128][1] = l_cell_wire[128];							inform_L[130][1] = l_cell_wire[129];							inform_L[129][1] = l_cell_wire[130];							inform_L[131][1] = l_cell_wire[131];							inform_L[132][1] = l_cell_wire[132];							inform_L[134][1] = l_cell_wire[133];							inform_L[133][1] = l_cell_wire[134];							inform_L[135][1] = l_cell_wire[135];							inform_L[136][1] = l_cell_wire[136];							inform_L[138][1] = l_cell_wire[137];							inform_L[137][1] = l_cell_wire[138];							inform_L[139][1] = l_cell_wire[139];							inform_L[140][1] = l_cell_wire[140];							inform_L[142][1] = l_cell_wire[141];							inform_L[141][1] = l_cell_wire[142];							inform_L[143][1] = l_cell_wire[143];							inform_L[144][1] = l_cell_wire[144];							inform_L[146][1] = l_cell_wire[145];							inform_L[145][1] = l_cell_wire[146];							inform_L[147][1] = l_cell_wire[147];							inform_L[148][1] = l_cell_wire[148];							inform_L[150][1] = l_cell_wire[149];							inform_L[149][1] = l_cell_wire[150];							inform_L[151][1] = l_cell_wire[151];							inform_L[152][1] = l_cell_wire[152];							inform_L[154][1] = l_cell_wire[153];							inform_L[153][1] = l_cell_wire[154];							inform_L[155][1] = l_cell_wire[155];							inform_L[156][1] = l_cell_wire[156];							inform_L[158][1] = l_cell_wire[157];							inform_L[157][1] = l_cell_wire[158];							inform_L[159][1] = l_cell_wire[159];							inform_L[160][1] = l_cell_wire[160];							inform_L[162][1] = l_cell_wire[161];							inform_L[161][1] = l_cell_wire[162];							inform_L[163][1] = l_cell_wire[163];							inform_L[164][1] = l_cell_wire[164];							inform_L[166][1] = l_cell_wire[165];							inform_L[165][1] = l_cell_wire[166];							inform_L[167][1] = l_cell_wire[167];							inform_L[168][1] = l_cell_wire[168];							inform_L[170][1] = l_cell_wire[169];							inform_L[169][1] = l_cell_wire[170];							inform_L[171][1] = l_cell_wire[171];							inform_L[172][1] = l_cell_wire[172];							inform_L[174][1] = l_cell_wire[173];							inform_L[173][1] = l_cell_wire[174];							inform_L[175][1] = l_cell_wire[175];							inform_L[176][1] = l_cell_wire[176];							inform_L[178][1] = l_cell_wire[177];							inform_L[177][1] = l_cell_wire[178];							inform_L[179][1] = l_cell_wire[179];							inform_L[180][1] = l_cell_wire[180];							inform_L[182][1] = l_cell_wire[181];							inform_L[181][1] = l_cell_wire[182];							inform_L[183][1] = l_cell_wire[183];							inform_L[184][1] = l_cell_wire[184];							inform_L[186][1] = l_cell_wire[185];							inform_L[185][1] = l_cell_wire[186];							inform_L[187][1] = l_cell_wire[187];							inform_L[188][1] = l_cell_wire[188];							inform_L[190][1] = l_cell_wire[189];							inform_L[189][1] = l_cell_wire[190];							inform_L[191][1] = l_cell_wire[191];							inform_L[192][1] = l_cell_wire[192];							inform_L[194][1] = l_cell_wire[193];							inform_L[193][1] = l_cell_wire[194];							inform_L[195][1] = l_cell_wire[195];							inform_L[196][1] = l_cell_wire[196];							inform_L[198][1] = l_cell_wire[197];							inform_L[197][1] = l_cell_wire[198];							inform_L[199][1] = l_cell_wire[199];							inform_L[200][1] = l_cell_wire[200];							inform_L[202][1] = l_cell_wire[201];							inform_L[201][1] = l_cell_wire[202];							inform_L[203][1] = l_cell_wire[203];							inform_L[204][1] = l_cell_wire[204];							inform_L[206][1] = l_cell_wire[205];							inform_L[205][1] = l_cell_wire[206];							inform_L[207][1] = l_cell_wire[207];							inform_L[208][1] = l_cell_wire[208];							inform_L[210][1] = l_cell_wire[209];							inform_L[209][1] = l_cell_wire[210];							inform_L[211][1] = l_cell_wire[211];							inform_L[212][1] = l_cell_wire[212];							inform_L[214][1] = l_cell_wire[213];							inform_L[213][1] = l_cell_wire[214];							inform_L[215][1] = l_cell_wire[215];							inform_L[216][1] = l_cell_wire[216];							inform_L[218][1] = l_cell_wire[217];							inform_L[217][1] = l_cell_wire[218];							inform_L[219][1] = l_cell_wire[219];							inform_L[220][1] = l_cell_wire[220];							inform_L[222][1] = l_cell_wire[221];							inform_L[221][1] = l_cell_wire[222];							inform_L[223][1] = l_cell_wire[223];							inform_L[224][1] = l_cell_wire[224];							inform_L[226][1] = l_cell_wire[225];							inform_L[225][1] = l_cell_wire[226];							inform_L[227][1] = l_cell_wire[227];							inform_L[228][1] = l_cell_wire[228];							inform_L[230][1] = l_cell_wire[229];							inform_L[229][1] = l_cell_wire[230];							inform_L[231][1] = l_cell_wire[231];							inform_L[232][1] = l_cell_wire[232];							inform_L[234][1] = l_cell_wire[233];							inform_L[233][1] = l_cell_wire[234];							inform_L[235][1] = l_cell_wire[235];							inform_L[236][1] = l_cell_wire[236];							inform_L[238][1] = l_cell_wire[237];							inform_L[237][1] = l_cell_wire[238];							inform_L[239][1] = l_cell_wire[239];							inform_L[240][1] = l_cell_wire[240];							inform_L[242][1] = l_cell_wire[241];							inform_L[241][1] = l_cell_wire[242];							inform_L[243][1] = l_cell_wire[243];							inform_L[244][1] = l_cell_wire[244];							inform_L[246][1] = l_cell_wire[245];							inform_L[245][1] = l_cell_wire[246];							inform_L[247][1] = l_cell_wire[247];							inform_L[248][1] = l_cell_wire[248];							inform_L[250][1] = l_cell_wire[249];							inform_L[249][1] = l_cell_wire[250];							inform_L[251][1] = l_cell_wire[251];							inform_L[252][1] = l_cell_wire[252];							inform_L[254][1] = l_cell_wire[253];							inform_L[253][1] = l_cell_wire[254];							inform_L[255][1] = l_cell_wire[255];						end
						3:						begin							inform_R[0][3] = r_cell_wire[0];							inform_R[4][3] = r_cell_wire[1];							inform_R[1][3] = r_cell_wire[2];							inform_R[5][3] = r_cell_wire[3];							inform_R[2][3] = r_cell_wire[4];							inform_R[6][3] = r_cell_wire[5];							inform_R[3][3] = r_cell_wire[6];							inform_R[7][3] = r_cell_wire[7];							inform_R[8][3] = r_cell_wire[8];							inform_R[12][3] = r_cell_wire[9];							inform_R[9][3] = r_cell_wire[10];							inform_R[13][3] = r_cell_wire[11];							inform_R[10][3] = r_cell_wire[12];							inform_R[14][3] = r_cell_wire[13];							inform_R[11][3] = r_cell_wire[14];							inform_R[15][3] = r_cell_wire[15];							inform_R[16][3] = r_cell_wire[16];							inform_R[20][3] = r_cell_wire[17];							inform_R[17][3] = r_cell_wire[18];							inform_R[21][3] = r_cell_wire[19];							inform_R[18][3] = r_cell_wire[20];							inform_R[22][3] = r_cell_wire[21];							inform_R[19][3] = r_cell_wire[22];							inform_R[23][3] = r_cell_wire[23];							inform_R[24][3] = r_cell_wire[24];							inform_R[28][3] = r_cell_wire[25];							inform_R[25][3] = r_cell_wire[26];							inform_R[29][3] = r_cell_wire[27];							inform_R[26][3] = r_cell_wire[28];							inform_R[30][3] = r_cell_wire[29];							inform_R[27][3] = r_cell_wire[30];							inform_R[31][3] = r_cell_wire[31];							inform_R[32][3] = r_cell_wire[32];							inform_R[36][3] = r_cell_wire[33];							inform_R[33][3] = r_cell_wire[34];							inform_R[37][3] = r_cell_wire[35];							inform_R[34][3] = r_cell_wire[36];							inform_R[38][3] = r_cell_wire[37];							inform_R[35][3] = r_cell_wire[38];							inform_R[39][3] = r_cell_wire[39];							inform_R[40][3] = r_cell_wire[40];							inform_R[44][3] = r_cell_wire[41];							inform_R[41][3] = r_cell_wire[42];							inform_R[45][3] = r_cell_wire[43];							inform_R[42][3] = r_cell_wire[44];							inform_R[46][3] = r_cell_wire[45];							inform_R[43][3] = r_cell_wire[46];							inform_R[47][3] = r_cell_wire[47];							inform_R[48][3] = r_cell_wire[48];							inform_R[52][3] = r_cell_wire[49];							inform_R[49][3] = r_cell_wire[50];							inform_R[53][3] = r_cell_wire[51];							inform_R[50][3] = r_cell_wire[52];							inform_R[54][3] = r_cell_wire[53];							inform_R[51][3] = r_cell_wire[54];							inform_R[55][3] = r_cell_wire[55];							inform_R[56][3] = r_cell_wire[56];							inform_R[60][3] = r_cell_wire[57];							inform_R[57][3] = r_cell_wire[58];							inform_R[61][3] = r_cell_wire[59];							inform_R[58][3] = r_cell_wire[60];							inform_R[62][3] = r_cell_wire[61];							inform_R[59][3] = r_cell_wire[62];							inform_R[63][3] = r_cell_wire[63];							inform_R[64][3] = r_cell_wire[64];							inform_R[68][3] = r_cell_wire[65];							inform_R[65][3] = r_cell_wire[66];							inform_R[69][3] = r_cell_wire[67];							inform_R[66][3] = r_cell_wire[68];							inform_R[70][3] = r_cell_wire[69];							inform_R[67][3] = r_cell_wire[70];							inform_R[71][3] = r_cell_wire[71];							inform_R[72][3] = r_cell_wire[72];							inform_R[76][3] = r_cell_wire[73];							inform_R[73][3] = r_cell_wire[74];							inform_R[77][3] = r_cell_wire[75];							inform_R[74][3] = r_cell_wire[76];							inform_R[78][3] = r_cell_wire[77];							inform_R[75][3] = r_cell_wire[78];							inform_R[79][3] = r_cell_wire[79];							inform_R[80][3] = r_cell_wire[80];							inform_R[84][3] = r_cell_wire[81];							inform_R[81][3] = r_cell_wire[82];							inform_R[85][3] = r_cell_wire[83];							inform_R[82][3] = r_cell_wire[84];							inform_R[86][3] = r_cell_wire[85];							inform_R[83][3] = r_cell_wire[86];							inform_R[87][3] = r_cell_wire[87];							inform_R[88][3] = r_cell_wire[88];							inform_R[92][3] = r_cell_wire[89];							inform_R[89][3] = r_cell_wire[90];							inform_R[93][3] = r_cell_wire[91];							inform_R[90][3] = r_cell_wire[92];							inform_R[94][3] = r_cell_wire[93];							inform_R[91][3] = r_cell_wire[94];							inform_R[95][3] = r_cell_wire[95];							inform_R[96][3] = r_cell_wire[96];							inform_R[100][3] = r_cell_wire[97];							inform_R[97][3] = r_cell_wire[98];							inform_R[101][3] = r_cell_wire[99];							inform_R[98][3] = r_cell_wire[100];							inform_R[102][3] = r_cell_wire[101];							inform_R[99][3] = r_cell_wire[102];							inform_R[103][3] = r_cell_wire[103];							inform_R[104][3] = r_cell_wire[104];							inform_R[108][3] = r_cell_wire[105];							inform_R[105][3] = r_cell_wire[106];							inform_R[109][3] = r_cell_wire[107];							inform_R[106][3] = r_cell_wire[108];							inform_R[110][3] = r_cell_wire[109];							inform_R[107][3] = r_cell_wire[110];							inform_R[111][3] = r_cell_wire[111];							inform_R[112][3] = r_cell_wire[112];							inform_R[116][3] = r_cell_wire[113];							inform_R[113][3] = r_cell_wire[114];							inform_R[117][3] = r_cell_wire[115];							inform_R[114][3] = r_cell_wire[116];							inform_R[118][3] = r_cell_wire[117];							inform_R[115][3] = r_cell_wire[118];							inform_R[119][3] = r_cell_wire[119];							inform_R[120][3] = r_cell_wire[120];							inform_R[124][3] = r_cell_wire[121];							inform_R[121][3] = r_cell_wire[122];							inform_R[125][3] = r_cell_wire[123];							inform_R[122][3] = r_cell_wire[124];							inform_R[126][3] = r_cell_wire[125];							inform_R[123][3] = r_cell_wire[126];							inform_R[127][3] = r_cell_wire[127];							inform_R[128][3] = r_cell_wire[128];							inform_R[132][3] = r_cell_wire[129];							inform_R[129][3] = r_cell_wire[130];							inform_R[133][3] = r_cell_wire[131];							inform_R[130][3] = r_cell_wire[132];							inform_R[134][3] = r_cell_wire[133];							inform_R[131][3] = r_cell_wire[134];							inform_R[135][3] = r_cell_wire[135];							inform_R[136][3] = r_cell_wire[136];							inform_R[140][3] = r_cell_wire[137];							inform_R[137][3] = r_cell_wire[138];							inform_R[141][3] = r_cell_wire[139];							inform_R[138][3] = r_cell_wire[140];							inform_R[142][3] = r_cell_wire[141];							inform_R[139][3] = r_cell_wire[142];							inform_R[143][3] = r_cell_wire[143];							inform_R[144][3] = r_cell_wire[144];							inform_R[148][3] = r_cell_wire[145];							inform_R[145][3] = r_cell_wire[146];							inform_R[149][3] = r_cell_wire[147];							inform_R[146][3] = r_cell_wire[148];							inform_R[150][3] = r_cell_wire[149];							inform_R[147][3] = r_cell_wire[150];							inform_R[151][3] = r_cell_wire[151];							inform_R[152][3] = r_cell_wire[152];							inform_R[156][3] = r_cell_wire[153];							inform_R[153][3] = r_cell_wire[154];							inform_R[157][3] = r_cell_wire[155];							inform_R[154][3] = r_cell_wire[156];							inform_R[158][3] = r_cell_wire[157];							inform_R[155][3] = r_cell_wire[158];							inform_R[159][3] = r_cell_wire[159];							inform_R[160][3] = r_cell_wire[160];							inform_R[164][3] = r_cell_wire[161];							inform_R[161][3] = r_cell_wire[162];							inform_R[165][3] = r_cell_wire[163];							inform_R[162][3] = r_cell_wire[164];							inform_R[166][3] = r_cell_wire[165];							inform_R[163][3] = r_cell_wire[166];							inform_R[167][3] = r_cell_wire[167];							inform_R[168][3] = r_cell_wire[168];							inform_R[172][3] = r_cell_wire[169];							inform_R[169][3] = r_cell_wire[170];							inform_R[173][3] = r_cell_wire[171];							inform_R[170][3] = r_cell_wire[172];							inform_R[174][3] = r_cell_wire[173];							inform_R[171][3] = r_cell_wire[174];							inform_R[175][3] = r_cell_wire[175];							inform_R[176][3] = r_cell_wire[176];							inform_R[180][3] = r_cell_wire[177];							inform_R[177][3] = r_cell_wire[178];							inform_R[181][3] = r_cell_wire[179];							inform_R[178][3] = r_cell_wire[180];							inform_R[182][3] = r_cell_wire[181];							inform_R[179][3] = r_cell_wire[182];							inform_R[183][3] = r_cell_wire[183];							inform_R[184][3] = r_cell_wire[184];							inform_R[188][3] = r_cell_wire[185];							inform_R[185][3] = r_cell_wire[186];							inform_R[189][3] = r_cell_wire[187];							inform_R[186][3] = r_cell_wire[188];							inform_R[190][3] = r_cell_wire[189];							inform_R[187][3] = r_cell_wire[190];							inform_R[191][3] = r_cell_wire[191];							inform_R[192][3] = r_cell_wire[192];							inform_R[196][3] = r_cell_wire[193];							inform_R[193][3] = r_cell_wire[194];							inform_R[197][3] = r_cell_wire[195];							inform_R[194][3] = r_cell_wire[196];							inform_R[198][3] = r_cell_wire[197];							inform_R[195][3] = r_cell_wire[198];							inform_R[199][3] = r_cell_wire[199];							inform_R[200][3] = r_cell_wire[200];							inform_R[204][3] = r_cell_wire[201];							inform_R[201][3] = r_cell_wire[202];							inform_R[205][3] = r_cell_wire[203];							inform_R[202][3] = r_cell_wire[204];							inform_R[206][3] = r_cell_wire[205];							inform_R[203][3] = r_cell_wire[206];							inform_R[207][3] = r_cell_wire[207];							inform_R[208][3] = r_cell_wire[208];							inform_R[212][3] = r_cell_wire[209];							inform_R[209][3] = r_cell_wire[210];							inform_R[213][3] = r_cell_wire[211];							inform_R[210][3] = r_cell_wire[212];							inform_R[214][3] = r_cell_wire[213];							inform_R[211][3] = r_cell_wire[214];							inform_R[215][3] = r_cell_wire[215];							inform_R[216][3] = r_cell_wire[216];							inform_R[220][3] = r_cell_wire[217];							inform_R[217][3] = r_cell_wire[218];							inform_R[221][3] = r_cell_wire[219];							inform_R[218][3] = r_cell_wire[220];							inform_R[222][3] = r_cell_wire[221];							inform_R[219][3] = r_cell_wire[222];							inform_R[223][3] = r_cell_wire[223];							inform_R[224][3] = r_cell_wire[224];							inform_R[228][3] = r_cell_wire[225];							inform_R[225][3] = r_cell_wire[226];							inform_R[229][3] = r_cell_wire[227];							inform_R[226][3] = r_cell_wire[228];							inform_R[230][3] = r_cell_wire[229];							inform_R[227][3] = r_cell_wire[230];							inform_R[231][3] = r_cell_wire[231];							inform_R[232][3] = r_cell_wire[232];							inform_R[236][3] = r_cell_wire[233];							inform_R[233][3] = r_cell_wire[234];							inform_R[237][3] = r_cell_wire[235];							inform_R[234][3] = r_cell_wire[236];							inform_R[238][3] = r_cell_wire[237];							inform_R[235][3] = r_cell_wire[238];							inform_R[239][3] = r_cell_wire[239];							inform_R[240][3] = r_cell_wire[240];							inform_R[244][3] = r_cell_wire[241];							inform_R[241][3] = r_cell_wire[242];							inform_R[245][3] = r_cell_wire[243];							inform_R[242][3] = r_cell_wire[244];							inform_R[246][3] = r_cell_wire[245];							inform_R[243][3] = r_cell_wire[246];							inform_R[247][3] = r_cell_wire[247];							inform_R[248][3] = r_cell_wire[248];							inform_R[252][3] = r_cell_wire[249];							inform_R[249][3] = r_cell_wire[250];							inform_R[253][3] = r_cell_wire[251];							inform_R[250][3] = r_cell_wire[252];							inform_R[254][3] = r_cell_wire[253];							inform_R[251][3] = r_cell_wire[254];							inform_R[255][3] = r_cell_wire[255];							inform_L[0][2] = l_cell_wire[0];							inform_L[4][2] = l_cell_wire[1];							inform_L[1][2] = l_cell_wire[2];							inform_L[5][2] = l_cell_wire[3];							inform_L[2][2] = l_cell_wire[4];							inform_L[6][2] = l_cell_wire[5];							inform_L[3][2] = l_cell_wire[6];							inform_L[7][2] = l_cell_wire[7];							inform_L[8][2] = l_cell_wire[8];							inform_L[12][2] = l_cell_wire[9];							inform_L[9][2] = l_cell_wire[10];							inform_L[13][2] = l_cell_wire[11];							inform_L[10][2] = l_cell_wire[12];							inform_L[14][2] = l_cell_wire[13];							inform_L[11][2] = l_cell_wire[14];							inform_L[15][2] = l_cell_wire[15];							inform_L[16][2] = l_cell_wire[16];							inform_L[20][2] = l_cell_wire[17];							inform_L[17][2] = l_cell_wire[18];							inform_L[21][2] = l_cell_wire[19];							inform_L[18][2] = l_cell_wire[20];							inform_L[22][2] = l_cell_wire[21];							inform_L[19][2] = l_cell_wire[22];							inform_L[23][2] = l_cell_wire[23];							inform_L[24][2] = l_cell_wire[24];							inform_L[28][2] = l_cell_wire[25];							inform_L[25][2] = l_cell_wire[26];							inform_L[29][2] = l_cell_wire[27];							inform_L[26][2] = l_cell_wire[28];							inform_L[30][2] = l_cell_wire[29];							inform_L[27][2] = l_cell_wire[30];							inform_L[31][2] = l_cell_wire[31];							inform_L[32][2] = l_cell_wire[32];							inform_L[36][2] = l_cell_wire[33];							inform_L[33][2] = l_cell_wire[34];							inform_L[37][2] = l_cell_wire[35];							inform_L[34][2] = l_cell_wire[36];							inform_L[38][2] = l_cell_wire[37];							inform_L[35][2] = l_cell_wire[38];							inform_L[39][2] = l_cell_wire[39];							inform_L[40][2] = l_cell_wire[40];							inform_L[44][2] = l_cell_wire[41];							inform_L[41][2] = l_cell_wire[42];							inform_L[45][2] = l_cell_wire[43];							inform_L[42][2] = l_cell_wire[44];							inform_L[46][2] = l_cell_wire[45];							inform_L[43][2] = l_cell_wire[46];							inform_L[47][2] = l_cell_wire[47];							inform_L[48][2] = l_cell_wire[48];							inform_L[52][2] = l_cell_wire[49];							inform_L[49][2] = l_cell_wire[50];							inform_L[53][2] = l_cell_wire[51];							inform_L[50][2] = l_cell_wire[52];							inform_L[54][2] = l_cell_wire[53];							inform_L[51][2] = l_cell_wire[54];							inform_L[55][2] = l_cell_wire[55];							inform_L[56][2] = l_cell_wire[56];							inform_L[60][2] = l_cell_wire[57];							inform_L[57][2] = l_cell_wire[58];							inform_L[61][2] = l_cell_wire[59];							inform_L[58][2] = l_cell_wire[60];							inform_L[62][2] = l_cell_wire[61];							inform_L[59][2] = l_cell_wire[62];							inform_L[63][2] = l_cell_wire[63];							inform_L[64][2] = l_cell_wire[64];							inform_L[68][2] = l_cell_wire[65];							inform_L[65][2] = l_cell_wire[66];							inform_L[69][2] = l_cell_wire[67];							inform_L[66][2] = l_cell_wire[68];							inform_L[70][2] = l_cell_wire[69];							inform_L[67][2] = l_cell_wire[70];							inform_L[71][2] = l_cell_wire[71];							inform_L[72][2] = l_cell_wire[72];							inform_L[76][2] = l_cell_wire[73];							inform_L[73][2] = l_cell_wire[74];							inform_L[77][2] = l_cell_wire[75];							inform_L[74][2] = l_cell_wire[76];							inform_L[78][2] = l_cell_wire[77];							inform_L[75][2] = l_cell_wire[78];							inform_L[79][2] = l_cell_wire[79];							inform_L[80][2] = l_cell_wire[80];							inform_L[84][2] = l_cell_wire[81];							inform_L[81][2] = l_cell_wire[82];							inform_L[85][2] = l_cell_wire[83];							inform_L[82][2] = l_cell_wire[84];							inform_L[86][2] = l_cell_wire[85];							inform_L[83][2] = l_cell_wire[86];							inform_L[87][2] = l_cell_wire[87];							inform_L[88][2] = l_cell_wire[88];							inform_L[92][2] = l_cell_wire[89];							inform_L[89][2] = l_cell_wire[90];							inform_L[93][2] = l_cell_wire[91];							inform_L[90][2] = l_cell_wire[92];							inform_L[94][2] = l_cell_wire[93];							inform_L[91][2] = l_cell_wire[94];							inform_L[95][2] = l_cell_wire[95];							inform_L[96][2] = l_cell_wire[96];							inform_L[100][2] = l_cell_wire[97];							inform_L[97][2] = l_cell_wire[98];							inform_L[101][2] = l_cell_wire[99];							inform_L[98][2] = l_cell_wire[100];							inform_L[102][2] = l_cell_wire[101];							inform_L[99][2] = l_cell_wire[102];							inform_L[103][2] = l_cell_wire[103];							inform_L[104][2] = l_cell_wire[104];							inform_L[108][2] = l_cell_wire[105];							inform_L[105][2] = l_cell_wire[106];							inform_L[109][2] = l_cell_wire[107];							inform_L[106][2] = l_cell_wire[108];							inform_L[110][2] = l_cell_wire[109];							inform_L[107][2] = l_cell_wire[110];							inform_L[111][2] = l_cell_wire[111];							inform_L[112][2] = l_cell_wire[112];							inform_L[116][2] = l_cell_wire[113];							inform_L[113][2] = l_cell_wire[114];							inform_L[117][2] = l_cell_wire[115];							inform_L[114][2] = l_cell_wire[116];							inform_L[118][2] = l_cell_wire[117];							inform_L[115][2] = l_cell_wire[118];							inform_L[119][2] = l_cell_wire[119];							inform_L[120][2] = l_cell_wire[120];							inform_L[124][2] = l_cell_wire[121];							inform_L[121][2] = l_cell_wire[122];							inform_L[125][2] = l_cell_wire[123];							inform_L[122][2] = l_cell_wire[124];							inform_L[126][2] = l_cell_wire[125];							inform_L[123][2] = l_cell_wire[126];							inform_L[127][2] = l_cell_wire[127];							inform_L[128][2] = l_cell_wire[128];							inform_L[132][2] = l_cell_wire[129];							inform_L[129][2] = l_cell_wire[130];							inform_L[133][2] = l_cell_wire[131];							inform_L[130][2] = l_cell_wire[132];							inform_L[134][2] = l_cell_wire[133];							inform_L[131][2] = l_cell_wire[134];							inform_L[135][2] = l_cell_wire[135];							inform_L[136][2] = l_cell_wire[136];							inform_L[140][2] = l_cell_wire[137];							inform_L[137][2] = l_cell_wire[138];							inform_L[141][2] = l_cell_wire[139];							inform_L[138][2] = l_cell_wire[140];							inform_L[142][2] = l_cell_wire[141];							inform_L[139][2] = l_cell_wire[142];							inform_L[143][2] = l_cell_wire[143];							inform_L[144][2] = l_cell_wire[144];							inform_L[148][2] = l_cell_wire[145];							inform_L[145][2] = l_cell_wire[146];							inform_L[149][2] = l_cell_wire[147];							inform_L[146][2] = l_cell_wire[148];							inform_L[150][2] = l_cell_wire[149];							inform_L[147][2] = l_cell_wire[150];							inform_L[151][2] = l_cell_wire[151];							inform_L[152][2] = l_cell_wire[152];							inform_L[156][2] = l_cell_wire[153];							inform_L[153][2] = l_cell_wire[154];							inform_L[157][2] = l_cell_wire[155];							inform_L[154][2] = l_cell_wire[156];							inform_L[158][2] = l_cell_wire[157];							inform_L[155][2] = l_cell_wire[158];							inform_L[159][2] = l_cell_wire[159];							inform_L[160][2] = l_cell_wire[160];							inform_L[164][2] = l_cell_wire[161];							inform_L[161][2] = l_cell_wire[162];							inform_L[165][2] = l_cell_wire[163];							inform_L[162][2] = l_cell_wire[164];							inform_L[166][2] = l_cell_wire[165];							inform_L[163][2] = l_cell_wire[166];							inform_L[167][2] = l_cell_wire[167];							inform_L[168][2] = l_cell_wire[168];							inform_L[172][2] = l_cell_wire[169];							inform_L[169][2] = l_cell_wire[170];							inform_L[173][2] = l_cell_wire[171];							inform_L[170][2] = l_cell_wire[172];							inform_L[174][2] = l_cell_wire[173];							inform_L[171][2] = l_cell_wire[174];							inform_L[175][2] = l_cell_wire[175];							inform_L[176][2] = l_cell_wire[176];							inform_L[180][2] = l_cell_wire[177];							inform_L[177][2] = l_cell_wire[178];							inform_L[181][2] = l_cell_wire[179];							inform_L[178][2] = l_cell_wire[180];							inform_L[182][2] = l_cell_wire[181];							inform_L[179][2] = l_cell_wire[182];							inform_L[183][2] = l_cell_wire[183];							inform_L[184][2] = l_cell_wire[184];							inform_L[188][2] = l_cell_wire[185];							inform_L[185][2] = l_cell_wire[186];							inform_L[189][2] = l_cell_wire[187];							inform_L[186][2] = l_cell_wire[188];							inform_L[190][2] = l_cell_wire[189];							inform_L[187][2] = l_cell_wire[190];							inform_L[191][2] = l_cell_wire[191];							inform_L[192][2] = l_cell_wire[192];							inform_L[196][2] = l_cell_wire[193];							inform_L[193][2] = l_cell_wire[194];							inform_L[197][2] = l_cell_wire[195];							inform_L[194][2] = l_cell_wire[196];							inform_L[198][2] = l_cell_wire[197];							inform_L[195][2] = l_cell_wire[198];							inform_L[199][2] = l_cell_wire[199];							inform_L[200][2] = l_cell_wire[200];							inform_L[204][2] = l_cell_wire[201];							inform_L[201][2] = l_cell_wire[202];							inform_L[205][2] = l_cell_wire[203];							inform_L[202][2] = l_cell_wire[204];							inform_L[206][2] = l_cell_wire[205];							inform_L[203][2] = l_cell_wire[206];							inform_L[207][2] = l_cell_wire[207];							inform_L[208][2] = l_cell_wire[208];							inform_L[212][2] = l_cell_wire[209];							inform_L[209][2] = l_cell_wire[210];							inform_L[213][2] = l_cell_wire[211];							inform_L[210][2] = l_cell_wire[212];							inform_L[214][2] = l_cell_wire[213];							inform_L[211][2] = l_cell_wire[214];							inform_L[215][2] = l_cell_wire[215];							inform_L[216][2] = l_cell_wire[216];							inform_L[220][2] = l_cell_wire[217];							inform_L[217][2] = l_cell_wire[218];							inform_L[221][2] = l_cell_wire[219];							inform_L[218][2] = l_cell_wire[220];							inform_L[222][2] = l_cell_wire[221];							inform_L[219][2] = l_cell_wire[222];							inform_L[223][2] = l_cell_wire[223];							inform_L[224][2] = l_cell_wire[224];							inform_L[228][2] = l_cell_wire[225];							inform_L[225][2] = l_cell_wire[226];							inform_L[229][2] = l_cell_wire[227];							inform_L[226][2] = l_cell_wire[228];							inform_L[230][2] = l_cell_wire[229];							inform_L[227][2] = l_cell_wire[230];							inform_L[231][2] = l_cell_wire[231];							inform_L[232][2] = l_cell_wire[232];							inform_L[236][2] = l_cell_wire[233];							inform_L[233][2] = l_cell_wire[234];							inform_L[237][2] = l_cell_wire[235];							inform_L[234][2] = l_cell_wire[236];							inform_L[238][2] = l_cell_wire[237];							inform_L[235][2] = l_cell_wire[238];							inform_L[239][2] = l_cell_wire[239];							inform_L[240][2] = l_cell_wire[240];							inform_L[244][2] = l_cell_wire[241];							inform_L[241][2] = l_cell_wire[242];							inform_L[245][2] = l_cell_wire[243];							inform_L[242][2] = l_cell_wire[244];							inform_L[246][2] = l_cell_wire[245];							inform_L[243][2] = l_cell_wire[246];							inform_L[247][2] = l_cell_wire[247];							inform_L[248][2] = l_cell_wire[248];							inform_L[252][2] = l_cell_wire[249];							inform_L[249][2] = l_cell_wire[250];							inform_L[253][2] = l_cell_wire[251];							inform_L[250][2] = l_cell_wire[252];							inform_L[254][2] = l_cell_wire[253];							inform_L[251][2] = l_cell_wire[254];							inform_L[255][2] = l_cell_wire[255];						end
						4:						begin							inform_R[0][4] = r_cell_wire[0];							inform_R[8][4] = r_cell_wire[1];							inform_R[1][4] = r_cell_wire[2];							inform_R[9][4] = r_cell_wire[3];							inform_R[2][4] = r_cell_wire[4];							inform_R[10][4] = r_cell_wire[5];							inform_R[3][4] = r_cell_wire[6];							inform_R[11][4] = r_cell_wire[7];							inform_R[4][4] = r_cell_wire[8];							inform_R[12][4] = r_cell_wire[9];							inform_R[5][4] = r_cell_wire[10];							inform_R[13][4] = r_cell_wire[11];							inform_R[6][4] = r_cell_wire[12];							inform_R[14][4] = r_cell_wire[13];							inform_R[7][4] = r_cell_wire[14];							inform_R[15][4] = r_cell_wire[15];							inform_R[16][4] = r_cell_wire[16];							inform_R[24][4] = r_cell_wire[17];							inform_R[17][4] = r_cell_wire[18];							inform_R[25][4] = r_cell_wire[19];							inform_R[18][4] = r_cell_wire[20];							inform_R[26][4] = r_cell_wire[21];							inform_R[19][4] = r_cell_wire[22];							inform_R[27][4] = r_cell_wire[23];							inform_R[20][4] = r_cell_wire[24];							inform_R[28][4] = r_cell_wire[25];							inform_R[21][4] = r_cell_wire[26];							inform_R[29][4] = r_cell_wire[27];							inform_R[22][4] = r_cell_wire[28];							inform_R[30][4] = r_cell_wire[29];							inform_R[23][4] = r_cell_wire[30];							inform_R[31][4] = r_cell_wire[31];							inform_R[32][4] = r_cell_wire[32];							inform_R[40][4] = r_cell_wire[33];							inform_R[33][4] = r_cell_wire[34];							inform_R[41][4] = r_cell_wire[35];							inform_R[34][4] = r_cell_wire[36];							inform_R[42][4] = r_cell_wire[37];							inform_R[35][4] = r_cell_wire[38];							inform_R[43][4] = r_cell_wire[39];							inform_R[36][4] = r_cell_wire[40];							inform_R[44][4] = r_cell_wire[41];							inform_R[37][4] = r_cell_wire[42];							inform_R[45][4] = r_cell_wire[43];							inform_R[38][4] = r_cell_wire[44];							inform_R[46][4] = r_cell_wire[45];							inform_R[39][4] = r_cell_wire[46];							inform_R[47][4] = r_cell_wire[47];							inform_R[48][4] = r_cell_wire[48];							inform_R[56][4] = r_cell_wire[49];							inform_R[49][4] = r_cell_wire[50];							inform_R[57][4] = r_cell_wire[51];							inform_R[50][4] = r_cell_wire[52];							inform_R[58][4] = r_cell_wire[53];							inform_R[51][4] = r_cell_wire[54];							inform_R[59][4] = r_cell_wire[55];							inform_R[52][4] = r_cell_wire[56];							inform_R[60][4] = r_cell_wire[57];							inform_R[53][4] = r_cell_wire[58];							inform_R[61][4] = r_cell_wire[59];							inform_R[54][4] = r_cell_wire[60];							inform_R[62][4] = r_cell_wire[61];							inform_R[55][4] = r_cell_wire[62];							inform_R[63][4] = r_cell_wire[63];							inform_R[64][4] = r_cell_wire[64];							inform_R[72][4] = r_cell_wire[65];							inform_R[65][4] = r_cell_wire[66];							inform_R[73][4] = r_cell_wire[67];							inform_R[66][4] = r_cell_wire[68];							inform_R[74][4] = r_cell_wire[69];							inform_R[67][4] = r_cell_wire[70];							inform_R[75][4] = r_cell_wire[71];							inform_R[68][4] = r_cell_wire[72];							inform_R[76][4] = r_cell_wire[73];							inform_R[69][4] = r_cell_wire[74];							inform_R[77][4] = r_cell_wire[75];							inform_R[70][4] = r_cell_wire[76];							inform_R[78][4] = r_cell_wire[77];							inform_R[71][4] = r_cell_wire[78];							inform_R[79][4] = r_cell_wire[79];							inform_R[80][4] = r_cell_wire[80];							inform_R[88][4] = r_cell_wire[81];							inform_R[81][4] = r_cell_wire[82];							inform_R[89][4] = r_cell_wire[83];							inform_R[82][4] = r_cell_wire[84];							inform_R[90][4] = r_cell_wire[85];							inform_R[83][4] = r_cell_wire[86];							inform_R[91][4] = r_cell_wire[87];							inform_R[84][4] = r_cell_wire[88];							inform_R[92][4] = r_cell_wire[89];							inform_R[85][4] = r_cell_wire[90];							inform_R[93][4] = r_cell_wire[91];							inform_R[86][4] = r_cell_wire[92];							inform_R[94][4] = r_cell_wire[93];							inform_R[87][4] = r_cell_wire[94];							inform_R[95][4] = r_cell_wire[95];							inform_R[96][4] = r_cell_wire[96];							inform_R[104][4] = r_cell_wire[97];							inform_R[97][4] = r_cell_wire[98];							inform_R[105][4] = r_cell_wire[99];							inform_R[98][4] = r_cell_wire[100];							inform_R[106][4] = r_cell_wire[101];							inform_R[99][4] = r_cell_wire[102];							inform_R[107][4] = r_cell_wire[103];							inform_R[100][4] = r_cell_wire[104];							inform_R[108][4] = r_cell_wire[105];							inform_R[101][4] = r_cell_wire[106];							inform_R[109][4] = r_cell_wire[107];							inform_R[102][4] = r_cell_wire[108];							inform_R[110][4] = r_cell_wire[109];							inform_R[103][4] = r_cell_wire[110];							inform_R[111][4] = r_cell_wire[111];							inform_R[112][4] = r_cell_wire[112];							inform_R[120][4] = r_cell_wire[113];							inform_R[113][4] = r_cell_wire[114];							inform_R[121][4] = r_cell_wire[115];							inform_R[114][4] = r_cell_wire[116];							inform_R[122][4] = r_cell_wire[117];							inform_R[115][4] = r_cell_wire[118];							inform_R[123][4] = r_cell_wire[119];							inform_R[116][4] = r_cell_wire[120];							inform_R[124][4] = r_cell_wire[121];							inform_R[117][4] = r_cell_wire[122];							inform_R[125][4] = r_cell_wire[123];							inform_R[118][4] = r_cell_wire[124];							inform_R[126][4] = r_cell_wire[125];							inform_R[119][4] = r_cell_wire[126];							inform_R[127][4] = r_cell_wire[127];							inform_R[128][4] = r_cell_wire[128];							inform_R[136][4] = r_cell_wire[129];							inform_R[129][4] = r_cell_wire[130];							inform_R[137][4] = r_cell_wire[131];							inform_R[130][4] = r_cell_wire[132];							inform_R[138][4] = r_cell_wire[133];							inform_R[131][4] = r_cell_wire[134];							inform_R[139][4] = r_cell_wire[135];							inform_R[132][4] = r_cell_wire[136];							inform_R[140][4] = r_cell_wire[137];							inform_R[133][4] = r_cell_wire[138];							inform_R[141][4] = r_cell_wire[139];							inform_R[134][4] = r_cell_wire[140];							inform_R[142][4] = r_cell_wire[141];							inform_R[135][4] = r_cell_wire[142];							inform_R[143][4] = r_cell_wire[143];							inform_R[144][4] = r_cell_wire[144];							inform_R[152][4] = r_cell_wire[145];							inform_R[145][4] = r_cell_wire[146];							inform_R[153][4] = r_cell_wire[147];							inform_R[146][4] = r_cell_wire[148];							inform_R[154][4] = r_cell_wire[149];							inform_R[147][4] = r_cell_wire[150];							inform_R[155][4] = r_cell_wire[151];							inform_R[148][4] = r_cell_wire[152];							inform_R[156][4] = r_cell_wire[153];							inform_R[149][4] = r_cell_wire[154];							inform_R[157][4] = r_cell_wire[155];							inform_R[150][4] = r_cell_wire[156];							inform_R[158][4] = r_cell_wire[157];							inform_R[151][4] = r_cell_wire[158];							inform_R[159][4] = r_cell_wire[159];							inform_R[160][4] = r_cell_wire[160];							inform_R[168][4] = r_cell_wire[161];							inform_R[161][4] = r_cell_wire[162];							inform_R[169][4] = r_cell_wire[163];							inform_R[162][4] = r_cell_wire[164];							inform_R[170][4] = r_cell_wire[165];							inform_R[163][4] = r_cell_wire[166];							inform_R[171][4] = r_cell_wire[167];							inform_R[164][4] = r_cell_wire[168];							inform_R[172][4] = r_cell_wire[169];							inform_R[165][4] = r_cell_wire[170];							inform_R[173][4] = r_cell_wire[171];							inform_R[166][4] = r_cell_wire[172];							inform_R[174][4] = r_cell_wire[173];							inform_R[167][4] = r_cell_wire[174];							inform_R[175][4] = r_cell_wire[175];							inform_R[176][4] = r_cell_wire[176];							inform_R[184][4] = r_cell_wire[177];							inform_R[177][4] = r_cell_wire[178];							inform_R[185][4] = r_cell_wire[179];							inform_R[178][4] = r_cell_wire[180];							inform_R[186][4] = r_cell_wire[181];							inform_R[179][4] = r_cell_wire[182];							inform_R[187][4] = r_cell_wire[183];							inform_R[180][4] = r_cell_wire[184];							inform_R[188][4] = r_cell_wire[185];							inform_R[181][4] = r_cell_wire[186];							inform_R[189][4] = r_cell_wire[187];							inform_R[182][4] = r_cell_wire[188];							inform_R[190][4] = r_cell_wire[189];							inform_R[183][4] = r_cell_wire[190];							inform_R[191][4] = r_cell_wire[191];							inform_R[192][4] = r_cell_wire[192];							inform_R[200][4] = r_cell_wire[193];							inform_R[193][4] = r_cell_wire[194];							inform_R[201][4] = r_cell_wire[195];							inform_R[194][4] = r_cell_wire[196];							inform_R[202][4] = r_cell_wire[197];							inform_R[195][4] = r_cell_wire[198];							inform_R[203][4] = r_cell_wire[199];							inform_R[196][4] = r_cell_wire[200];							inform_R[204][4] = r_cell_wire[201];							inform_R[197][4] = r_cell_wire[202];							inform_R[205][4] = r_cell_wire[203];							inform_R[198][4] = r_cell_wire[204];							inform_R[206][4] = r_cell_wire[205];							inform_R[199][4] = r_cell_wire[206];							inform_R[207][4] = r_cell_wire[207];							inform_R[208][4] = r_cell_wire[208];							inform_R[216][4] = r_cell_wire[209];							inform_R[209][4] = r_cell_wire[210];							inform_R[217][4] = r_cell_wire[211];							inform_R[210][4] = r_cell_wire[212];							inform_R[218][4] = r_cell_wire[213];							inform_R[211][4] = r_cell_wire[214];							inform_R[219][4] = r_cell_wire[215];							inform_R[212][4] = r_cell_wire[216];							inform_R[220][4] = r_cell_wire[217];							inform_R[213][4] = r_cell_wire[218];							inform_R[221][4] = r_cell_wire[219];							inform_R[214][4] = r_cell_wire[220];							inform_R[222][4] = r_cell_wire[221];							inform_R[215][4] = r_cell_wire[222];							inform_R[223][4] = r_cell_wire[223];							inform_R[224][4] = r_cell_wire[224];							inform_R[232][4] = r_cell_wire[225];							inform_R[225][4] = r_cell_wire[226];							inform_R[233][4] = r_cell_wire[227];							inform_R[226][4] = r_cell_wire[228];							inform_R[234][4] = r_cell_wire[229];							inform_R[227][4] = r_cell_wire[230];							inform_R[235][4] = r_cell_wire[231];							inform_R[228][4] = r_cell_wire[232];							inform_R[236][4] = r_cell_wire[233];							inform_R[229][4] = r_cell_wire[234];							inform_R[237][4] = r_cell_wire[235];							inform_R[230][4] = r_cell_wire[236];							inform_R[238][4] = r_cell_wire[237];							inform_R[231][4] = r_cell_wire[238];							inform_R[239][4] = r_cell_wire[239];							inform_R[240][4] = r_cell_wire[240];							inform_R[248][4] = r_cell_wire[241];							inform_R[241][4] = r_cell_wire[242];							inform_R[249][4] = r_cell_wire[243];							inform_R[242][4] = r_cell_wire[244];							inform_R[250][4] = r_cell_wire[245];							inform_R[243][4] = r_cell_wire[246];							inform_R[251][4] = r_cell_wire[247];							inform_R[244][4] = r_cell_wire[248];							inform_R[252][4] = r_cell_wire[249];							inform_R[245][4] = r_cell_wire[250];							inform_R[253][4] = r_cell_wire[251];							inform_R[246][4] = r_cell_wire[252];							inform_R[254][4] = r_cell_wire[253];							inform_R[247][4] = r_cell_wire[254];							inform_R[255][4] = r_cell_wire[255];							inform_L[0][3] = l_cell_wire[0];							inform_L[8][3] = l_cell_wire[1];							inform_L[1][3] = l_cell_wire[2];							inform_L[9][3] = l_cell_wire[3];							inform_L[2][3] = l_cell_wire[4];							inform_L[10][3] = l_cell_wire[5];							inform_L[3][3] = l_cell_wire[6];							inform_L[11][3] = l_cell_wire[7];							inform_L[4][3] = l_cell_wire[8];							inform_L[12][3] = l_cell_wire[9];							inform_L[5][3] = l_cell_wire[10];							inform_L[13][3] = l_cell_wire[11];							inform_L[6][3] = l_cell_wire[12];							inform_L[14][3] = l_cell_wire[13];							inform_L[7][3] = l_cell_wire[14];							inform_L[15][3] = l_cell_wire[15];							inform_L[16][3] = l_cell_wire[16];							inform_L[24][3] = l_cell_wire[17];							inform_L[17][3] = l_cell_wire[18];							inform_L[25][3] = l_cell_wire[19];							inform_L[18][3] = l_cell_wire[20];							inform_L[26][3] = l_cell_wire[21];							inform_L[19][3] = l_cell_wire[22];							inform_L[27][3] = l_cell_wire[23];							inform_L[20][3] = l_cell_wire[24];							inform_L[28][3] = l_cell_wire[25];							inform_L[21][3] = l_cell_wire[26];							inform_L[29][3] = l_cell_wire[27];							inform_L[22][3] = l_cell_wire[28];							inform_L[30][3] = l_cell_wire[29];							inform_L[23][3] = l_cell_wire[30];							inform_L[31][3] = l_cell_wire[31];							inform_L[32][3] = l_cell_wire[32];							inform_L[40][3] = l_cell_wire[33];							inform_L[33][3] = l_cell_wire[34];							inform_L[41][3] = l_cell_wire[35];							inform_L[34][3] = l_cell_wire[36];							inform_L[42][3] = l_cell_wire[37];							inform_L[35][3] = l_cell_wire[38];							inform_L[43][3] = l_cell_wire[39];							inform_L[36][3] = l_cell_wire[40];							inform_L[44][3] = l_cell_wire[41];							inform_L[37][3] = l_cell_wire[42];							inform_L[45][3] = l_cell_wire[43];							inform_L[38][3] = l_cell_wire[44];							inform_L[46][3] = l_cell_wire[45];							inform_L[39][3] = l_cell_wire[46];							inform_L[47][3] = l_cell_wire[47];							inform_L[48][3] = l_cell_wire[48];							inform_L[56][3] = l_cell_wire[49];							inform_L[49][3] = l_cell_wire[50];							inform_L[57][3] = l_cell_wire[51];							inform_L[50][3] = l_cell_wire[52];							inform_L[58][3] = l_cell_wire[53];							inform_L[51][3] = l_cell_wire[54];							inform_L[59][3] = l_cell_wire[55];							inform_L[52][3] = l_cell_wire[56];							inform_L[60][3] = l_cell_wire[57];							inform_L[53][3] = l_cell_wire[58];							inform_L[61][3] = l_cell_wire[59];							inform_L[54][3] = l_cell_wire[60];							inform_L[62][3] = l_cell_wire[61];							inform_L[55][3] = l_cell_wire[62];							inform_L[63][3] = l_cell_wire[63];							inform_L[64][3] = l_cell_wire[64];							inform_L[72][3] = l_cell_wire[65];							inform_L[65][3] = l_cell_wire[66];							inform_L[73][3] = l_cell_wire[67];							inform_L[66][3] = l_cell_wire[68];							inform_L[74][3] = l_cell_wire[69];							inform_L[67][3] = l_cell_wire[70];							inform_L[75][3] = l_cell_wire[71];							inform_L[68][3] = l_cell_wire[72];							inform_L[76][3] = l_cell_wire[73];							inform_L[69][3] = l_cell_wire[74];							inform_L[77][3] = l_cell_wire[75];							inform_L[70][3] = l_cell_wire[76];							inform_L[78][3] = l_cell_wire[77];							inform_L[71][3] = l_cell_wire[78];							inform_L[79][3] = l_cell_wire[79];							inform_L[80][3] = l_cell_wire[80];							inform_L[88][3] = l_cell_wire[81];							inform_L[81][3] = l_cell_wire[82];							inform_L[89][3] = l_cell_wire[83];							inform_L[82][3] = l_cell_wire[84];							inform_L[90][3] = l_cell_wire[85];							inform_L[83][3] = l_cell_wire[86];							inform_L[91][3] = l_cell_wire[87];							inform_L[84][3] = l_cell_wire[88];							inform_L[92][3] = l_cell_wire[89];							inform_L[85][3] = l_cell_wire[90];							inform_L[93][3] = l_cell_wire[91];							inform_L[86][3] = l_cell_wire[92];							inform_L[94][3] = l_cell_wire[93];							inform_L[87][3] = l_cell_wire[94];							inform_L[95][3] = l_cell_wire[95];							inform_L[96][3] = l_cell_wire[96];							inform_L[104][3] = l_cell_wire[97];							inform_L[97][3] = l_cell_wire[98];							inform_L[105][3] = l_cell_wire[99];							inform_L[98][3] = l_cell_wire[100];							inform_L[106][3] = l_cell_wire[101];							inform_L[99][3] = l_cell_wire[102];							inform_L[107][3] = l_cell_wire[103];							inform_L[100][3] = l_cell_wire[104];							inform_L[108][3] = l_cell_wire[105];							inform_L[101][3] = l_cell_wire[106];							inform_L[109][3] = l_cell_wire[107];							inform_L[102][3] = l_cell_wire[108];							inform_L[110][3] = l_cell_wire[109];							inform_L[103][3] = l_cell_wire[110];							inform_L[111][3] = l_cell_wire[111];							inform_L[112][3] = l_cell_wire[112];							inform_L[120][3] = l_cell_wire[113];							inform_L[113][3] = l_cell_wire[114];							inform_L[121][3] = l_cell_wire[115];							inform_L[114][3] = l_cell_wire[116];							inform_L[122][3] = l_cell_wire[117];							inform_L[115][3] = l_cell_wire[118];							inform_L[123][3] = l_cell_wire[119];							inform_L[116][3] = l_cell_wire[120];							inform_L[124][3] = l_cell_wire[121];							inform_L[117][3] = l_cell_wire[122];							inform_L[125][3] = l_cell_wire[123];							inform_L[118][3] = l_cell_wire[124];							inform_L[126][3] = l_cell_wire[125];							inform_L[119][3] = l_cell_wire[126];							inform_L[127][3] = l_cell_wire[127];							inform_L[128][3] = l_cell_wire[128];							inform_L[136][3] = l_cell_wire[129];							inform_L[129][3] = l_cell_wire[130];							inform_L[137][3] = l_cell_wire[131];							inform_L[130][3] = l_cell_wire[132];							inform_L[138][3] = l_cell_wire[133];							inform_L[131][3] = l_cell_wire[134];							inform_L[139][3] = l_cell_wire[135];							inform_L[132][3] = l_cell_wire[136];							inform_L[140][3] = l_cell_wire[137];							inform_L[133][3] = l_cell_wire[138];							inform_L[141][3] = l_cell_wire[139];							inform_L[134][3] = l_cell_wire[140];							inform_L[142][3] = l_cell_wire[141];							inform_L[135][3] = l_cell_wire[142];							inform_L[143][3] = l_cell_wire[143];							inform_L[144][3] = l_cell_wire[144];							inform_L[152][3] = l_cell_wire[145];							inform_L[145][3] = l_cell_wire[146];							inform_L[153][3] = l_cell_wire[147];							inform_L[146][3] = l_cell_wire[148];							inform_L[154][3] = l_cell_wire[149];							inform_L[147][3] = l_cell_wire[150];							inform_L[155][3] = l_cell_wire[151];							inform_L[148][3] = l_cell_wire[152];							inform_L[156][3] = l_cell_wire[153];							inform_L[149][3] = l_cell_wire[154];							inform_L[157][3] = l_cell_wire[155];							inform_L[150][3] = l_cell_wire[156];							inform_L[158][3] = l_cell_wire[157];							inform_L[151][3] = l_cell_wire[158];							inform_L[159][3] = l_cell_wire[159];							inform_L[160][3] = l_cell_wire[160];							inform_L[168][3] = l_cell_wire[161];							inform_L[161][3] = l_cell_wire[162];							inform_L[169][3] = l_cell_wire[163];							inform_L[162][3] = l_cell_wire[164];							inform_L[170][3] = l_cell_wire[165];							inform_L[163][3] = l_cell_wire[166];							inform_L[171][3] = l_cell_wire[167];							inform_L[164][3] = l_cell_wire[168];							inform_L[172][3] = l_cell_wire[169];							inform_L[165][3] = l_cell_wire[170];							inform_L[173][3] = l_cell_wire[171];							inform_L[166][3] = l_cell_wire[172];							inform_L[174][3] = l_cell_wire[173];							inform_L[167][3] = l_cell_wire[174];							inform_L[175][3] = l_cell_wire[175];							inform_L[176][3] = l_cell_wire[176];							inform_L[184][3] = l_cell_wire[177];							inform_L[177][3] = l_cell_wire[178];							inform_L[185][3] = l_cell_wire[179];							inform_L[178][3] = l_cell_wire[180];							inform_L[186][3] = l_cell_wire[181];							inform_L[179][3] = l_cell_wire[182];							inform_L[187][3] = l_cell_wire[183];							inform_L[180][3] = l_cell_wire[184];							inform_L[188][3] = l_cell_wire[185];							inform_L[181][3] = l_cell_wire[186];							inform_L[189][3] = l_cell_wire[187];							inform_L[182][3] = l_cell_wire[188];							inform_L[190][3] = l_cell_wire[189];							inform_L[183][3] = l_cell_wire[190];							inform_L[191][3] = l_cell_wire[191];							inform_L[192][3] = l_cell_wire[192];							inform_L[200][3] = l_cell_wire[193];							inform_L[193][3] = l_cell_wire[194];							inform_L[201][3] = l_cell_wire[195];							inform_L[194][3] = l_cell_wire[196];							inform_L[202][3] = l_cell_wire[197];							inform_L[195][3] = l_cell_wire[198];							inform_L[203][3] = l_cell_wire[199];							inform_L[196][3] = l_cell_wire[200];							inform_L[204][3] = l_cell_wire[201];							inform_L[197][3] = l_cell_wire[202];							inform_L[205][3] = l_cell_wire[203];							inform_L[198][3] = l_cell_wire[204];							inform_L[206][3] = l_cell_wire[205];							inform_L[199][3] = l_cell_wire[206];							inform_L[207][3] = l_cell_wire[207];							inform_L[208][3] = l_cell_wire[208];							inform_L[216][3] = l_cell_wire[209];							inform_L[209][3] = l_cell_wire[210];							inform_L[217][3] = l_cell_wire[211];							inform_L[210][3] = l_cell_wire[212];							inform_L[218][3] = l_cell_wire[213];							inform_L[211][3] = l_cell_wire[214];							inform_L[219][3] = l_cell_wire[215];							inform_L[212][3] = l_cell_wire[216];							inform_L[220][3] = l_cell_wire[217];							inform_L[213][3] = l_cell_wire[218];							inform_L[221][3] = l_cell_wire[219];							inform_L[214][3] = l_cell_wire[220];							inform_L[222][3] = l_cell_wire[221];							inform_L[215][3] = l_cell_wire[222];							inform_L[223][3] = l_cell_wire[223];							inform_L[224][3] = l_cell_wire[224];							inform_L[232][3] = l_cell_wire[225];							inform_L[225][3] = l_cell_wire[226];							inform_L[233][3] = l_cell_wire[227];							inform_L[226][3] = l_cell_wire[228];							inform_L[234][3] = l_cell_wire[229];							inform_L[227][3] = l_cell_wire[230];							inform_L[235][3] = l_cell_wire[231];							inform_L[228][3] = l_cell_wire[232];							inform_L[236][3] = l_cell_wire[233];							inform_L[229][3] = l_cell_wire[234];							inform_L[237][3] = l_cell_wire[235];							inform_L[230][3] = l_cell_wire[236];							inform_L[238][3] = l_cell_wire[237];							inform_L[231][3] = l_cell_wire[238];							inform_L[239][3] = l_cell_wire[239];							inform_L[240][3] = l_cell_wire[240];							inform_L[248][3] = l_cell_wire[241];							inform_L[241][3] = l_cell_wire[242];							inform_L[249][3] = l_cell_wire[243];							inform_L[242][3] = l_cell_wire[244];							inform_L[250][3] = l_cell_wire[245];							inform_L[243][3] = l_cell_wire[246];							inform_L[251][3] = l_cell_wire[247];							inform_L[244][3] = l_cell_wire[248];							inform_L[252][3] = l_cell_wire[249];							inform_L[245][3] = l_cell_wire[250];							inform_L[253][3] = l_cell_wire[251];							inform_L[246][3] = l_cell_wire[252];							inform_L[254][3] = l_cell_wire[253];							inform_L[247][3] = l_cell_wire[254];							inform_L[255][3] = l_cell_wire[255];						end
						5:						begin							inform_R[0][5] = r_cell_wire[0];							inform_R[16][5] = r_cell_wire[1];							inform_R[1][5] = r_cell_wire[2];							inform_R[17][5] = r_cell_wire[3];							inform_R[2][5] = r_cell_wire[4];							inform_R[18][5] = r_cell_wire[5];							inform_R[3][5] = r_cell_wire[6];							inform_R[19][5] = r_cell_wire[7];							inform_R[4][5] = r_cell_wire[8];							inform_R[20][5] = r_cell_wire[9];							inform_R[5][5] = r_cell_wire[10];							inform_R[21][5] = r_cell_wire[11];							inform_R[6][5] = r_cell_wire[12];							inform_R[22][5] = r_cell_wire[13];							inform_R[7][5] = r_cell_wire[14];							inform_R[23][5] = r_cell_wire[15];							inform_R[8][5] = r_cell_wire[16];							inform_R[24][5] = r_cell_wire[17];							inform_R[9][5] = r_cell_wire[18];							inform_R[25][5] = r_cell_wire[19];							inform_R[10][5] = r_cell_wire[20];							inform_R[26][5] = r_cell_wire[21];							inform_R[11][5] = r_cell_wire[22];							inform_R[27][5] = r_cell_wire[23];							inform_R[12][5] = r_cell_wire[24];							inform_R[28][5] = r_cell_wire[25];							inform_R[13][5] = r_cell_wire[26];							inform_R[29][5] = r_cell_wire[27];							inform_R[14][5] = r_cell_wire[28];							inform_R[30][5] = r_cell_wire[29];							inform_R[15][5] = r_cell_wire[30];							inform_R[31][5] = r_cell_wire[31];							inform_R[32][5] = r_cell_wire[32];							inform_R[48][5] = r_cell_wire[33];							inform_R[33][5] = r_cell_wire[34];							inform_R[49][5] = r_cell_wire[35];							inform_R[34][5] = r_cell_wire[36];							inform_R[50][5] = r_cell_wire[37];							inform_R[35][5] = r_cell_wire[38];							inform_R[51][5] = r_cell_wire[39];							inform_R[36][5] = r_cell_wire[40];							inform_R[52][5] = r_cell_wire[41];							inform_R[37][5] = r_cell_wire[42];							inform_R[53][5] = r_cell_wire[43];							inform_R[38][5] = r_cell_wire[44];							inform_R[54][5] = r_cell_wire[45];							inform_R[39][5] = r_cell_wire[46];							inform_R[55][5] = r_cell_wire[47];							inform_R[40][5] = r_cell_wire[48];							inform_R[56][5] = r_cell_wire[49];							inform_R[41][5] = r_cell_wire[50];							inform_R[57][5] = r_cell_wire[51];							inform_R[42][5] = r_cell_wire[52];							inform_R[58][5] = r_cell_wire[53];							inform_R[43][5] = r_cell_wire[54];							inform_R[59][5] = r_cell_wire[55];							inform_R[44][5] = r_cell_wire[56];							inform_R[60][5] = r_cell_wire[57];							inform_R[45][5] = r_cell_wire[58];							inform_R[61][5] = r_cell_wire[59];							inform_R[46][5] = r_cell_wire[60];							inform_R[62][5] = r_cell_wire[61];							inform_R[47][5] = r_cell_wire[62];							inform_R[63][5] = r_cell_wire[63];							inform_R[64][5] = r_cell_wire[64];							inform_R[80][5] = r_cell_wire[65];							inform_R[65][5] = r_cell_wire[66];							inform_R[81][5] = r_cell_wire[67];							inform_R[66][5] = r_cell_wire[68];							inform_R[82][5] = r_cell_wire[69];							inform_R[67][5] = r_cell_wire[70];							inform_R[83][5] = r_cell_wire[71];							inform_R[68][5] = r_cell_wire[72];							inform_R[84][5] = r_cell_wire[73];							inform_R[69][5] = r_cell_wire[74];							inform_R[85][5] = r_cell_wire[75];							inform_R[70][5] = r_cell_wire[76];							inform_R[86][5] = r_cell_wire[77];							inform_R[71][5] = r_cell_wire[78];							inform_R[87][5] = r_cell_wire[79];							inform_R[72][5] = r_cell_wire[80];							inform_R[88][5] = r_cell_wire[81];							inform_R[73][5] = r_cell_wire[82];							inform_R[89][5] = r_cell_wire[83];							inform_R[74][5] = r_cell_wire[84];							inform_R[90][5] = r_cell_wire[85];							inform_R[75][5] = r_cell_wire[86];							inform_R[91][5] = r_cell_wire[87];							inform_R[76][5] = r_cell_wire[88];							inform_R[92][5] = r_cell_wire[89];							inform_R[77][5] = r_cell_wire[90];							inform_R[93][5] = r_cell_wire[91];							inform_R[78][5] = r_cell_wire[92];							inform_R[94][5] = r_cell_wire[93];							inform_R[79][5] = r_cell_wire[94];							inform_R[95][5] = r_cell_wire[95];							inform_R[96][5] = r_cell_wire[96];							inform_R[112][5] = r_cell_wire[97];							inform_R[97][5] = r_cell_wire[98];							inform_R[113][5] = r_cell_wire[99];							inform_R[98][5] = r_cell_wire[100];							inform_R[114][5] = r_cell_wire[101];							inform_R[99][5] = r_cell_wire[102];							inform_R[115][5] = r_cell_wire[103];							inform_R[100][5] = r_cell_wire[104];							inform_R[116][5] = r_cell_wire[105];							inform_R[101][5] = r_cell_wire[106];							inform_R[117][5] = r_cell_wire[107];							inform_R[102][5] = r_cell_wire[108];							inform_R[118][5] = r_cell_wire[109];							inform_R[103][5] = r_cell_wire[110];							inform_R[119][5] = r_cell_wire[111];							inform_R[104][5] = r_cell_wire[112];							inform_R[120][5] = r_cell_wire[113];							inform_R[105][5] = r_cell_wire[114];							inform_R[121][5] = r_cell_wire[115];							inform_R[106][5] = r_cell_wire[116];							inform_R[122][5] = r_cell_wire[117];							inform_R[107][5] = r_cell_wire[118];							inform_R[123][5] = r_cell_wire[119];							inform_R[108][5] = r_cell_wire[120];							inform_R[124][5] = r_cell_wire[121];							inform_R[109][5] = r_cell_wire[122];							inform_R[125][5] = r_cell_wire[123];							inform_R[110][5] = r_cell_wire[124];							inform_R[126][5] = r_cell_wire[125];							inform_R[111][5] = r_cell_wire[126];							inform_R[127][5] = r_cell_wire[127];							inform_R[128][5] = r_cell_wire[128];							inform_R[144][5] = r_cell_wire[129];							inform_R[129][5] = r_cell_wire[130];							inform_R[145][5] = r_cell_wire[131];							inform_R[130][5] = r_cell_wire[132];							inform_R[146][5] = r_cell_wire[133];							inform_R[131][5] = r_cell_wire[134];							inform_R[147][5] = r_cell_wire[135];							inform_R[132][5] = r_cell_wire[136];							inform_R[148][5] = r_cell_wire[137];							inform_R[133][5] = r_cell_wire[138];							inform_R[149][5] = r_cell_wire[139];							inform_R[134][5] = r_cell_wire[140];							inform_R[150][5] = r_cell_wire[141];							inform_R[135][5] = r_cell_wire[142];							inform_R[151][5] = r_cell_wire[143];							inform_R[136][5] = r_cell_wire[144];							inform_R[152][5] = r_cell_wire[145];							inform_R[137][5] = r_cell_wire[146];							inform_R[153][5] = r_cell_wire[147];							inform_R[138][5] = r_cell_wire[148];							inform_R[154][5] = r_cell_wire[149];							inform_R[139][5] = r_cell_wire[150];							inform_R[155][5] = r_cell_wire[151];							inform_R[140][5] = r_cell_wire[152];							inform_R[156][5] = r_cell_wire[153];							inform_R[141][5] = r_cell_wire[154];							inform_R[157][5] = r_cell_wire[155];							inform_R[142][5] = r_cell_wire[156];							inform_R[158][5] = r_cell_wire[157];							inform_R[143][5] = r_cell_wire[158];							inform_R[159][5] = r_cell_wire[159];							inform_R[160][5] = r_cell_wire[160];							inform_R[176][5] = r_cell_wire[161];							inform_R[161][5] = r_cell_wire[162];							inform_R[177][5] = r_cell_wire[163];							inform_R[162][5] = r_cell_wire[164];							inform_R[178][5] = r_cell_wire[165];							inform_R[163][5] = r_cell_wire[166];							inform_R[179][5] = r_cell_wire[167];							inform_R[164][5] = r_cell_wire[168];							inform_R[180][5] = r_cell_wire[169];							inform_R[165][5] = r_cell_wire[170];							inform_R[181][5] = r_cell_wire[171];							inform_R[166][5] = r_cell_wire[172];							inform_R[182][5] = r_cell_wire[173];							inform_R[167][5] = r_cell_wire[174];							inform_R[183][5] = r_cell_wire[175];							inform_R[168][5] = r_cell_wire[176];							inform_R[184][5] = r_cell_wire[177];							inform_R[169][5] = r_cell_wire[178];							inform_R[185][5] = r_cell_wire[179];							inform_R[170][5] = r_cell_wire[180];							inform_R[186][5] = r_cell_wire[181];							inform_R[171][5] = r_cell_wire[182];							inform_R[187][5] = r_cell_wire[183];							inform_R[172][5] = r_cell_wire[184];							inform_R[188][5] = r_cell_wire[185];							inform_R[173][5] = r_cell_wire[186];							inform_R[189][5] = r_cell_wire[187];							inform_R[174][5] = r_cell_wire[188];							inform_R[190][5] = r_cell_wire[189];							inform_R[175][5] = r_cell_wire[190];							inform_R[191][5] = r_cell_wire[191];							inform_R[192][5] = r_cell_wire[192];							inform_R[208][5] = r_cell_wire[193];							inform_R[193][5] = r_cell_wire[194];							inform_R[209][5] = r_cell_wire[195];							inform_R[194][5] = r_cell_wire[196];							inform_R[210][5] = r_cell_wire[197];							inform_R[195][5] = r_cell_wire[198];							inform_R[211][5] = r_cell_wire[199];							inform_R[196][5] = r_cell_wire[200];							inform_R[212][5] = r_cell_wire[201];							inform_R[197][5] = r_cell_wire[202];							inform_R[213][5] = r_cell_wire[203];							inform_R[198][5] = r_cell_wire[204];							inform_R[214][5] = r_cell_wire[205];							inform_R[199][5] = r_cell_wire[206];							inform_R[215][5] = r_cell_wire[207];							inform_R[200][5] = r_cell_wire[208];							inform_R[216][5] = r_cell_wire[209];							inform_R[201][5] = r_cell_wire[210];							inform_R[217][5] = r_cell_wire[211];							inform_R[202][5] = r_cell_wire[212];							inform_R[218][5] = r_cell_wire[213];							inform_R[203][5] = r_cell_wire[214];							inform_R[219][5] = r_cell_wire[215];							inform_R[204][5] = r_cell_wire[216];							inform_R[220][5] = r_cell_wire[217];							inform_R[205][5] = r_cell_wire[218];							inform_R[221][5] = r_cell_wire[219];							inform_R[206][5] = r_cell_wire[220];							inform_R[222][5] = r_cell_wire[221];							inform_R[207][5] = r_cell_wire[222];							inform_R[223][5] = r_cell_wire[223];							inform_R[224][5] = r_cell_wire[224];							inform_R[240][5] = r_cell_wire[225];							inform_R[225][5] = r_cell_wire[226];							inform_R[241][5] = r_cell_wire[227];							inform_R[226][5] = r_cell_wire[228];							inform_R[242][5] = r_cell_wire[229];							inform_R[227][5] = r_cell_wire[230];							inform_R[243][5] = r_cell_wire[231];							inform_R[228][5] = r_cell_wire[232];							inform_R[244][5] = r_cell_wire[233];							inform_R[229][5] = r_cell_wire[234];							inform_R[245][5] = r_cell_wire[235];							inform_R[230][5] = r_cell_wire[236];							inform_R[246][5] = r_cell_wire[237];							inform_R[231][5] = r_cell_wire[238];							inform_R[247][5] = r_cell_wire[239];							inform_R[232][5] = r_cell_wire[240];							inform_R[248][5] = r_cell_wire[241];							inform_R[233][5] = r_cell_wire[242];							inform_R[249][5] = r_cell_wire[243];							inform_R[234][5] = r_cell_wire[244];							inform_R[250][5] = r_cell_wire[245];							inform_R[235][5] = r_cell_wire[246];							inform_R[251][5] = r_cell_wire[247];							inform_R[236][5] = r_cell_wire[248];							inform_R[252][5] = r_cell_wire[249];							inform_R[237][5] = r_cell_wire[250];							inform_R[253][5] = r_cell_wire[251];							inform_R[238][5] = r_cell_wire[252];							inform_R[254][5] = r_cell_wire[253];							inform_R[239][5] = r_cell_wire[254];							inform_R[255][5] = r_cell_wire[255];							inform_L[0][4] = l_cell_wire[0];							inform_L[16][4] = l_cell_wire[1];							inform_L[1][4] = l_cell_wire[2];							inform_L[17][4] = l_cell_wire[3];							inform_L[2][4] = l_cell_wire[4];							inform_L[18][4] = l_cell_wire[5];							inform_L[3][4] = l_cell_wire[6];							inform_L[19][4] = l_cell_wire[7];							inform_L[4][4] = l_cell_wire[8];							inform_L[20][4] = l_cell_wire[9];							inform_L[5][4] = l_cell_wire[10];							inform_L[21][4] = l_cell_wire[11];							inform_L[6][4] = l_cell_wire[12];							inform_L[22][4] = l_cell_wire[13];							inform_L[7][4] = l_cell_wire[14];							inform_L[23][4] = l_cell_wire[15];							inform_L[8][4] = l_cell_wire[16];							inform_L[24][4] = l_cell_wire[17];							inform_L[9][4] = l_cell_wire[18];							inform_L[25][4] = l_cell_wire[19];							inform_L[10][4] = l_cell_wire[20];							inform_L[26][4] = l_cell_wire[21];							inform_L[11][4] = l_cell_wire[22];							inform_L[27][4] = l_cell_wire[23];							inform_L[12][4] = l_cell_wire[24];							inform_L[28][4] = l_cell_wire[25];							inform_L[13][4] = l_cell_wire[26];							inform_L[29][4] = l_cell_wire[27];							inform_L[14][4] = l_cell_wire[28];							inform_L[30][4] = l_cell_wire[29];							inform_L[15][4] = l_cell_wire[30];							inform_L[31][4] = l_cell_wire[31];							inform_L[32][4] = l_cell_wire[32];							inform_L[48][4] = l_cell_wire[33];							inform_L[33][4] = l_cell_wire[34];							inform_L[49][4] = l_cell_wire[35];							inform_L[34][4] = l_cell_wire[36];							inform_L[50][4] = l_cell_wire[37];							inform_L[35][4] = l_cell_wire[38];							inform_L[51][4] = l_cell_wire[39];							inform_L[36][4] = l_cell_wire[40];							inform_L[52][4] = l_cell_wire[41];							inform_L[37][4] = l_cell_wire[42];							inform_L[53][4] = l_cell_wire[43];							inform_L[38][4] = l_cell_wire[44];							inform_L[54][4] = l_cell_wire[45];							inform_L[39][4] = l_cell_wire[46];							inform_L[55][4] = l_cell_wire[47];							inform_L[40][4] = l_cell_wire[48];							inform_L[56][4] = l_cell_wire[49];							inform_L[41][4] = l_cell_wire[50];							inform_L[57][4] = l_cell_wire[51];							inform_L[42][4] = l_cell_wire[52];							inform_L[58][4] = l_cell_wire[53];							inform_L[43][4] = l_cell_wire[54];							inform_L[59][4] = l_cell_wire[55];							inform_L[44][4] = l_cell_wire[56];							inform_L[60][4] = l_cell_wire[57];							inform_L[45][4] = l_cell_wire[58];							inform_L[61][4] = l_cell_wire[59];							inform_L[46][4] = l_cell_wire[60];							inform_L[62][4] = l_cell_wire[61];							inform_L[47][4] = l_cell_wire[62];							inform_L[63][4] = l_cell_wire[63];							inform_L[64][4] = l_cell_wire[64];							inform_L[80][4] = l_cell_wire[65];							inform_L[65][4] = l_cell_wire[66];							inform_L[81][4] = l_cell_wire[67];							inform_L[66][4] = l_cell_wire[68];							inform_L[82][4] = l_cell_wire[69];							inform_L[67][4] = l_cell_wire[70];							inform_L[83][4] = l_cell_wire[71];							inform_L[68][4] = l_cell_wire[72];							inform_L[84][4] = l_cell_wire[73];							inform_L[69][4] = l_cell_wire[74];							inform_L[85][4] = l_cell_wire[75];							inform_L[70][4] = l_cell_wire[76];							inform_L[86][4] = l_cell_wire[77];							inform_L[71][4] = l_cell_wire[78];							inform_L[87][4] = l_cell_wire[79];							inform_L[72][4] = l_cell_wire[80];							inform_L[88][4] = l_cell_wire[81];							inform_L[73][4] = l_cell_wire[82];							inform_L[89][4] = l_cell_wire[83];							inform_L[74][4] = l_cell_wire[84];							inform_L[90][4] = l_cell_wire[85];							inform_L[75][4] = l_cell_wire[86];							inform_L[91][4] = l_cell_wire[87];							inform_L[76][4] = l_cell_wire[88];							inform_L[92][4] = l_cell_wire[89];							inform_L[77][4] = l_cell_wire[90];							inform_L[93][4] = l_cell_wire[91];							inform_L[78][4] = l_cell_wire[92];							inform_L[94][4] = l_cell_wire[93];							inform_L[79][4] = l_cell_wire[94];							inform_L[95][4] = l_cell_wire[95];							inform_L[96][4] = l_cell_wire[96];							inform_L[112][4] = l_cell_wire[97];							inform_L[97][4] = l_cell_wire[98];							inform_L[113][4] = l_cell_wire[99];							inform_L[98][4] = l_cell_wire[100];							inform_L[114][4] = l_cell_wire[101];							inform_L[99][4] = l_cell_wire[102];							inform_L[115][4] = l_cell_wire[103];							inform_L[100][4] = l_cell_wire[104];							inform_L[116][4] = l_cell_wire[105];							inform_L[101][4] = l_cell_wire[106];							inform_L[117][4] = l_cell_wire[107];							inform_L[102][4] = l_cell_wire[108];							inform_L[118][4] = l_cell_wire[109];							inform_L[103][4] = l_cell_wire[110];							inform_L[119][4] = l_cell_wire[111];							inform_L[104][4] = l_cell_wire[112];							inform_L[120][4] = l_cell_wire[113];							inform_L[105][4] = l_cell_wire[114];							inform_L[121][4] = l_cell_wire[115];							inform_L[106][4] = l_cell_wire[116];							inform_L[122][4] = l_cell_wire[117];							inform_L[107][4] = l_cell_wire[118];							inform_L[123][4] = l_cell_wire[119];							inform_L[108][4] = l_cell_wire[120];							inform_L[124][4] = l_cell_wire[121];							inform_L[109][4] = l_cell_wire[122];							inform_L[125][4] = l_cell_wire[123];							inform_L[110][4] = l_cell_wire[124];							inform_L[126][4] = l_cell_wire[125];							inform_L[111][4] = l_cell_wire[126];							inform_L[127][4] = l_cell_wire[127];							inform_L[128][4] = l_cell_wire[128];							inform_L[144][4] = l_cell_wire[129];							inform_L[129][4] = l_cell_wire[130];							inform_L[145][4] = l_cell_wire[131];							inform_L[130][4] = l_cell_wire[132];							inform_L[146][4] = l_cell_wire[133];							inform_L[131][4] = l_cell_wire[134];							inform_L[147][4] = l_cell_wire[135];							inform_L[132][4] = l_cell_wire[136];							inform_L[148][4] = l_cell_wire[137];							inform_L[133][4] = l_cell_wire[138];							inform_L[149][4] = l_cell_wire[139];							inform_L[134][4] = l_cell_wire[140];							inform_L[150][4] = l_cell_wire[141];							inform_L[135][4] = l_cell_wire[142];							inform_L[151][4] = l_cell_wire[143];							inform_L[136][4] = l_cell_wire[144];							inform_L[152][4] = l_cell_wire[145];							inform_L[137][4] = l_cell_wire[146];							inform_L[153][4] = l_cell_wire[147];							inform_L[138][4] = l_cell_wire[148];							inform_L[154][4] = l_cell_wire[149];							inform_L[139][4] = l_cell_wire[150];							inform_L[155][4] = l_cell_wire[151];							inform_L[140][4] = l_cell_wire[152];							inform_L[156][4] = l_cell_wire[153];							inform_L[141][4] = l_cell_wire[154];							inform_L[157][4] = l_cell_wire[155];							inform_L[142][4] = l_cell_wire[156];							inform_L[158][4] = l_cell_wire[157];							inform_L[143][4] = l_cell_wire[158];							inform_L[159][4] = l_cell_wire[159];							inform_L[160][4] = l_cell_wire[160];							inform_L[176][4] = l_cell_wire[161];							inform_L[161][4] = l_cell_wire[162];							inform_L[177][4] = l_cell_wire[163];							inform_L[162][4] = l_cell_wire[164];							inform_L[178][4] = l_cell_wire[165];							inform_L[163][4] = l_cell_wire[166];							inform_L[179][4] = l_cell_wire[167];							inform_L[164][4] = l_cell_wire[168];							inform_L[180][4] = l_cell_wire[169];							inform_L[165][4] = l_cell_wire[170];							inform_L[181][4] = l_cell_wire[171];							inform_L[166][4] = l_cell_wire[172];							inform_L[182][4] = l_cell_wire[173];							inform_L[167][4] = l_cell_wire[174];							inform_L[183][4] = l_cell_wire[175];							inform_L[168][4] = l_cell_wire[176];							inform_L[184][4] = l_cell_wire[177];							inform_L[169][4] = l_cell_wire[178];							inform_L[185][4] = l_cell_wire[179];							inform_L[170][4] = l_cell_wire[180];							inform_L[186][4] = l_cell_wire[181];							inform_L[171][4] = l_cell_wire[182];							inform_L[187][4] = l_cell_wire[183];							inform_L[172][4] = l_cell_wire[184];							inform_L[188][4] = l_cell_wire[185];							inform_L[173][4] = l_cell_wire[186];							inform_L[189][4] = l_cell_wire[187];							inform_L[174][4] = l_cell_wire[188];							inform_L[190][4] = l_cell_wire[189];							inform_L[175][4] = l_cell_wire[190];							inform_L[191][4] = l_cell_wire[191];							inform_L[192][4] = l_cell_wire[192];							inform_L[208][4] = l_cell_wire[193];							inform_L[193][4] = l_cell_wire[194];							inform_L[209][4] = l_cell_wire[195];							inform_L[194][4] = l_cell_wire[196];							inform_L[210][4] = l_cell_wire[197];							inform_L[195][4] = l_cell_wire[198];							inform_L[211][4] = l_cell_wire[199];							inform_L[196][4] = l_cell_wire[200];							inform_L[212][4] = l_cell_wire[201];							inform_L[197][4] = l_cell_wire[202];							inform_L[213][4] = l_cell_wire[203];							inform_L[198][4] = l_cell_wire[204];							inform_L[214][4] = l_cell_wire[205];							inform_L[199][4] = l_cell_wire[206];							inform_L[215][4] = l_cell_wire[207];							inform_L[200][4] = l_cell_wire[208];							inform_L[216][4] = l_cell_wire[209];							inform_L[201][4] = l_cell_wire[210];							inform_L[217][4] = l_cell_wire[211];							inform_L[202][4] = l_cell_wire[212];							inform_L[218][4] = l_cell_wire[213];							inform_L[203][4] = l_cell_wire[214];							inform_L[219][4] = l_cell_wire[215];							inform_L[204][4] = l_cell_wire[216];							inform_L[220][4] = l_cell_wire[217];							inform_L[205][4] = l_cell_wire[218];							inform_L[221][4] = l_cell_wire[219];							inform_L[206][4] = l_cell_wire[220];							inform_L[222][4] = l_cell_wire[221];							inform_L[207][4] = l_cell_wire[222];							inform_L[223][4] = l_cell_wire[223];							inform_L[224][4] = l_cell_wire[224];							inform_L[240][4] = l_cell_wire[225];							inform_L[225][4] = l_cell_wire[226];							inform_L[241][4] = l_cell_wire[227];							inform_L[226][4] = l_cell_wire[228];							inform_L[242][4] = l_cell_wire[229];							inform_L[227][4] = l_cell_wire[230];							inform_L[243][4] = l_cell_wire[231];							inform_L[228][4] = l_cell_wire[232];							inform_L[244][4] = l_cell_wire[233];							inform_L[229][4] = l_cell_wire[234];							inform_L[245][4] = l_cell_wire[235];							inform_L[230][4] = l_cell_wire[236];							inform_L[246][4] = l_cell_wire[237];							inform_L[231][4] = l_cell_wire[238];							inform_L[247][4] = l_cell_wire[239];							inform_L[232][4] = l_cell_wire[240];							inform_L[248][4] = l_cell_wire[241];							inform_L[233][4] = l_cell_wire[242];							inform_L[249][4] = l_cell_wire[243];							inform_L[234][4] = l_cell_wire[244];							inform_L[250][4] = l_cell_wire[245];							inform_L[235][4] = l_cell_wire[246];							inform_L[251][4] = l_cell_wire[247];							inform_L[236][4] = l_cell_wire[248];							inform_L[252][4] = l_cell_wire[249];							inform_L[237][4] = l_cell_wire[250];							inform_L[253][4] = l_cell_wire[251];							inform_L[238][4] = l_cell_wire[252];							inform_L[254][4] = l_cell_wire[253];							inform_L[239][4] = l_cell_wire[254];							inform_L[255][4] = l_cell_wire[255];						end
						6:						begin							inform_R[0][6] = r_cell_wire[0];							inform_R[32][6] = r_cell_wire[1];							inform_R[1][6] = r_cell_wire[2];							inform_R[33][6] = r_cell_wire[3];							inform_R[2][6] = r_cell_wire[4];							inform_R[34][6] = r_cell_wire[5];							inform_R[3][6] = r_cell_wire[6];							inform_R[35][6] = r_cell_wire[7];							inform_R[4][6] = r_cell_wire[8];							inform_R[36][6] = r_cell_wire[9];							inform_R[5][6] = r_cell_wire[10];							inform_R[37][6] = r_cell_wire[11];							inform_R[6][6] = r_cell_wire[12];							inform_R[38][6] = r_cell_wire[13];							inform_R[7][6] = r_cell_wire[14];							inform_R[39][6] = r_cell_wire[15];							inform_R[8][6] = r_cell_wire[16];							inform_R[40][6] = r_cell_wire[17];							inform_R[9][6] = r_cell_wire[18];							inform_R[41][6] = r_cell_wire[19];							inform_R[10][6] = r_cell_wire[20];							inform_R[42][6] = r_cell_wire[21];							inform_R[11][6] = r_cell_wire[22];							inform_R[43][6] = r_cell_wire[23];							inform_R[12][6] = r_cell_wire[24];							inform_R[44][6] = r_cell_wire[25];							inform_R[13][6] = r_cell_wire[26];							inform_R[45][6] = r_cell_wire[27];							inform_R[14][6] = r_cell_wire[28];							inform_R[46][6] = r_cell_wire[29];							inform_R[15][6] = r_cell_wire[30];							inform_R[47][6] = r_cell_wire[31];							inform_R[16][6] = r_cell_wire[32];							inform_R[48][6] = r_cell_wire[33];							inform_R[17][6] = r_cell_wire[34];							inform_R[49][6] = r_cell_wire[35];							inform_R[18][6] = r_cell_wire[36];							inform_R[50][6] = r_cell_wire[37];							inform_R[19][6] = r_cell_wire[38];							inform_R[51][6] = r_cell_wire[39];							inform_R[20][6] = r_cell_wire[40];							inform_R[52][6] = r_cell_wire[41];							inform_R[21][6] = r_cell_wire[42];							inform_R[53][6] = r_cell_wire[43];							inform_R[22][6] = r_cell_wire[44];							inform_R[54][6] = r_cell_wire[45];							inform_R[23][6] = r_cell_wire[46];							inform_R[55][6] = r_cell_wire[47];							inform_R[24][6] = r_cell_wire[48];							inform_R[56][6] = r_cell_wire[49];							inform_R[25][6] = r_cell_wire[50];							inform_R[57][6] = r_cell_wire[51];							inform_R[26][6] = r_cell_wire[52];							inform_R[58][6] = r_cell_wire[53];							inform_R[27][6] = r_cell_wire[54];							inform_R[59][6] = r_cell_wire[55];							inform_R[28][6] = r_cell_wire[56];							inform_R[60][6] = r_cell_wire[57];							inform_R[29][6] = r_cell_wire[58];							inform_R[61][6] = r_cell_wire[59];							inform_R[30][6] = r_cell_wire[60];							inform_R[62][6] = r_cell_wire[61];							inform_R[31][6] = r_cell_wire[62];							inform_R[63][6] = r_cell_wire[63];							inform_R[64][6] = r_cell_wire[64];							inform_R[96][6] = r_cell_wire[65];							inform_R[65][6] = r_cell_wire[66];							inform_R[97][6] = r_cell_wire[67];							inform_R[66][6] = r_cell_wire[68];							inform_R[98][6] = r_cell_wire[69];							inform_R[67][6] = r_cell_wire[70];							inform_R[99][6] = r_cell_wire[71];							inform_R[68][6] = r_cell_wire[72];							inform_R[100][6] = r_cell_wire[73];							inform_R[69][6] = r_cell_wire[74];							inform_R[101][6] = r_cell_wire[75];							inform_R[70][6] = r_cell_wire[76];							inform_R[102][6] = r_cell_wire[77];							inform_R[71][6] = r_cell_wire[78];							inform_R[103][6] = r_cell_wire[79];							inform_R[72][6] = r_cell_wire[80];							inform_R[104][6] = r_cell_wire[81];							inform_R[73][6] = r_cell_wire[82];							inform_R[105][6] = r_cell_wire[83];							inform_R[74][6] = r_cell_wire[84];							inform_R[106][6] = r_cell_wire[85];							inform_R[75][6] = r_cell_wire[86];							inform_R[107][6] = r_cell_wire[87];							inform_R[76][6] = r_cell_wire[88];							inform_R[108][6] = r_cell_wire[89];							inform_R[77][6] = r_cell_wire[90];							inform_R[109][6] = r_cell_wire[91];							inform_R[78][6] = r_cell_wire[92];							inform_R[110][6] = r_cell_wire[93];							inform_R[79][6] = r_cell_wire[94];							inform_R[111][6] = r_cell_wire[95];							inform_R[80][6] = r_cell_wire[96];							inform_R[112][6] = r_cell_wire[97];							inform_R[81][6] = r_cell_wire[98];							inform_R[113][6] = r_cell_wire[99];							inform_R[82][6] = r_cell_wire[100];							inform_R[114][6] = r_cell_wire[101];							inform_R[83][6] = r_cell_wire[102];							inform_R[115][6] = r_cell_wire[103];							inform_R[84][6] = r_cell_wire[104];							inform_R[116][6] = r_cell_wire[105];							inform_R[85][6] = r_cell_wire[106];							inform_R[117][6] = r_cell_wire[107];							inform_R[86][6] = r_cell_wire[108];							inform_R[118][6] = r_cell_wire[109];							inform_R[87][6] = r_cell_wire[110];							inform_R[119][6] = r_cell_wire[111];							inform_R[88][6] = r_cell_wire[112];							inform_R[120][6] = r_cell_wire[113];							inform_R[89][6] = r_cell_wire[114];							inform_R[121][6] = r_cell_wire[115];							inform_R[90][6] = r_cell_wire[116];							inform_R[122][6] = r_cell_wire[117];							inform_R[91][6] = r_cell_wire[118];							inform_R[123][6] = r_cell_wire[119];							inform_R[92][6] = r_cell_wire[120];							inform_R[124][6] = r_cell_wire[121];							inform_R[93][6] = r_cell_wire[122];							inform_R[125][6] = r_cell_wire[123];							inform_R[94][6] = r_cell_wire[124];							inform_R[126][6] = r_cell_wire[125];							inform_R[95][6] = r_cell_wire[126];							inform_R[127][6] = r_cell_wire[127];							inform_R[128][6] = r_cell_wire[128];							inform_R[160][6] = r_cell_wire[129];							inform_R[129][6] = r_cell_wire[130];							inform_R[161][6] = r_cell_wire[131];							inform_R[130][6] = r_cell_wire[132];							inform_R[162][6] = r_cell_wire[133];							inform_R[131][6] = r_cell_wire[134];							inform_R[163][6] = r_cell_wire[135];							inform_R[132][6] = r_cell_wire[136];							inform_R[164][6] = r_cell_wire[137];							inform_R[133][6] = r_cell_wire[138];							inform_R[165][6] = r_cell_wire[139];							inform_R[134][6] = r_cell_wire[140];							inform_R[166][6] = r_cell_wire[141];							inform_R[135][6] = r_cell_wire[142];							inform_R[167][6] = r_cell_wire[143];							inform_R[136][6] = r_cell_wire[144];							inform_R[168][6] = r_cell_wire[145];							inform_R[137][6] = r_cell_wire[146];							inform_R[169][6] = r_cell_wire[147];							inform_R[138][6] = r_cell_wire[148];							inform_R[170][6] = r_cell_wire[149];							inform_R[139][6] = r_cell_wire[150];							inform_R[171][6] = r_cell_wire[151];							inform_R[140][6] = r_cell_wire[152];							inform_R[172][6] = r_cell_wire[153];							inform_R[141][6] = r_cell_wire[154];							inform_R[173][6] = r_cell_wire[155];							inform_R[142][6] = r_cell_wire[156];							inform_R[174][6] = r_cell_wire[157];							inform_R[143][6] = r_cell_wire[158];							inform_R[175][6] = r_cell_wire[159];							inform_R[144][6] = r_cell_wire[160];							inform_R[176][6] = r_cell_wire[161];							inform_R[145][6] = r_cell_wire[162];							inform_R[177][6] = r_cell_wire[163];							inform_R[146][6] = r_cell_wire[164];							inform_R[178][6] = r_cell_wire[165];							inform_R[147][6] = r_cell_wire[166];							inform_R[179][6] = r_cell_wire[167];							inform_R[148][6] = r_cell_wire[168];							inform_R[180][6] = r_cell_wire[169];							inform_R[149][6] = r_cell_wire[170];							inform_R[181][6] = r_cell_wire[171];							inform_R[150][6] = r_cell_wire[172];							inform_R[182][6] = r_cell_wire[173];							inform_R[151][6] = r_cell_wire[174];							inform_R[183][6] = r_cell_wire[175];							inform_R[152][6] = r_cell_wire[176];							inform_R[184][6] = r_cell_wire[177];							inform_R[153][6] = r_cell_wire[178];							inform_R[185][6] = r_cell_wire[179];							inform_R[154][6] = r_cell_wire[180];							inform_R[186][6] = r_cell_wire[181];							inform_R[155][6] = r_cell_wire[182];							inform_R[187][6] = r_cell_wire[183];							inform_R[156][6] = r_cell_wire[184];							inform_R[188][6] = r_cell_wire[185];							inform_R[157][6] = r_cell_wire[186];							inform_R[189][6] = r_cell_wire[187];							inform_R[158][6] = r_cell_wire[188];							inform_R[190][6] = r_cell_wire[189];							inform_R[159][6] = r_cell_wire[190];							inform_R[191][6] = r_cell_wire[191];							inform_R[192][6] = r_cell_wire[192];							inform_R[224][6] = r_cell_wire[193];							inform_R[193][6] = r_cell_wire[194];							inform_R[225][6] = r_cell_wire[195];							inform_R[194][6] = r_cell_wire[196];							inform_R[226][6] = r_cell_wire[197];							inform_R[195][6] = r_cell_wire[198];							inform_R[227][6] = r_cell_wire[199];							inform_R[196][6] = r_cell_wire[200];							inform_R[228][6] = r_cell_wire[201];							inform_R[197][6] = r_cell_wire[202];							inform_R[229][6] = r_cell_wire[203];							inform_R[198][6] = r_cell_wire[204];							inform_R[230][6] = r_cell_wire[205];							inform_R[199][6] = r_cell_wire[206];							inform_R[231][6] = r_cell_wire[207];							inform_R[200][6] = r_cell_wire[208];							inform_R[232][6] = r_cell_wire[209];							inform_R[201][6] = r_cell_wire[210];							inform_R[233][6] = r_cell_wire[211];							inform_R[202][6] = r_cell_wire[212];							inform_R[234][6] = r_cell_wire[213];							inform_R[203][6] = r_cell_wire[214];							inform_R[235][6] = r_cell_wire[215];							inform_R[204][6] = r_cell_wire[216];							inform_R[236][6] = r_cell_wire[217];							inform_R[205][6] = r_cell_wire[218];							inform_R[237][6] = r_cell_wire[219];							inform_R[206][6] = r_cell_wire[220];							inform_R[238][6] = r_cell_wire[221];							inform_R[207][6] = r_cell_wire[222];							inform_R[239][6] = r_cell_wire[223];							inform_R[208][6] = r_cell_wire[224];							inform_R[240][6] = r_cell_wire[225];							inform_R[209][6] = r_cell_wire[226];							inform_R[241][6] = r_cell_wire[227];							inform_R[210][6] = r_cell_wire[228];							inform_R[242][6] = r_cell_wire[229];							inform_R[211][6] = r_cell_wire[230];							inform_R[243][6] = r_cell_wire[231];							inform_R[212][6] = r_cell_wire[232];							inform_R[244][6] = r_cell_wire[233];							inform_R[213][6] = r_cell_wire[234];							inform_R[245][6] = r_cell_wire[235];							inform_R[214][6] = r_cell_wire[236];							inform_R[246][6] = r_cell_wire[237];							inform_R[215][6] = r_cell_wire[238];							inform_R[247][6] = r_cell_wire[239];							inform_R[216][6] = r_cell_wire[240];							inform_R[248][6] = r_cell_wire[241];							inform_R[217][6] = r_cell_wire[242];							inform_R[249][6] = r_cell_wire[243];							inform_R[218][6] = r_cell_wire[244];							inform_R[250][6] = r_cell_wire[245];							inform_R[219][6] = r_cell_wire[246];							inform_R[251][6] = r_cell_wire[247];							inform_R[220][6] = r_cell_wire[248];							inform_R[252][6] = r_cell_wire[249];							inform_R[221][6] = r_cell_wire[250];							inform_R[253][6] = r_cell_wire[251];							inform_R[222][6] = r_cell_wire[252];							inform_R[254][6] = r_cell_wire[253];							inform_R[223][6] = r_cell_wire[254];							inform_R[255][6] = r_cell_wire[255];							inform_L[0][5] = l_cell_wire[0];							inform_L[32][5] = l_cell_wire[1];							inform_L[1][5] = l_cell_wire[2];							inform_L[33][5] = l_cell_wire[3];							inform_L[2][5] = l_cell_wire[4];							inform_L[34][5] = l_cell_wire[5];							inform_L[3][5] = l_cell_wire[6];							inform_L[35][5] = l_cell_wire[7];							inform_L[4][5] = l_cell_wire[8];							inform_L[36][5] = l_cell_wire[9];							inform_L[5][5] = l_cell_wire[10];							inform_L[37][5] = l_cell_wire[11];							inform_L[6][5] = l_cell_wire[12];							inform_L[38][5] = l_cell_wire[13];							inform_L[7][5] = l_cell_wire[14];							inform_L[39][5] = l_cell_wire[15];							inform_L[8][5] = l_cell_wire[16];							inform_L[40][5] = l_cell_wire[17];							inform_L[9][5] = l_cell_wire[18];							inform_L[41][5] = l_cell_wire[19];							inform_L[10][5] = l_cell_wire[20];							inform_L[42][5] = l_cell_wire[21];							inform_L[11][5] = l_cell_wire[22];							inform_L[43][5] = l_cell_wire[23];							inform_L[12][5] = l_cell_wire[24];							inform_L[44][5] = l_cell_wire[25];							inform_L[13][5] = l_cell_wire[26];							inform_L[45][5] = l_cell_wire[27];							inform_L[14][5] = l_cell_wire[28];							inform_L[46][5] = l_cell_wire[29];							inform_L[15][5] = l_cell_wire[30];							inform_L[47][5] = l_cell_wire[31];							inform_L[16][5] = l_cell_wire[32];							inform_L[48][5] = l_cell_wire[33];							inform_L[17][5] = l_cell_wire[34];							inform_L[49][5] = l_cell_wire[35];							inform_L[18][5] = l_cell_wire[36];							inform_L[50][5] = l_cell_wire[37];							inform_L[19][5] = l_cell_wire[38];							inform_L[51][5] = l_cell_wire[39];							inform_L[20][5] = l_cell_wire[40];							inform_L[52][5] = l_cell_wire[41];							inform_L[21][5] = l_cell_wire[42];							inform_L[53][5] = l_cell_wire[43];							inform_L[22][5] = l_cell_wire[44];							inform_L[54][5] = l_cell_wire[45];							inform_L[23][5] = l_cell_wire[46];							inform_L[55][5] = l_cell_wire[47];							inform_L[24][5] = l_cell_wire[48];							inform_L[56][5] = l_cell_wire[49];							inform_L[25][5] = l_cell_wire[50];							inform_L[57][5] = l_cell_wire[51];							inform_L[26][5] = l_cell_wire[52];							inform_L[58][5] = l_cell_wire[53];							inform_L[27][5] = l_cell_wire[54];							inform_L[59][5] = l_cell_wire[55];							inform_L[28][5] = l_cell_wire[56];							inform_L[60][5] = l_cell_wire[57];							inform_L[29][5] = l_cell_wire[58];							inform_L[61][5] = l_cell_wire[59];							inform_L[30][5] = l_cell_wire[60];							inform_L[62][5] = l_cell_wire[61];							inform_L[31][5] = l_cell_wire[62];							inform_L[63][5] = l_cell_wire[63];							inform_L[64][5] = l_cell_wire[64];							inform_L[96][5] = l_cell_wire[65];							inform_L[65][5] = l_cell_wire[66];							inform_L[97][5] = l_cell_wire[67];							inform_L[66][5] = l_cell_wire[68];							inform_L[98][5] = l_cell_wire[69];							inform_L[67][5] = l_cell_wire[70];							inform_L[99][5] = l_cell_wire[71];							inform_L[68][5] = l_cell_wire[72];							inform_L[100][5] = l_cell_wire[73];							inform_L[69][5] = l_cell_wire[74];							inform_L[101][5] = l_cell_wire[75];							inform_L[70][5] = l_cell_wire[76];							inform_L[102][5] = l_cell_wire[77];							inform_L[71][5] = l_cell_wire[78];							inform_L[103][5] = l_cell_wire[79];							inform_L[72][5] = l_cell_wire[80];							inform_L[104][5] = l_cell_wire[81];							inform_L[73][5] = l_cell_wire[82];							inform_L[105][5] = l_cell_wire[83];							inform_L[74][5] = l_cell_wire[84];							inform_L[106][5] = l_cell_wire[85];							inform_L[75][5] = l_cell_wire[86];							inform_L[107][5] = l_cell_wire[87];							inform_L[76][5] = l_cell_wire[88];							inform_L[108][5] = l_cell_wire[89];							inform_L[77][5] = l_cell_wire[90];							inform_L[109][5] = l_cell_wire[91];							inform_L[78][5] = l_cell_wire[92];							inform_L[110][5] = l_cell_wire[93];							inform_L[79][5] = l_cell_wire[94];							inform_L[111][5] = l_cell_wire[95];							inform_L[80][5] = l_cell_wire[96];							inform_L[112][5] = l_cell_wire[97];							inform_L[81][5] = l_cell_wire[98];							inform_L[113][5] = l_cell_wire[99];							inform_L[82][5] = l_cell_wire[100];							inform_L[114][5] = l_cell_wire[101];							inform_L[83][5] = l_cell_wire[102];							inform_L[115][5] = l_cell_wire[103];							inform_L[84][5] = l_cell_wire[104];							inform_L[116][5] = l_cell_wire[105];							inform_L[85][5] = l_cell_wire[106];							inform_L[117][5] = l_cell_wire[107];							inform_L[86][5] = l_cell_wire[108];							inform_L[118][5] = l_cell_wire[109];							inform_L[87][5] = l_cell_wire[110];							inform_L[119][5] = l_cell_wire[111];							inform_L[88][5] = l_cell_wire[112];							inform_L[120][5] = l_cell_wire[113];							inform_L[89][5] = l_cell_wire[114];							inform_L[121][5] = l_cell_wire[115];							inform_L[90][5] = l_cell_wire[116];							inform_L[122][5] = l_cell_wire[117];							inform_L[91][5] = l_cell_wire[118];							inform_L[123][5] = l_cell_wire[119];							inform_L[92][5] = l_cell_wire[120];							inform_L[124][5] = l_cell_wire[121];							inform_L[93][5] = l_cell_wire[122];							inform_L[125][5] = l_cell_wire[123];							inform_L[94][5] = l_cell_wire[124];							inform_L[126][5] = l_cell_wire[125];							inform_L[95][5] = l_cell_wire[126];							inform_L[127][5] = l_cell_wire[127];							inform_L[128][5] = l_cell_wire[128];							inform_L[160][5] = l_cell_wire[129];							inform_L[129][5] = l_cell_wire[130];							inform_L[161][5] = l_cell_wire[131];							inform_L[130][5] = l_cell_wire[132];							inform_L[162][5] = l_cell_wire[133];							inform_L[131][5] = l_cell_wire[134];							inform_L[163][5] = l_cell_wire[135];							inform_L[132][5] = l_cell_wire[136];							inform_L[164][5] = l_cell_wire[137];							inform_L[133][5] = l_cell_wire[138];							inform_L[165][5] = l_cell_wire[139];							inform_L[134][5] = l_cell_wire[140];							inform_L[166][5] = l_cell_wire[141];							inform_L[135][5] = l_cell_wire[142];							inform_L[167][5] = l_cell_wire[143];							inform_L[136][5] = l_cell_wire[144];							inform_L[168][5] = l_cell_wire[145];							inform_L[137][5] = l_cell_wire[146];							inform_L[169][5] = l_cell_wire[147];							inform_L[138][5] = l_cell_wire[148];							inform_L[170][5] = l_cell_wire[149];							inform_L[139][5] = l_cell_wire[150];							inform_L[171][5] = l_cell_wire[151];							inform_L[140][5] = l_cell_wire[152];							inform_L[172][5] = l_cell_wire[153];							inform_L[141][5] = l_cell_wire[154];							inform_L[173][5] = l_cell_wire[155];							inform_L[142][5] = l_cell_wire[156];							inform_L[174][5] = l_cell_wire[157];							inform_L[143][5] = l_cell_wire[158];							inform_L[175][5] = l_cell_wire[159];							inform_L[144][5] = l_cell_wire[160];							inform_L[176][5] = l_cell_wire[161];							inform_L[145][5] = l_cell_wire[162];							inform_L[177][5] = l_cell_wire[163];							inform_L[146][5] = l_cell_wire[164];							inform_L[178][5] = l_cell_wire[165];							inform_L[147][5] = l_cell_wire[166];							inform_L[179][5] = l_cell_wire[167];							inform_L[148][5] = l_cell_wire[168];							inform_L[180][5] = l_cell_wire[169];							inform_L[149][5] = l_cell_wire[170];							inform_L[181][5] = l_cell_wire[171];							inform_L[150][5] = l_cell_wire[172];							inform_L[182][5] = l_cell_wire[173];							inform_L[151][5] = l_cell_wire[174];							inform_L[183][5] = l_cell_wire[175];							inform_L[152][5] = l_cell_wire[176];							inform_L[184][5] = l_cell_wire[177];							inform_L[153][5] = l_cell_wire[178];							inform_L[185][5] = l_cell_wire[179];							inform_L[154][5] = l_cell_wire[180];							inform_L[186][5] = l_cell_wire[181];							inform_L[155][5] = l_cell_wire[182];							inform_L[187][5] = l_cell_wire[183];							inform_L[156][5] = l_cell_wire[184];							inform_L[188][5] = l_cell_wire[185];							inform_L[157][5] = l_cell_wire[186];							inform_L[189][5] = l_cell_wire[187];							inform_L[158][5] = l_cell_wire[188];							inform_L[190][5] = l_cell_wire[189];							inform_L[159][5] = l_cell_wire[190];							inform_L[191][5] = l_cell_wire[191];							inform_L[192][5] = l_cell_wire[192];							inform_L[224][5] = l_cell_wire[193];							inform_L[193][5] = l_cell_wire[194];							inform_L[225][5] = l_cell_wire[195];							inform_L[194][5] = l_cell_wire[196];							inform_L[226][5] = l_cell_wire[197];							inform_L[195][5] = l_cell_wire[198];							inform_L[227][5] = l_cell_wire[199];							inform_L[196][5] = l_cell_wire[200];							inform_L[228][5] = l_cell_wire[201];							inform_L[197][5] = l_cell_wire[202];							inform_L[229][5] = l_cell_wire[203];							inform_L[198][5] = l_cell_wire[204];							inform_L[230][5] = l_cell_wire[205];							inform_L[199][5] = l_cell_wire[206];							inform_L[231][5] = l_cell_wire[207];							inform_L[200][5] = l_cell_wire[208];							inform_L[232][5] = l_cell_wire[209];							inform_L[201][5] = l_cell_wire[210];							inform_L[233][5] = l_cell_wire[211];							inform_L[202][5] = l_cell_wire[212];							inform_L[234][5] = l_cell_wire[213];							inform_L[203][5] = l_cell_wire[214];							inform_L[235][5] = l_cell_wire[215];							inform_L[204][5] = l_cell_wire[216];							inform_L[236][5] = l_cell_wire[217];							inform_L[205][5] = l_cell_wire[218];							inform_L[237][5] = l_cell_wire[219];							inform_L[206][5] = l_cell_wire[220];							inform_L[238][5] = l_cell_wire[221];							inform_L[207][5] = l_cell_wire[222];							inform_L[239][5] = l_cell_wire[223];							inform_L[208][5] = l_cell_wire[224];							inform_L[240][5] = l_cell_wire[225];							inform_L[209][5] = l_cell_wire[226];							inform_L[241][5] = l_cell_wire[227];							inform_L[210][5] = l_cell_wire[228];							inform_L[242][5] = l_cell_wire[229];							inform_L[211][5] = l_cell_wire[230];							inform_L[243][5] = l_cell_wire[231];							inform_L[212][5] = l_cell_wire[232];							inform_L[244][5] = l_cell_wire[233];							inform_L[213][5] = l_cell_wire[234];							inform_L[245][5] = l_cell_wire[235];							inform_L[214][5] = l_cell_wire[236];							inform_L[246][5] = l_cell_wire[237];							inform_L[215][5] = l_cell_wire[238];							inform_L[247][5] = l_cell_wire[239];							inform_L[216][5] = l_cell_wire[240];							inform_L[248][5] = l_cell_wire[241];							inform_L[217][5] = l_cell_wire[242];							inform_L[249][5] = l_cell_wire[243];							inform_L[218][5] = l_cell_wire[244];							inform_L[250][5] = l_cell_wire[245];							inform_L[219][5] = l_cell_wire[246];							inform_L[251][5] = l_cell_wire[247];							inform_L[220][5] = l_cell_wire[248];							inform_L[252][5] = l_cell_wire[249];							inform_L[221][5] = l_cell_wire[250];							inform_L[253][5] = l_cell_wire[251];							inform_L[222][5] = l_cell_wire[252];							inform_L[254][5] = l_cell_wire[253];							inform_L[223][5] = l_cell_wire[254];							inform_L[255][5] = l_cell_wire[255];						end
						7:						begin							inform_R[0][7] = r_cell_wire[0];							inform_R[64][7] = r_cell_wire[1];							inform_R[1][7] = r_cell_wire[2];							inform_R[65][7] = r_cell_wire[3];							inform_R[2][7] = r_cell_wire[4];							inform_R[66][7] = r_cell_wire[5];							inform_R[3][7] = r_cell_wire[6];							inform_R[67][7] = r_cell_wire[7];							inform_R[4][7] = r_cell_wire[8];							inform_R[68][7] = r_cell_wire[9];							inform_R[5][7] = r_cell_wire[10];							inform_R[69][7] = r_cell_wire[11];							inform_R[6][7] = r_cell_wire[12];							inform_R[70][7] = r_cell_wire[13];							inform_R[7][7] = r_cell_wire[14];							inform_R[71][7] = r_cell_wire[15];							inform_R[8][7] = r_cell_wire[16];							inform_R[72][7] = r_cell_wire[17];							inform_R[9][7] = r_cell_wire[18];							inform_R[73][7] = r_cell_wire[19];							inform_R[10][7] = r_cell_wire[20];							inform_R[74][7] = r_cell_wire[21];							inform_R[11][7] = r_cell_wire[22];							inform_R[75][7] = r_cell_wire[23];							inform_R[12][7] = r_cell_wire[24];							inform_R[76][7] = r_cell_wire[25];							inform_R[13][7] = r_cell_wire[26];							inform_R[77][7] = r_cell_wire[27];							inform_R[14][7] = r_cell_wire[28];							inform_R[78][7] = r_cell_wire[29];							inform_R[15][7] = r_cell_wire[30];							inform_R[79][7] = r_cell_wire[31];							inform_R[16][7] = r_cell_wire[32];							inform_R[80][7] = r_cell_wire[33];							inform_R[17][7] = r_cell_wire[34];							inform_R[81][7] = r_cell_wire[35];							inform_R[18][7] = r_cell_wire[36];							inform_R[82][7] = r_cell_wire[37];							inform_R[19][7] = r_cell_wire[38];							inform_R[83][7] = r_cell_wire[39];							inform_R[20][7] = r_cell_wire[40];							inform_R[84][7] = r_cell_wire[41];							inform_R[21][7] = r_cell_wire[42];							inform_R[85][7] = r_cell_wire[43];							inform_R[22][7] = r_cell_wire[44];							inform_R[86][7] = r_cell_wire[45];							inform_R[23][7] = r_cell_wire[46];							inform_R[87][7] = r_cell_wire[47];							inform_R[24][7] = r_cell_wire[48];							inform_R[88][7] = r_cell_wire[49];							inform_R[25][7] = r_cell_wire[50];							inform_R[89][7] = r_cell_wire[51];							inform_R[26][7] = r_cell_wire[52];							inform_R[90][7] = r_cell_wire[53];							inform_R[27][7] = r_cell_wire[54];							inform_R[91][7] = r_cell_wire[55];							inform_R[28][7] = r_cell_wire[56];							inform_R[92][7] = r_cell_wire[57];							inform_R[29][7] = r_cell_wire[58];							inform_R[93][7] = r_cell_wire[59];							inform_R[30][7] = r_cell_wire[60];							inform_R[94][7] = r_cell_wire[61];							inform_R[31][7] = r_cell_wire[62];							inform_R[95][7] = r_cell_wire[63];							inform_R[32][7] = r_cell_wire[64];							inform_R[96][7] = r_cell_wire[65];							inform_R[33][7] = r_cell_wire[66];							inform_R[97][7] = r_cell_wire[67];							inform_R[34][7] = r_cell_wire[68];							inform_R[98][7] = r_cell_wire[69];							inform_R[35][7] = r_cell_wire[70];							inform_R[99][7] = r_cell_wire[71];							inform_R[36][7] = r_cell_wire[72];							inform_R[100][7] = r_cell_wire[73];							inform_R[37][7] = r_cell_wire[74];							inform_R[101][7] = r_cell_wire[75];							inform_R[38][7] = r_cell_wire[76];							inform_R[102][7] = r_cell_wire[77];							inform_R[39][7] = r_cell_wire[78];							inform_R[103][7] = r_cell_wire[79];							inform_R[40][7] = r_cell_wire[80];							inform_R[104][7] = r_cell_wire[81];							inform_R[41][7] = r_cell_wire[82];							inform_R[105][7] = r_cell_wire[83];							inform_R[42][7] = r_cell_wire[84];							inform_R[106][7] = r_cell_wire[85];							inform_R[43][7] = r_cell_wire[86];							inform_R[107][7] = r_cell_wire[87];							inform_R[44][7] = r_cell_wire[88];							inform_R[108][7] = r_cell_wire[89];							inform_R[45][7] = r_cell_wire[90];							inform_R[109][7] = r_cell_wire[91];							inform_R[46][7] = r_cell_wire[92];							inform_R[110][7] = r_cell_wire[93];							inform_R[47][7] = r_cell_wire[94];							inform_R[111][7] = r_cell_wire[95];							inform_R[48][7] = r_cell_wire[96];							inform_R[112][7] = r_cell_wire[97];							inform_R[49][7] = r_cell_wire[98];							inform_R[113][7] = r_cell_wire[99];							inform_R[50][7] = r_cell_wire[100];							inform_R[114][7] = r_cell_wire[101];							inform_R[51][7] = r_cell_wire[102];							inform_R[115][7] = r_cell_wire[103];							inform_R[52][7] = r_cell_wire[104];							inform_R[116][7] = r_cell_wire[105];							inform_R[53][7] = r_cell_wire[106];							inform_R[117][7] = r_cell_wire[107];							inform_R[54][7] = r_cell_wire[108];							inform_R[118][7] = r_cell_wire[109];							inform_R[55][7] = r_cell_wire[110];							inform_R[119][7] = r_cell_wire[111];							inform_R[56][7] = r_cell_wire[112];							inform_R[120][7] = r_cell_wire[113];							inform_R[57][7] = r_cell_wire[114];							inform_R[121][7] = r_cell_wire[115];							inform_R[58][7] = r_cell_wire[116];							inform_R[122][7] = r_cell_wire[117];							inform_R[59][7] = r_cell_wire[118];							inform_R[123][7] = r_cell_wire[119];							inform_R[60][7] = r_cell_wire[120];							inform_R[124][7] = r_cell_wire[121];							inform_R[61][7] = r_cell_wire[122];							inform_R[125][7] = r_cell_wire[123];							inform_R[62][7] = r_cell_wire[124];							inform_R[126][7] = r_cell_wire[125];							inform_R[63][7] = r_cell_wire[126];							inform_R[127][7] = r_cell_wire[127];							inform_R[128][7] = r_cell_wire[128];							inform_R[192][7] = r_cell_wire[129];							inform_R[129][7] = r_cell_wire[130];							inform_R[193][7] = r_cell_wire[131];							inform_R[130][7] = r_cell_wire[132];							inform_R[194][7] = r_cell_wire[133];							inform_R[131][7] = r_cell_wire[134];							inform_R[195][7] = r_cell_wire[135];							inform_R[132][7] = r_cell_wire[136];							inform_R[196][7] = r_cell_wire[137];							inform_R[133][7] = r_cell_wire[138];							inform_R[197][7] = r_cell_wire[139];							inform_R[134][7] = r_cell_wire[140];							inform_R[198][7] = r_cell_wire[141];							inform_R[135][7] = r_cell_wire[142];							inform_R[199][7] = r_cell_wire[143];							inform_R[136][7] = r_cell_wire[144];							inform_R[200][7] = r_cell_wire[145];							inform_R[137][7] = r_cell_wire[146];							inform_R[201][7] = r_cell_wire[147];							inform_R[138][7] = r_cell_wire[148];							inform_R[202][7] = r_cell_wire[149];							inform_R[139][7] = r_cell_wire[150];							inform_R[203][7] = r_cell_wire[151];							inform_R[140][7] = r_cell_wire[152];							inform_R[204][7] = r_cell_wire[153];							inform_R[141][7] = r_cell_wire[154];							inform_R[205][7] = r_cell_wire[155];							inform_R[142][7] = r_cell_wire[156];							inform_R[206][7] = r_cell_wire[157];							inform_R[143][7] = r_cell_wire[158];							inform_R[207][7] = r_cell_wire[159];							inform_R[144][7] = r_cell_wire[160];							inform_R[208][7] = r_cell_wire[161];							inform_R[145][7] = r_cell_wire[162];							inform_R[209][7] = r_cell_wire[163];							inform_R[146][7] = r_cell_wire[164];							inform_R[210][7] = r_cell_wire[165];							inform_R[147][7] = r_cell_wire[166];							inform_R[211][7] = r_cell_wire[167];							inform_R[148][7] = r_cell_wire[168];							inform_R[212][7] = r_cell_wire[169];							inform_R[149][7] = r_cell_wire[170];							inform_R[213][7] = r_cell_wire[171];							inform_R[150][7] = r_cell_wire[172];							inform_R[214][7] = r_cell_wire[173];							inform_R[151][7] = r_cell_wire[174];							inform_R[215][7] = r_cell_wire[175];							inform_R[152][7] = r_cell_wire[176];							inform_R[216][7] = r_cell_wire[177];							inform_R[153][7] = r_cell_wire[178];							inform_R[217][7] = r_cell_wire[179];							inform_R[154][7] = r_cell_wire[180];							inform_R[218][7] = r_cell_wire[181];							inform_R[155][7] = r_cell_wire[182];							inform_R[219][7] = r_cell_wire[183];							inform_R[156][7] = r_cell_wire[184];							inform_R[220][7] = r_cell_wire[185];							inform_R[157][7] = r_cell_wire[186];							inform_R[221][7] = r_cell_wire[187];							inform_R[158][7] = r_cell_wire[188];							inform_R[222][7] = r_cell_wire[189];							inform_R[159][7] = r_cell_wire[190];							inform_R[223][7] = r_cell_wire[191];							inform_R[160][7] = r_cell_wire[192];							inform_R[224][7] = r_cell_wire[193];							inform_R[161][7] = r_cell_wire[194];							inform_R[225][7] = r_cell_wire[195];							inform_R[162][7] = r_cell_wire[196];							inform_R[226][7] = r_cell_wire[197];							inform_R[163][7] = r_cell_wire[198];							inform_R[227][7] = r_cell_wire[199];							inform_R[164][7] = r_cell_wire[200];							inform_R[228][7] = r_cell_wire[201];							inform_R[165][7] = r_cell_wire[202];							inform_R[229][7] = r_cell_wire[203];							inform_R[166][7] = r_cell_wire[204];							inform_R[230][7] = r_cell_wire[205];							inform_R[167][7] = r_cell_wire[206];							inform_R[231][7] = r_cell_wire[207];							inform_R[168][7] = r_cell_wire[208];							inform_R[232][7] = r_cell_wire[209];							inform_R[169][7] = r_cell_wire[210];							inform_R[233][7] = r_cell_wire[211];							inform_R[170][7] = r_cell_wire[212];							inform_R[234][7] = r_cell_wire[213];							inform_R[171][7] = r_cell_wire[214];							inform_R[235][7] = r_cell_wire[215];							inform_R[172][7] = r_cell_wire[216];							inform_R[236][7] = r_cell_wire[217];							inform_R[173][7] = r_cell_wire[218];							inform_R[237][7] = r_cell_wire[219];							inform_R[174][7] = r_cell_wire[220];							inform_R[238][7] = r_cell_wire[221];							inform_R[175][7] = r_cell_wire[222];							inform_R[239][7] = r_cell_wire[223];							inform_R[176][7] = r_cell_wire[224];							inform_R[240][7] = r_cell_wire[225];							inform_R[177][7] = r_cell_wire[226];							inform_R[241][7] = r_cell_wire[227];							inform_R[178][7] = r_cell_wire[228];							inform_R[242][7] = r_cell_wire[229];							inform_R[179][7] = r_cell_wire[230];							inform_R[243][7] = r_cell_wire[231];							inform_R[180][7] = r_cell_wire[232];							inform_R[244][7] = r_cell_wire[233];							inform_R[181][7] = r_cell_wire[234];							inform_R[245][7] = r_cell_wire[235];							inform_R[182][7] = r_cell_wire[236];							inform_R[246][7] = r_cell_wire[237];							inform_R[183][7] = r_cell_wire[238];							inform_R[247][7] = r_cell_wire[239];							inform_R[184][7] = r_cell_wire[240];							inform_R[248][7] = r_cell_wire[241];							inform_R[185][7] = r_cell_wire[242];							inform_R[249][7] = r_cell_wire[243];							inform_R[186][7] = r_cell_wire[244];							inform_R[250][7] = r_cell_wire[245];							inform_R[187][7] = r_cell_wire[246];							inform_R[251][7] = r_cell_wire[247];							inform_R[188][7] = r_cell_wire[248];							inform_R[252][7] = r_cell_wire[249];							inform_R[189][7] = r_cell_wire[250];							inform_R[253][7] = r_cell_wire[251];							inform_R[190][7] = r_cell_wire[252];							inform_R[254][7] = r_cell_wire[253];							inform_R[191][7] = r_cell_wire[254];							inform_R[255][7] = r_cell_wire[255];							inform_L[0][6] = l_cell_wire[0];							inform_L[64][6] = l_cell_wire[1];							inform_L[1][6] = l_cell_wire[2];							inform_L[65][6] = l_cell_wire[3];							inform_L[2][6] = l_cell_wire[4];							inform_L[66][6] = l_cell_wire[5];							inform_L[3][6] = l_cell_wire[6];							inform_L[67][6] = l_cell_wire[7];							inform_L[4][6] = l_cell_wire[8];							inform_L[68][6] = l_cell_wire[9];							inform_L[5][6] = l_cell_wire[10];							inform_L[69][6] = l_cell_wire[11];							inform_L[6][6] = l_cell_wire[12];							inform_L[70][6] = l_cell_wire[13];							inform_L[7][6] = l_cell_wire[14];							inform_L[71][6] = l_cell_wire[15];							inform_L[8][6] = l_cell_wire[16];							inform_L[72][6] = l_cell_wire[17];							inform_L[9][6] = l_cell_wire[18];							inform_L[73][6] = l_cell_wire[19];							inform_L[10][6] = l_cell_wire[20];							inform_L[74][6] = l_cell_wire[21];							inform_L[11][6] = l_cell_wire[22];							inform_L[75][6] = l_cell_wire[23];							inform_L[12][6] = l_cell_wire[24];							inform_L[76][6] = l_cell_wire[25];							inform_L[13][6] = l_cell_wire[26];							inform_L[77][6] = l_cell_wire[27];							inform_L[14][6] = l_cell_wire[28];							inform_L[78][6] = l_cell_wire[29];							inform_L[15][6] = l_cell_wire[30];							inform_L[79][6] = l_cell_wire[31];							inform_L[16][6] = l_cell_wire[32];							inform_L[80][6] = l_cell_wire[33];							inform_L[17][6] = l_cell_wire[34];							inform_L[81][6] = l_cell_wire[35];							inform_L[18][6] = l_cell_wire[36];							inform_L[82][6] = l_cell_wire[37];							inform_L[19][6] = l_cell_wire[38];							inform_L[83][6] = l_cell_wire[39];							inform_L[20][6] = l_cell_wire[40];							inform_L[84][6] = l_cell_wire[41];							inform_L[21][6] = l_cell_wire[42];							inform_L[85][6] = l_cell_wire[43];							inform_L[22][6] = l_cell_wire[44];							inform_L[86][6] = l_cell_wire[45];							inform_L[23][6] = l_cell_wire[46];							inform_L[87][6] = l_cell_wire[47];							inform_L[24][6] = l_cell_wire[48];							inform_L[88][6] = l_cell_wire[49];							inform_L[25][6] = l_cell_wire[50];							inform_L[89][6] = l_cell_wire[51];							inform_L[26][6] = l_cell_wire[52];							inform_L[90][6] = l_cell_wire[53];							inform_L[27][6] = l_cell_wire[54];							inform_L[91][6] = l_cell_wire[55];							inform_L[28][6] = l_cell_wire[56];							inform_L[92][6] = l_cell_wire[57];							inform_L[29][6] = l_cell_wire[58];							inform_L[93][6] = l_cell_wire[59];							inform_L[30][6] = l_cell_wire[60];							inform_L[94][6] = l_cell_wire[61];							inform_L[31][6] = l_cell_wire[62];							inform_L[95][6] = l_cell_wire[63];							inform_L[32][6] = l_cell_wire[64];							inform_L[96][6] = l_cell_wire[65];							inform_L[33][6] = l_cell_wire[66];							inform_L[97][6] = l_cell_wire[67];							inform_L[34][6] = l_cell_wire[68];							inform_L[98][6] = l_cell_wire[69];							inform_L[35][6] = l_cell_wire[70];							inform_L[99][6] = l_cell_wire[71];							inform_L[36][6] = l_cell_wire[72];							inform_L[100][6] = l_cell_wire[73];							inform_L[37][6] = l_cell_wire[74];							inform_L[101][6] = l_cell_wire[75];							inform_L[38][6] = l_cell_wire[76];							inform_L[102][6] = l_cell_wire[77];							inform_L[39][6] = l_cell_wire[78];							inform_L[103][6] = l_cell_wire[79];							inform_L[40][6] = l_cell_wire[80];							inform_L[104][6] = l_cell_wire[81];							inform_L[41][6] = l_cell_wire[82];							inform_L[105][6] = l_cell_wire[83];							inform_L[42][6] = l_cell_wire[84];							inform_L[106][6] = l_cell_wire[85];							inform_L[43][6] = l_cell_wire[86];							inform_L[107][6] = l_cell_wire[87];							inform_L[44][6] = l_cell_wire[88];							inform_L[108][6] = l_cell_wire[89];							inform_L[45][6] = l_cell_wire[90];							inform_L[109][6] = l_cell_wire[91];							inform_L[46][6] = l_cell_wire[92];							inform_L[110][6] = l_cell_wire[93];							inform_L[47][6] = l_cell_wire[94];							inform_L[111][6] = l_cell_wire[95];							inform_L[48][6] = l_cell_wire[96];							inform_L[112][6] = l_cell_wire[97];							inform_L[49][6] = l_cell_wire[98];							inform_L[113][6] = l_cell_wire[99];							inform_L[50][6] = l_cell_wire[100];							inform_L[114][6] = l_cell_wire[101];							inform_L[51][6] = l_cell_wire[102];							inform_L[115][6] = l_cell_wire[103];							inform_L[52][6] = l_cell_wire[104];							inform_L[116][6] = l_cell_wire[105];							inform_L[53][6] = l_cell_wire[106];							inform_L[117][6] = l_cell_wire[107];							inform_L[54][6] = l_cell_wire[108];							inform_L[118][6] = l_cell_wire[109];							inform_L[55][6] = l_cell_wire[110];							inform_L[119][6] = l_cell_wire[111];							inform_L[56][6] = l_cell_wire[112];							inform_L[120][6] = l_cell_wire[113];							inform_L[57][6] = l_cell_wire[114];							inform_L[121][6] = l_cell_wire[115];							inform_L[58][6] = l_cell_wire[116];							inform_L[122][6] = l_cell_wire[117];							inform_L[59][6] = l_cell_wire[118];							inform_L[123][6] = l_cell_wire[119];							inform_L[60][6] = l_cell_wire[120];							inform_L[124][6] = l_cell_wire[121];							inform_L[61][6] = l_cell_wire[122];							inform_L[125][6] = l_cell_wire[123];							inform_L[62][6] = l_cell_wire[124];							inform_L[126][6] = l_cell_wire[125];							inform_L[63][6] = l_cell_wire[126];							inform_L[127][6] = l_cell_wire[127];							inform_L[128][6] = l_cell_wire[128];							inform_L[192][6] = l_cell_wire[129];							inform_L[129][6] = l_cell_wire[130];							inform_L[193][6] = l_cell_wire[131];							inform_L[130][6] = l_cell_wire[132];							inform_L[194][6] = l_cell_wire[133];							inform_L[131][6] = l_cell_wire[134];							inform_L[195][6] = l_cell_wire[135];							inform_L[132][6] = l_cell_wire[136];							inform_L[196][6] = l_cell_wire[137];							inform_L[133][6] = l_cell_wire[138];							inform_L[197][6] = l_cell_wire[139];							inform_L[134][6] = l_cell_wire[140];							inform_L[198][6] = l_cell_wire[141];							inform_L[135][6] = l_cell_wire[142];							inform_L[199][6] = l_cell_wire[143];							inform_L[136][6] = l_cell_wire[144];							inform_L[200][6] = l_cell_wire[145];							inform_L[137][6] = l_cell_wire[146];							inform_L[201][6] = l_cell_wire[147];							inform_L[138][6] = l_cell_wire[148];							inform_L[202][6] = l_cell_wire[149];							inform_L[139][6] = l_cell_wire[150];							inform_L[203][6] = l_cell_wire[151];							inform_L[140][6] = l_cell_wire[152];							inform_L[204][6] = l_cell_wire[153];							inform_L[141][6] = l_cell_wire[154];							inform_L[205][6] = l_cell_wire[155];							inform_L[142][6] = l_cell_wire[156];							inform_L[206][6] = l_cell_wire[157];							inform_L[143][6] = l_cell_wire[158];							inform_L[207][6] = l_cell_wire[159];							inform_L[144][6] = l_cell_wire[160];							inform_L[208][6] = l_cell_wire[161];							inform_L[145][6] = l_cell_wire[162];							inform_L[209][6] = l_cell_wire[163];							inform_L[146][6] = l_cell_wire[164];							inform_L[210][6] = l_cell_wire[165];							inform_L[147][6] = l_cell_wire[166];							inform_L[211][6] = l_cell_wire[167];							inform_L[148][6] = l_cell_wire[168];							inform_L[212][6] = l_cell_wire[169];							inform_L[149][6] = l_cell_wire[170];							inform_L[213][6] = l_cell_wire[171];							inform_L[150][6] = l_cell_wire[172];							inform_L[214][6] = l_cell_wire[173];							inform_L[151][6] = l_cell_wire[174];							inform_L[215][6] = l_cell_wire[175];							inform_L[152][6] = l_cell_wire[176];							inform_L[216][6] = l_cell_wire[177];							inform_L[153][6] = l_cell_wire[178];							inform_L[217][6] = l_cell_wire[179];							inform_L[154][6] = l_cell_wire[180];							inform_L[218][6] = l_cell_wire[181];							inform_L[155][6] = l_cell_wire[182];							inform_L[219][6] = l_cell_wire[183];							inform_L[156][6] = l_cell_wire[184];							inform_L[220][6] = l_cell_wire[185];							inform_L[157][6] = l_cell_wire[186];							inform_L[221][6] = l_cell_wire[187];							inform_L[158][6] = l_cell_wire[188];							inform_L[222][6] = l_cell_wire[189];							inform_L[159][6] = l_cell_wire[190];							inform_L[223][6] = l_cell_wire[191];							inform_L[160][6] = l_cell_wire[192];							inform_L[224][6] = l_cell_wire[193];							inform_L[161][6] = l_cell_wire[194];							inform_L[225][6] = l_cell_wire[195];							inform_L[162][6] = l_cell_wire[196];							inform_L[226][6] = l_cell_wire[197];							inform_L[163][6] = l_cell_wire[198];							inform_L[227][6] = l_cell_wire[199];							inform_L[164][6] = l_cell_wire[200];							inform_L[228][6] = l_cell_wire[201];							inform_L[165][6] = l_cell_wire[202];							inform_L[229][6] = l_cell_wire[203];							inform_L[166][6] = l_cell_wire[204];							inform_L[230][6] = l_cell_wire[205];							inform_L[167][6] = l_cell_wire[206];							inform_L[231][6] = l_cell_wire[207];							inform_L[168][6] = l_cell_wire[208];							inform_L[232][6] = l_cell_wire[209];							inform_L[169][6] = l_cell_wire[210];							inform_L[233][6] = l_cell_wire[211];							inform_L[170][6] = l_cell_wire[212];							inform_L[234][6] = l_cell_wire[213];							inform_L[171][6] = l_cell_wire[214];							inform_L[235][6] = l_cell_wire[215];							inform_L[172][6] = l_cell_wire[216];							inform_L[236][6] = l_cell_wire[217];							inform_L[173][6] = l_cell_wire[218];							inform_L[237][6] = l_cell_wire[219];							inform_L[174][6] = l_cell_wire[220];							inform_L[238][6] = l_cell_wire[221];							inform_L[175][6] = l_cell_wire[222];							inform_L[239][6] = l_cell_wire[223];							inform_L[176][6] = l_cell_wire[224];							inform_L[240][6] = l_cell_wire[225];							inform_L[177][6] = l_cell_wire[226];							inform_L[241][6] = l_cell_wire[227];							inform_L[178][6] = l_cell_wire[228];							inform_L[242][6] = l_cell_wire[229];							inform_L[179][6] = l_cell_wire[230];							inform_L[243][6] = l_cell_wire[231];							inform_L[180][6] = l_cell_wire[232];							inform_L[244][6] = l_cell_wire[233];							inform_L[181][6] = l_cell_wire[234];							inform_L[245][6] = l_cell_wire[235];							inform_L[182][6] = l_cell_wire[236];							inform_L[246][6] = l_cell_wire[237];							inform_L[183][6] = l_cell_wire[238];							inform_L[247][6] = l_cell_wire[239];							inform_L[184][6] = l_cell_wire[240];							inform_L[248][6] = l_cell_wire[241];							inform_L[185][6] = l_cell_wire[242];							inform_L[249][6] = l_cell_wire[243];							inform_L[186][6] = l_cell_wire[244];							inform_L[250][6] = l_cell_wire[245];							inform_L[187][6] = l_cell_wire[246];							inform_L[251][6] = l_cell_wire[247];							inform_L[188][6] = l_cell_wire[248];							inform_L[252][6] = l_cell_wire[249];							inform_L[189][6] = l_cell_wire[250];							inform_L[253][6] = l_cell_wire[251];							inform_L[190][6] = l_cell_wire[252];							inform_L[254][6] = l_cell_wire[253];							inform_L[191][6] = l_cell_wire[254];							inform_L[255][6] = l_cell_wire[255];						end
						8:						begin							inform_R[0][8] = r_cell_wire[0];							inform_R[128][8] = r_cell_wire[1];							inform_R[1][8] = r_cell_wire[2];							inform_R[129][8] = r_cell_wire[3];							inform_R[2][8] = r_cell_wire[4];							inform_R[130][8] = r_cell_wire[5];							inform_R[3][8] = r_cell_wire[6];							inform_R[131][8] = r_cell_wire[7];							inform_R[4][8] = r_cell_wire[8];							inform_R[132][8] = r_cell_wire[9];							inform_R[5][8] = r_cell_wire[10];							inform_R[133][8] = r_cell_wire[11];							inform_R[6][8] = r_cell_wire[12];							inform_R[134][8] = r_cell_wire[13];							inform_R[7][8] = r_cell_wire[14];							inform_R[135][8] = r_cell_wire[15];							inform_R[8][8] = r_cell_wire[16];							inform_R[136][8] = r_cell_wire[17];							inform_R[9][8] = r_cell_wire[18];							inform_R[137][8] = r_cell_wire[19];							inform_R[10][8] = r_cell_wire[20];							inform_R[138][8] = r_cell_wire[21];							inform_R[11][8] = r_cell_wire[22];							inform_R[139][8] = r_cell_wire[23];							inform_R[12][8] = r_cell_wire[24];							inform_R[140][8] = r_cell_wire[25];							inform_R[13][8] = r_cell_wire[26];							inform_R[141][8] = r_cell_wire[27];							inform_R[14][8] = r_cell_wire[28];							inform_R[142][8] = r_cell_wire[29];							inform_R[15][8] = r_cell_wire[30];							inform_R[143][8] = r_cell_wire[31];							inform_R[16][8] = r_cell_wire[32];							inform_R[144][8] = r_cell_wire[33];							inform_R[17][8] = r_cell_wire[34];							inform_R[145][8] = r_cell_wire[35];							inform_R[18][8] = r_cell_wire[36];							inform_R[146][8] = r_cell_wire[37];							inform_R[19][8] = r_cell_wire[38];							inform_R[147][8] = r_cell_wire[39];							inform_R[20][8] = r_cell_wire[40];							inform_R[148][8] = r_cell_wire[41];							inform_R[21][8] = r_cell_wire[42];							inform_R[149][8] = r_cell_wire[43];							inform_R[22][8] = r_cell_wire[44];							inform_R[150][8] = r_cell_wire[45];							inform_R[23][8] = r_cell_wire[46];							inform_R[151][8] = r_cell_wire[47];							inform_R[24][8] = r_cell_wire[48];							inform_R[152][8] = r_cell_wire[49];							inform_R[25][8] = r_cell_wire[50];							inform_R[153][8] = r_cell_wire[51];							inform_R[26][8] = r_cell_wire[52];							inform_R[154][8] = r_cell_wire[53];							inform_R[27][8] = r_cell_wire[54];							inform_R[155][8] = r_cell_wire[55];							inform_R[28][8] = r_cell_wire[56];							inform_R[156][8] = r_cell_wire[57];							inform_R[29][8] = r_cell_wire[58];							inform_R[157][8] = r_cell_wire[59];							inform_R[30][8] = r_cell_wire[60];							inform_R[158][8] = r_cell_wire[61];							inform_R[31][8] = r_cell_wire[62];							inform_R[159][8] = r_cell_wire[63];							inform_R[32][8] = r_cell_wire[64];							inform_R[160][8] = r_cell_wire[65];							inform_R[33][8] = r_cell_wire[66];							inform_R[161][8] = r_cell_wire[67];							inform_R[34][8] = r_cell_wire[68];							inform_R[162][8] = r_cell_wire[69];							inform_R[35][8] = r_cell_wire[70];							inform_R[163][8] = r_cell_wire[71];							inform_R[36][8] = r_cell_wire[72];							inform_R[164][8] = r_cell_wire[73];							inform_R[37][8] = r_cell_wire[74];							inform_R[165][8] = r_cell_wire[75];							inform_R[38][8] = r_cell_wire[76];							inform_R[166][8] = r_cell_wire[77];							inform_R[39][8] = r_cell_wire[78];							inform_R[167][8] = r_cell_wire[79];							inform_R[40][8] = r_cell_wire[80];							inform_R[168][8] = r_cell_wire[81];							inform_R[41][8] = r_cell_wire[82];							inform_R[169][8] = r_cell_wire[83];							inform_R[42][8] = r_cell_wire[84];							inform_R[170][8] = r_cell_wire[85];							inform_R[43][8] = r_cell_wire[86];							inform_R[171][8] = r_cell_wire[87];							inform_R[44][8] = r_cell_wire[88];							inform_R[172][8] = r_cell_wire[89];							inform_R[45][8] = r_cell_wire[90];							inform_R[173][8] = r_cell_wire[91];							inform_R[46][8] = r_cell_wire[92];							inform_R[174][8] = r_cell_wire[93];							inform_R[47][8] = r_cell_wire[94];							inform_R[175][8] = r_cell_wire[95];							inform_R[48][8] = r_cell_wire[96];							inform_R[176][8] = r_cell_wire[97];							inform_R[49][8] = r_cell_wire[98];							inform_R[177][8] = r_cell_wire[99];							inform_R[50][8] = r_cell_wire[100];							inform_R[178][8] = r_cell_wire[101];							inform_R[51][8] = r_cell_wire[102];							inform_R[179][8] = r_cell_wire[103];							inform_R[52][8] = r_cell_wire[104];							inform_R[180][8] = r_cell_wire[105];							inform_R[53][8] = r_cell_wire[106];							inform_R[181][8] = r_cell_wire[107];							inform_R[54][8] = r_cell_wire[108];							inform_R[182][8] = r_cell_wire[109];							inform_R[55][8] = r_cell_wire[110];							inform_R[183][8] = r_cell_wire[111];							inform_R[56][8] = r_cell_wire[112];							inform_R[184][8] = r_cell_wire[113];							inform_R[57][8] = r_cell_wire[114];							inform_R[185][8] = r_cell_wire[115];							inform_R[58][8] = r_cell_wire[116];							inform_R[186][8] = r_cell_wire[117];							inform_R[59][8] = r_cell_wire[118];							inform_R[187][8] = r_cell_wire[119];							inform_R[60][8] = r_cell_wire[120];							inform_R[188][8] = r_cell_wire[121];							inform_R[61][8] = r_cell_wire[122];							inform_R[189][8] = r_cell_wire[123];							inform_R[62][8] = r_cell_wire[124];							inform_R[190][8] = r_cell_wire[125];							inform_R[63][8] = r_cell_wire[126];							inform_R[191][8] = r_cell_wire[127];							inform_R[64][8] = r_cell_wire[128];							inform_R[192][8] = r_cell_wire[129];							inform_R[65][8] = r_cell_wire[130];							inform_R[193][8] = r_cell_wire[131];							inform_R[66][8] = r_cell_wire[132];							inform_R[194][8] = r_cell_wire[133];							inform_R[67][8] = r_cell_wire[134];							inform_R[195][8] = r_cell_wire[135];							inform_R[68][8] = r_cell_wire[136];							inform_R[196][8] = r_cell_wire[137];							inform_R[69][8] = r_cell_wire[138];							inform_R[197][8] = r_cell_wire[139];							inform_R[70][8] = r_cell_wire[140];							inform_R[198][8] = r_cell_wire[141];							inform_R[71][8] = r_cell_wire[142];							inform_R[199][8] = r_cell_wire[143];							inform_R[72][8] = r_cell_wire[144];							inform_R[200][8] = r_cell_wire[145];							inform_R[73][8] = r_cell_wire[146];							inform_R[201][8] = r_cell_wire[147];							inform_R[74][8] = r_cell_wire[148];							inform_R[202][8] = r_cell_wire[149];							inform_R[75][8] = r_cell_wire[150];							inform_R[203][8] = r_cell_wire[151];							inform_R[76][8] = r_cell_wire[152];							inform_R[204][8] = r_cell_wire[153];							inform_R[77][8] = r_cell_wire[154];							inform_R[205][8] = r_cell_wire[155];							inform_R[78][8] = r_cell_wire[156];							inform_R[206][8] = r_cell_wire[157];							inform_R[79][8] = r_cell_wire[158];							inform_R[207][8] = r_cell_wire[159];							inform_R[80][8] = r_cell_wire[160];							inform_R[208][8] = r_cell_wire[161];							inform_R[81][8] = r_cell_wire[162];							inform_R[209][8] = r_cell_wire[163];							inform_R[82][8] = r_cell_wire[164];							inform_R[210][8] = r_cell_wire[165];							inform_R[83][8] = r_cell_wire[166];							inform_R[211][8] = r_cell_wire[167];							inform_R[84][8] = r_cell_wire[168];							inform_R[212][8] = r_cell_wire[169];							inform_R[85][8] = r_cell_wire[170];							inform_R[213][8] = r_cell_wire[171];							inform_R[86][8] = r_cell_wire[172];							inform_R[214][8] = r_cell_wire[173];							inform_R[87][8] = r_cell_wire[174];							inform_R[215][8] = r_cell_wire[175];							inform_R[88][8] = r_cell_wire[176];							inform_R[216][8] = r_cell_wire[177];							inform_R[89][8] = r_cell_wire[178];							inform_R[217][8] = r_cell_wire[179];							inform_R[90][8] = r_cell_wire[180];							inform_R[218][8] = r_cell_wire[181];							inform_R[91][8] = r_cell_wire[182];							inform_R[219][8] = r_cell_wire[183];							inform_R[92][8] = r_cell_wire[184];							inform_R[220][8] = r_cell_wire[185];							inform_R[93][8] = r_cell_wire[186];							inform_R[221][8] = r_cell_wire[187];							inform_R[94][8] = r_cell_wire[188];							inform_R[222][8] = r_cell_wire[189];							inform_R[95][8] = r_cell_wire[190];							inform_R[223][8] = r_cell_wire[191];							inform_R[96][8] = r_cell_wire[192];							inform_R[224][8] = r_cell_wire[193];							inform_R[97][8] = r_cell_wire[194];							inform_R[225][8] = r_cell_wire[195];							inform_R[98][8] = r_cell_wire[196];							inform_R[226][8] = r_cell_wire[197];							inform_R[99][8] = r_cell_wire[198];							inform_R[227][8] = r_cell_wire[199];							inform_R[100][8] = r_cell_wire[200];							inform_R[228][8] = r_cell_wire[201];							inform_R[101][8] = r_cell_wire[202];							inform_R[229][8] = r_cell_wire[203];							inform_R[102][8] = r_cell_wire[204];							inform_R[230][8] = r_cell_wire[205];							inform_R[103][8] = r_cell_wire[206];							inform_R[231][8] = r_cell_wire[207];							inform_R[104][8] = r_cell_wire[208];							inform_R[232][8] = r_cell_wire[209];							inform_R[105][8] = r_cell_wire[210];							inform_R[233][8] = r_cell_wire[211];							inform_R[106][8] = r_cell_wire[212];							inform_R[234][8] = r_cell_wire[213];							inform_R[107][8] = r_cell_wire[214];							inform_R[235][8] = r_cell_wire[215];							inform_R[108][8] = r_cell_wire[216];							inform_R[236][8] = r_cell_wire[217];							inform_R[109][8] = r_cell_wire[218];							inform_R[237][8] = r_cell_wire[219];							inform_R[110][8] = r_cell_wire[220];							inform_R[238][8] = r_cell_wire[221];							inform_R[111][8] = r_cell_wire[222];							inform_R[239][8] = r_cell_wire[223];							inform_R[112][8] = r_cell_wire[224];							inform_R[240][8] = r_cell_wire[225];							inform_R[113][8] = r_cell_wire[226];							inform_R[241][8] = r_cell_wire[227];							inform_R[114][8] = r_cell_wire[228];							inform_R[242][8] = r_cell_wire[229];							inform_R[115][8] = r_cell_wire[230];							inform_R[243][8] = r_cell_wire[231];							inform_R[116][8] = r_cell_wire[232];							inform_R[244][8] = r_cell_wire[233];							inform_R[117][8] = r_cell_wire[234];							inform_R[245][8] = r_cell_wire[235];							inform_R[118][8] = r_cell_wire[236];							inform_R[246][8] = r_cell_wire[237];							inform_R[119][8] = r_cell_wire[238];							inform_R[247][8] = r_cell_wire[239];							inform_R[120][8] = r_cell_wire[240];							inform_R[248][8] = r_cell_wire[241];							inform_R[121][8] = r_cell_wire[242];							inform_R[249][8] = r_cell_wire[243];							inform_R[122][8] = r_cell_wire[244];							inform_R[250][8] = r_cell_wire[245];							inform_R[123][8] = r_cell_wire[246];							inform_R[251][8] = r_cell_wire[247];							inform_R[124][8] = r_cell_wire[248];							inform_R[252][8] = r_cell_wire[249];							inform_R[125][8] = r_cell_wire[250];							inform_R[253][8] = r_cell_wire[251];							inform_R[126][8] = r_cell_wire[252];							inform_R[254][8] = r_cell_wire[253];							inform_R[127][8] = r_cell_wire[254];							inform_R[255][8] = r_cell_wire[255];							inform_L[0][7] = l_cell_wire[0];							inform_L[128][7] = l_cell_wire[1];							inform_L[1][7] = l_cell_wire[2];							inform_L[129][7] = l_cell_wire[3];							inform_L[2][7] = l_cell_wire[4];							inform_L[130][7] = l_cell_wire[5];							inform_L[3][7] = l_cell_wire[6];							inform_L[131][7] = l_cell_wire[7];							inform_L[4][7] = l_cell_wire[8];							inform_L[132][7] = l_cell_wire[9];							inform_L[5][7] = l_cell_wire[10];							inform_L[133][7] = l_cell_wire[11];							inform_L[6][7] = l_cell_wire[12];							inform_L[134][7] = l_cell_wire[13];							inform_L[7][7] = l_cell_wire[14];							inform_L[135][7] = l_cell_wire[15];							inform_L[8][7] = l_cell_wire[16];							inform_L[136][7] = l_cell_wire[17];							inform_L[9][7] = l_cell_wire[18];							inform_L[137][7] = l_cell_wire[19];							inform_L[10][7] = l_cell_wire[20];							inform_L[138][7] = l_cell_wire[21];							inform_L[11][7] = l_cell_wire[22];							inform_L[139][7] = l_cell_wire[23];							inform_L[12][7] = l_cell_wire[24];							inform_L[140][7] = l_cell_wire[25];							inform_L[13][7] = l_cell_wire[26];							inform_L[141][7] = l_cell_wire[27];							inform_L[14][7] = l_cell_wire[28];							inform_L[142][7] = l_cell_wire[29];							inform_L[15][7] = l_cell_wire[30];							inform_L[143][7] = l_cell_wire[31];							inform_L[16][7] = l_cell_wire[32];							inform_L[144][7] = l_cell_wire[33];							inform_L[17][7] = l_cell_wire[34];							inform_L[145][7] = l_cell_wire[35];							inform_L[18][7] = l_cell_wire[36];							inform_L[146][7] = l_cell_wire[37];							inform_L[19][7] = l_cell_wire[38];							inform_L[147][7] = l_cell_wire[39];							inform_L[20][7] = l_cell_wire[40];							inform_L[148][7] = l_cell_wire[41];							inform_L[21][7] = l_cell_wire[42];							inform_L[149][7] = l_cell_wire[43];							inform_L[22][7] = l_cell_wire[44];							inform_L[150][7] = l_cell_wire[45];							inform_L[23][7] = l_cell_wire[46];							inform_L[151][7] = l_cell_wire[47];							inform_L[24][7] = l_cell_wire[48];							inform_L[152][7] = l_cell_wire[49];							inform_L[25][7] = l_cell_wire[50];							inform_L[153][7] = l_cell_wire[51];							inform_L[26][7] = l_cell_wire[52];							inform_L[154][7] = l_cell_wire[53];							inform_L[27][7] = l_cell_wire[54];							inform_L[155][7] = l_cell_wire[55];							inform_L[28][7] = l_cell_wire[56];							inform_L[156][7] = l_cell_wire[57];							inform_L[29][7] = l_cell_wire[58];							inform_L[157][7] = l_cell_wire[59];							inform_L[30][7] = l_cell_wire[60];							inform_L[158][7] = l_cell_wire[61];							inform_L[31][7] = l_cell_wire[62];							inform_L[159][7] = l_cell_wire[63];							inform_L[32][7] = l_cell_wire[64];							inform_L[160][7] = l_cell_wire[65];							inform_L[33][7] = l_cell_wire[66];							inform_L[161][7] = l_cell_wire[67];							inform_L[34][7] = l_cell_wire[68];							inform_L[162][7] = l_cell_wire[69];							inform_L[35][7] = l_cell_wire[70];							inform_L[163][7] = l_cell_wire[71];							inform_L[36][7] = l_cell_wire[72];							inform_L[164][7] = l_cell_wire[73];							inform_L[37][7] = l_cell_wire[74];							inform_L[165][7] = l_cell_wire[75];							inform_L[38][7] = l_cell_wire[76];							inform_L[166][7] = l_cell_wire[77];							inform_L[39][7] = l_cell_wire[78];							inform_L[167][7] = l_cell_wire[79];							inform_L[40][7] = l_cell_wire[80];							inform_L[168][7] = l_cell_wire[81];							inform_L[41][7] = l_cell_wire[82];							inform_L[169][7] = l_cell_wire[83];							inform_L[42][7] = l_cell_wire[84];							inform_L[170][7] = l_cell_wire[85];							inform_L[43][7] = l_cell_wire[86];							inform_L[171][7] = l_cell_wire[87];							inform_L[44][7] = l_cell_wire[88];							inform_L[172][7] = l_cell_wire[89];							inform_L[45][7] = l_cell_wire[90];							inform_L[173][7] = l_cell_wire[91];							inform_L[46][7] = l_cell_wire[92];							inform_L[174][7] = l_cell_wire[93];							inform_L[47][7] = l_cell_wire[94];							inform_L[175][7] = l_cell_wire[95];							inform_L[48][7] = l_cell_wire[96];							inform_L[176][7] = l_cell_wire[97];							inform_L[49][7] = l_cell_wire[98];							inform_L[177][7] = l_cell_wire[99];							inform_L[50][7] = l_cell_wire[100];							inform_L[178][7] = l_cell_wire[101];							inform_L[51][7] = l_cell_wire[102];							inform_L[179][7] = l_cell_wire[103];							inform_L[52][7] = l_cell_wire[104];							inform_L[180][7] = l_cell_wire[105];							inform_L[53][7] = l_cell_wire[106];							inform_L[181][7] = l_cell_wire[107];							inform_L[54][7] = l_cell_wire[108];							inform_L[182][7] = l_cell_wire[109];							inform_L[55][7] = l_cell_wire[110];							inform_L[183][7] = l_cell_wire[111];							inform_L[56][7] = l_cell_wire[112];							inform_L[184][7] = l_cell_wire[113];							inform_L[57][7] = l_cell_wire[114];							inform_L[185][7] = l_cell_wire[115];							inform_L[58][7] = l_cell_wire[116];							inform_L[186][7] = l_cell_wire[117];							inform_L[59][7] = l_cell_wire[118];							inform_L[187][7] = l_cell_wire[119];							inform_L[60][7] = l_cell_wire[120];							inform_L[188][7] = l_cell_wire[121];							inform_L[61][7] = l_cell_wire[122];							inform_L[189][7] = l_cell_wire[123];							inform_L[62][7] = l_cell_wire[124];							inform_L[190][7] = l_cell_wire[125];							inform_L[63][7] = l_cell_wire[126];							inform_L[191][7] = l_cell_wire[127];							inform_L[64][7] = l_cell_wire[128];							inform_L[192][7] = l_cell_wire[129];							inform_L[65][7] = l_cell_wire[130];							inform_L[193][7] = l_cell_wire[131];							inform_L[66][7] = l_cell_wire[132];							inform_L[194][7] = l_cell_wire[133];							inform_L[67][7] = l_cell_wire[134];							inform_L[195][7] = l_cell_wire[135];							inform_L[68][7] = l_cell_wire[136];							inform_L[196][7] = l_cell_wire[137];							inform_L[69][7] = l_cell_wire[138];							inform_L[197][7] = l_cell_wire[139];							inform_L[70][7] = l_cell_wire[140];							inform_L[198][7] = l_cell_wire[141];							inform_L[71][7] = l_cell_wire[142];							inform_L[199][7] = l_cell_wire[143];							inform_L[72][7] = l_cell_wire[144];							inform_L[200][7] = l_cell_wire[145];							inform_L[73][7] = l_cell_wire[146];							inform_L[201][7] = l_cell_wire[147];							inform_L[74][7] = l_cell_wire[148];							inform_L[202][7] = l_cell_wire[149];							inform_L[75][7] = l_cell_wire[150];							inform_L[203][7] = l_cell_wire[151];							inform_L[76][7] = l_cell_wire[152];							inform_L[204][7] = l_cell_wire[153];							inform_L[77][7] = l_cell_wire[154];							inform_L[205][7] = l_cell_wire[155];							inform_L[78][7] = l_cell_wire[156];							inform_L[206][7] = l_cell_wire[157];							inform_L[79][7] = l_cell_wire[158];							inform_L[207][7] = l_cell_wire[159];							inform_L[80][7] = l_cell_wire[160];							inform_L[208][7] = l_cell_wire[161];							inform_L[81][7] = l_cell_wire[162];							inform_L[209][7] = l_cell_wire[163];							inform_L[82][7] = l_cell_wire[164];							inform_L[210][7] = l_cell_wire[165];							inform_L[83][7] = l_cell_wire[166];							inform_L[211][7] = l_cell_wire[167];							inform_L[84][7] = l_cell_wire[168];							inform_L[212][7] = l_cell_wire[169];							inform_L[85][7] = l_cell_wire[170];							inform_L[213][7] = l_cell_wire[171];							inform_L[86][7] = l_cell_wire[172];							inform_L[214][7] = l_cell_wire[173];							inform_L[87][7] = l_cell_wire[174];							inform_L[215][7] = l_cell_wire[175];							inform_L[88][7] = l_cell_wire[176];							inform_L[216][7] = l_cell_wire[177];							inform_L[89][7] = l_cell_wire[178];							inform_L[217][7] = l_cell_wire[179];							inform_L[90][7] = l_cell_wire[180];							inform_L[218][7] = l_cell_wire[181];							inform_L[91][7] = l_cell_wire[182];							inform_L[219][7] = l_cell_wire[183];							inform_L[92][7] = l_cell_wire[184];							inform_L[220][7] = l_cell_wire[185];							inform_L[93][7] = l_cell_wire[186];							inform_L[221][7] = l_cell_wire[187];							inform_L[94][7] = l_cell_wire[188];							inform_L[222][7] = l_cell_wire[189];							inform_L[95][7] = l_cell_wire[190];							inform_L[223][7] = l_cell_wire[191];							inform_L[96][7] = l_cell_wire[192];							inform_L[224][7] = l_cell_wire[193];							inform_L[97][7] = l_cell_wire[194];							inform_L[225][7] = l_cell_wire[195];							inform_L[98][7] = l_cell_wire[196];							inform_L[226][7] = l_cell_wire[197];							inform_L[99][7] = l_cell_wire[198];							inform_L[227][7] = l_cell_wire[199];							inform_L[100][7] = l_cell_wire[200];							inform_L[228][7] = l_cell_wire[201];							inform_L[101][7] = l_cell_wire[202];							inform_L[229][7] = l_cell_wire[203];							inform_L[102][7] = l_cell_wire[204];							inform_L[230][7] = l_cell_wire[205];							inform_L[103][7] = l_cell_wire[206];							inform_L[231][7] = l_cell_wire[207];							inform_L[104][7] = l_cell_wire[208];							inform_L[232][7] = l_cell_wire[209];							inform_L[105][7] = l_cell_wire[210];							inform_L[233][7] = l_cell_wire[211];							inform_L[106][7] = l_cell_wire[212];							inform_L[234][7] = l_cell_wire[213];							inform_L[107][7] = l_cell_wire[214];							inform_L[235][7] = l_cell_wire[215];							inform_L[108][7] = l_cell_wire[216];							inform_L[236][7] = l_cell_wire[217];							inform_L[109][7] = l_cell_wire[218];							inform_L[237][7] = l_cell_wire[219];							inform_L[110][7] = l_cell_wire[220];							inform_L[238][7] = l_cell_wire[221];							inform_L[111][7] = l_cell_wire[222];							inform_L[239][7] = l_cell_wire[223];							inform_L[112][7] = l_cell_wire[224];							inform_L[240][7] = l_cell_wire[225];							inform_L[113][7] = l_cell_wire[226];							inform_L[241][7] = l_cell_wire[227];							inform_L[114][7] = l_cell_wire[228];							inform_L[242][7] = l_cell_wire[229];							inform_L[115][7] = l_cell_wire[230];							inform_L[243][7] = l_cell_wire[231];							inform_L[116][7] = l_cell_wire[232];							inform_L[244][7] = l_cell_wire[233];							inform_L[117][7] = l_cell_wire[234];							inform_L[245][7] = l_cell_wire[235];							inform_L[118][7] = l_cell_wire[236];							inform_L[246][7] = l_cell_wire[237];							inform_L[119][7] = l_cell_wire[238];							inform_L[247][7] = l_cell_wire[239];							inform_L[120][7] = l_cell_wire[240];							inform_L[248][7] = l_cell_wire[241];							inform_L[121][7] = l_cell_wire[242];							inform_L[249][7] = l_cell_wire[243];							inform_L[122][7] = l_cell_wire[244];							inform_L[250][7] = l_cell_wire[245];							inform_L[123][7] = l_cell_wire[246];							inform_L[251][7] = l_cell_wire[247];							inform_L[124][7] = l_cell_wire[248];							inform_L[252][7] = l_cell_wire[249];							inform_L[125][7] = l_cell_wire[250];							inform_L[253][7] = l_cell_wire[251];							inform_L[126][7] = l_cell_wire[252];							inform_L[254][7] = l_cell_wire[253];							inform_L[127][7] = l_cell_wire[254];							inform_L[255][7] = l_cell_wire[255];						end
						default:							for (x = 0; x < 256; x = x + 1)								for (y = 0; y < 8; y = y + 1)								begin									inform_R[x][y+1] <= 8'd0;									inform_L[x][y] <= 8'd0;								end					endcase				end			end
				default:				begin				if (start) begin					inform_R [0][0] <= 8'b0111_1111;					inform_R [1][0] <= 8'b0111_1111;					inform_R [2][0] <= 8'b0111_1111;					inform_R [3][0] <= 8'b0111_1111;					inform_R [4][0] <= 8'b0111_1111;					inform_R [5][0] <= 8'b0111_1111;					inform_R [6][0] <= 8'b0111_1111;					inform_R [7][0] <= 8'b0111_1111;					inform_R [8][0] <= 8'b0111_1111;					inform_R [9][0] <= 8'b0111_1111;					inform_R [10][0] <= 8'b0111_1111;					inform_R [11][0] <= 8'b0111_1111;					inform_R [12][0] <= 8'b0111_1111;					inform_R [13][0] <= 8'b0111_1111;					inform_R [14][0] <= 8'b0111_1111;					inform_R [15][0] <= 8'b0111_1111;					inform_R [16][0] <= 8'b0111_1111;					inform_R [17][0] <= 8'b0111_1111;					inform_R [18][0] <= 8'b0111_1111;					inform_R [19][0] <= 8'b0111_1111;					inform_R [20][0] <= 8'b0111_1111;					inform_R [21][0] <= 8'b0111_1111;					inform_R [22][0] <= 8'b0111_1111;					inform_R [23][0] <= 8'b0111_1111;					inform_R [24][0] <= 8'b0111_1111;					inform_R [25][0] <= 8'b0111_1111;					inform_R [26][0] <= 8'b0111_1111;					inform_R [27][0] <= 8'b0111_1111;					inform_R [28][0] <= 8'b0111_1111;					inform_R [29][0] <= 8'b0111_1111;					inform_R [30][0] <= 8'b0111_1111;					inform_R [31][0] <= 8'b0111_1111;					inform_R [32][0] <= 8'b0111_1111;					inform_R [33][0] <= 8'b0111_1111;					inform_R [34][0] <= 8'b0111_1111;					inform_R [35][0] <= 8'b0111_1111;					inform_R [36][0] <= 8'b0111_1111;					inform_R [37][0] <= 8'b0111_1111;					inform_R [38][0] <= 8'b0111_1111;					inform_R [39][0] <= 8'b0111_1111;					inform_R [40][0] <= 8'b0111_1111;					inform_R [41][0] <= 8'b0111_1111;					inform_R [42][0] <= 8'b0111_1111;					inform_R [43][0] <= 8'b0111_1111;					inform_R [44][0] <= 8'b0111_1111;					inform_R [45][0] <= 8'b0111_1111;					inform_R [46][0] <= 8'b0111_1111;					inform_R [47][0] <= 8'b0111_1111;					inform_R [48][0] <= 8'b0111_1111;					inform_R [49][0] <= 8'b0111_1111;					inform_R [50][0] <= 8'b0111_1111;					inform_R [51][0] <= 8'b0111_1111;					inform_R [52][0] <= 8'b0111_1111;					inform_R [53][0] <= 8'b0111_1111;					inform_R [54][0] <= 8'b0111_1111;					inform_R [55][0] <= 8'b0111_1111;					inform_R [56][0] <= 8'b0111_1111;					inform_R [57][0] <= 8'b0111_1111;					inform_R [58][0] <= 8'b0111_1111;					inform_R [59][0] <= 8'b0000_0000;					inform_R [60][0] <= 8'b0111_1111;					inform_R [61][0] <= 8'b0000_0000;					inform_R [62][0] <= 8'b0000_0000;					inform_R [63][0] <= 8'b0000_0000;					inform_R [64][0] <= 8'b0111_1111;					inform_R [65][0] <= 8'b0111_1111;					inform_R [66][0] <= 8'b0111_1111;					inform_R [67][0] <= 8'b0111_1111;					inform_R [68][0] <= 8'b0111_1111;					inform_R [69][0] <= 8'b0111_1111;					inform_R [70][0] <= 8'b0111_1111;					inform_R [71][0] <= 8'b0111_1111;					inform_R [72][0] <= 8'b0111_1111;					inform_R [73][0] <= 8'b0111_1111;					inform_R [74][0] <= 8'b0111_1111;					inform_R [75][0] <= 8'b0111_1111;					inform_R [76][0] <= 8'b0111_1111;					inform_R [77][0] <= 8'b0111_1111;					inform_R [78][0] <= 8'b0111_1111;					inform_R [79][0] <= 8'b0111_1111;					inform_R [80][0] <= 8'b0111_1111;					inform_R [81][0] <= 8'b0111_1111;					inform_R [82][0] <= 8'b0111_1111;					inform_R [83][0] <= 8'b0111_1111;					inform_R [84][0] <= 8'b0111_1111;					inform_R [85][0] <= 8'b0111_1111;					inform_R [86][0] <= 8'b0111_1111;					inform_R [87][0] <= 8'b0000_0000;					inform_R [88][0] <= 8'b0111_1111;					inform_R [89][0] <= 8'b0111_1111;					inform_R [90][0] <= 8'b0111_1111;					inform_R [91][0] <= 8'b0000_0000;					inform_R [92][0] <= 8'b0111_1111;					inform_R [93][0] <= 8'b0000_0000;					inform_R [94][0] <= 8'b0000_0000;					inform_R [95][0] <= 8'b0000_0000;					inform_R [96][0] <= 8'b0111_1111;					inform_R [97][0] <= 8'b0111_1111;					inform_R [98][0] <= 8'b0111_1111;					inform_R [99][0] <= 8'b0111_1111;					inform_R [100][0] <= 8'b0111_1111;					inform_R [101][0] <= 8'b0111_1111;					inform_R [102][0] <= 8'b0111_1111;					inform_R [103][0] <= 8'b0000_0000;					inform_R [104][0] <= 8'b0111_1111;					inform_R [105][0] <= 8'b0111_1111;					inform_R [106][0] <= 8'b0000_0000;					inform_R [107][0] <= 8'b0000_0000;					inform_R [108][0] <= 8'b0000_0000;					inform_R [109][0] <= 8'b0000_0000;					inform_R [110][0] <= 8'b0000_0000;					inform_R [111][0] <= 8'b0000_0000;					inform_R [112][0] <= 8'b0111_1111;					inform_R [113][0] <= 8'b0000_0000;					inform_R [114][0] <= 8'b0000_0000;					inform_R [115][0] <= 8'b0000_0000;					inform_R [116][0] <= 8'b0000_0000;					inform_R [117][0] <= 8'b0000_0000;					inform_R [118][0] <= 8'b0000_0000;					inform_R [119][0] <= 8'b0000_0000;					inform_R [120][0] <= 8'b0000_0000;					inform_R [121][0] <= 8'b0000_0000;					inform_R [122][0] <= 8'b0000_0000;					inform_R [123][0] <= 8'b0000_0000;					inform_R [124][0] <= 8'b0000_0000;					inform_R [125][0] <= 8'b0000_0000;					inform_R [126][0] <= 8'b0000_0000;					inform_R [127][0] <= 8'b0000_0000;					inform_R [128][0] <= 8'b0111_1111;					inform_R [129][0] <= 8'b0111_1111;					inform_R [130][0] <= 8'b0111_1111;					inform_R [131][0] <= 8'b0111_1111;					inform_R [132][0] <= 8'b0111_1111;					inform_R [133][0] <= 8'b0111_1111;					inform_R [134][0] <= 8'b0111_1111;					inform_R [135][0] <= 8'b0111_1111;					inform_R [136][0] <= 8'b0111_1111;					inform_R [137][0] <= 8'b0111_1111;					inform_R [138][0] <= 8'b0111_1111;					inform_R [139][0] <= 8'b0111_1111;					inform_R [140][0] <= 8'b0111_1111;					inform_R [141][0] <= 8'b0111_1111;					inform_R [142][0] <= 8'b0111_1111;					inform_R [143][0] <= 8'b0000_0000;					inform_R [144][0] <= 8'b0111_1111;					inform_R [145][0] <= 8'b0111_1111;					inform_R [146][0] <= 8'b0111_1111;					inform_R [147][0] <= 8'b0111_1111;					inform_R [148][0] <= 8'b0111_1111;					inform_R [149][0] <= 8'b0111_1111;					inform_R [150][0] <= 8'b0000_0000;					inform_R [151][0] <= 8'b0000_0000;					inform_R [152][0] <= 8'b0111_1111;					inform_R [153][0] <= 8'b0000_0000;					inform_R [154][0] <= 8'b0000_0000;					inform_R [155][0] <= 8'b0000_0000;					inform_R [156][0] <= 8'b0000_0000;					inform_R [157][0] <= 8'b0000_0000;					inform_R [158][0] <= 8'b0000_0000;					inform_R [159][0] <= 8'b0000_0000;					inform_R [160][0] <= 8'b0111_1111;					inform_R [161][0] <= 8'b0111_1111;					inform_R [162][0] <= 8'b0111_1111;					inform_R [163][0] <= 8'b0000_0000;					inform_R [164][0] <= 8'b0111_1111;					inform_R [165][0] <= 8'b0000_0000;					inform_R [166][0] <= 8'b0000_0000;					inform_R [167][0] <= 8'b0000_0000;					inform_R [168][0] <= 8'b0111_1111;					inform_R [169][0] <= 8'b0000_0000;					inform_R [170][0] <= 8'b0000_0000;					inform_R [171][0] <= 8'b0000_0000;					inform_R [172][0] <= 8'b0000_0000;					inform_R [173][0] <= 8'b0000_0000;					inform_R [174][0] <= 8'b0000_0000;					inform_R [175][0] <= 8'b0000_0000;					inform_R [176][0] <= 8'b0000_0000;					inform_R [177][0] <= 8'b0000_0000;					inform_R [178][0] <= 8'b0000_0000;					inform_R [179][0] <= 8'b0000_0000;					inform_R [180][0] <= 8'b0000_0000;					inform_R [181][0] <= 8'b0000_0000;					inform_R [182][0] <= 8'b0000_0000;					inform_R [183][0] <= 8'b0000_0000;					inform_R [184][0] <= 8'b0000_0000;					inform_R [185][0] <= 8'b0000_0000;					inform_R [186][0] <= 8'b0000_0000;					inform_R [187][0] <= 8'b0000_0000;					inform_R [188][0] <= 8'b0000_0000;					inform_R [189][0] <= 8'b0000_0000;					inform_R [190][0] <= 8'b0000_0000;					inform_R [191][0] <= 8'b0000_0000;					inform_R [192][0] <= 8'b0111_1111;					inform_R [193][0] <= 8'b0111_1111;					inform_R [194][0] <= 8'b0111_1111;					inform_R [195][0] <= 8'b0000_0000;					inform_R [196][0] <= 8'b0111_1111;					inform_R [197][0] <= 8'b0000_0000;					inform_R [198][0] <= 8'b0000_0000;					inform_R [199][0] <= 8'b0000_0000;					inform_R [200][0] <= 8'b0000_0000;					inform_R [201][0] <= 8'b0000_0000;					inform_R [202][0] <= 8'b0000_0000;					inform_R [203][0] <= 8'b0000_0000;					inform_R [204][0] <= 8'b0000_0000;					inform_R [205][0] <= 8'b0000_0000;					inform_R [206][0] <= 8'b0000_0000;					inform_R [207][0] <= 8'b0000_0000;					inform_R [208][0] <= 8'b0000_0000;					inform_R [209][0] <= 8'b0000_0000;					inform_R [210][0] <= 8'b0000_0000;					inform_R [211][0] <= 8'b0000_0000;					inform_R [212][0] <= 8'b0000_0000;					inform_R [213][0] <= 8'b0000_0000;					inform_R [214][0] <= 8'b0000_0000;					inform_R [215][0] <= 8'b0000_0000;					inform_R [216][0] <= 8'b0000_0000;					inform_R [217][0] <= 8'b0000_0000;					inform_R [218][0] <= 8'b0000_0000;					inform_R [219][0] <= 8'b0000_0000;					inform_R [220][0] <= 8'b0000_0000;					inform_R [221][0] <= 8'b0000_0000;					inform_R [222][0] <= 8'b0000_0000;					inform_R [223][0] <= 8'b0000_0000;					inform_R [224][0] <= 8'b0000_0000;					inform_R [225][0] <= 8'b0000_0000;					inform_R [226][0] <= 8'b0000_0000;					inform_R [227][0] <= 8'b0000_0000;					inform_R [228][0] <= 8'b0000_0000;					inform_R [229][0] <= 8'b0000_0000;					inform_R [230][0] <= 8'b0000_0000;					inform_R [231][0] <= 8'b0000_0000;					inform_R [232][0] <= 8'b0000_0000;					inform_R [233][0] <= 8'b0000_0000;					inform_R [234][0] <= 8'b0000_0000;					inform_R [235][0] <= 8'b0000_0000;					inform_R [236][0] <= 8'b0000_0000;					inform_R [237][0] <= 8'b0000_0000;					inform_R [238][0] <= 8'b0000_0000;					inform_R [239][0] <= 8'b0000_0000;					inform_R [240][0] <= 8'b0000_0000;					inform_R [241][0] <= 8'b0000_0000;					inform_R [242][0] <= 8'b0000_0000;					inform_R [243][0] <= 8'b0000_0000;					inform_R [244][0] <= 8'b0000_0000;					inform_R [245][0] <= 8'b0000_0000;					inform_R [246][0] <= 8'b0000_0000;					inform_R [247][0] <= 8'b0000_0000;					inform_R [248][0] <= 8'b0000_0000;					inform_R [249][0] <= 8'b0000_0000;					inform_R [250][0] <= 8'b0000_0000;					inform_R [251][0] <= 8'b0000_0000;					inform_R [252][0] <= 8'b0000_0000;					inform_R [253][0] <= 8'b0000_0000;					inform_R [254][0] <= 8'b0000_0000;					inform_R [255][0] <= 8'b0000_0000;					inform_L [0][8] <= LLR_1;					inform_L [1][8] <= LLR_2;					inform_L [2][8] <= LLR_3;					inform_L [3][8] <= LLR_4;					inform_L [4][8] <= LLR_5;					inform_L [5][8] <= LLR_6;					inform_L [6][8] <= LLR_7;					inform_L [7][8] <= LLR_8;					inform_L [8][8] <= LLR_9;					inform_L [9][8] <= LLR_10;					inform_L [10][8] <= LLR_11;					inform_L [11][8] <= LLR_12;					inform_L [12][8] <= LLR_13;					inform_L [13][8] <= LLR_14;					inform_L [14][8] <= LLR_15;					inform_L [15][8] <= LLR_16;					inform_L [16][8] <= LLR_17;					inform_L [17][8] <= LLR_18;					inform_L [18][8] <= LLR_19;					inform_L [19][8] <= LLR_20;					inform_L [20][8] <= LLR_21;					inform_L [21][8] <= LLR_22;					inform_L [22][8] <= LLR_23;					inform_L [23][8] <= LLR_24;					inform_L [24][8] <= LLR_25;					inform_L [25][8] <= LLR_26;					inform_L [26][8] <= LLR_27;					inform_L [27][8] <= LLR_28;					inform_L [28][8] <= LLR_29;					inform_L [29][8] <= LLR_30;					inform_L [30][8] <= LLR_31;					inform_L [31][8] <= LLR_32;					inform_L [32][8] <= LLR_33;					inform_L [33][8] <= LLR_34;					inform_L [34][8] <= LLR_35;					inform_L [35][8] <= LLR_36;					inform_L [36][8] <= LLR_37;					inform_L [37][8] <= LLR_38;					inform_L [38][8] <= LLR_39;					inform_L [39][8] <= LLR_40;					inform_L [40][8] <= LLR_41;					inform_L [41][8] <= LLR_42;					inform_L [42][8] <= LLR_43;					inform_L [43][8] <= LLR_44;					inform_L [44][8] <= LLR_45;					inform_L [45][8] <= LLR_46;					inform_L [46][8] <= LLR_47;					inform_L [47][8] <= LLR_48;					inform_L [48][8] <= LLR_49;					inform_L [49][8] <= LLR_50;					inform_L [50][8] <= LLR_51;					inform_L [51][8] <= LLR_52;					inform_L [52][8] <= LLR_53;					inform_L [53][8] <= LLR_54;					inform_L [54][8] <= LLR_55;					inform_L [55][8] <= LLR_56;					inform_L [56][8] <= LLR_57;					inform_L [57][8] <= LLR_58;					inform_L [58][8] <= LLR_59;					inform_L [59][8] <= LLR_60;					inform_L [60][8] <= LLR_61;					inform_L [61][8] <= LLR_62;					inform_L [62][8] <= LLR_63;					inform_L [63][8] <= LLR_64;					inform_L [64][8] <= LLR_65;					inform_L [65][8] <= LLR_66;					inform_L [66][8] <= LLR_67;					inform_L [67][8] <= LLR_68;					inform_L [68][8] <= LLR_69;					inform_L [69][8] <= LLR_70;					inform_L [70][8] <= LLR_71;					inform_L [71][8] <= LLR_72;					inform_L [72][8] <= LLR_73;					inform_L [73][8] <= LLR_74;					inform_L [74][8] <= LLR_75;					inform_L [75][8] <= LLR_76;					inform_L [76][8] <= LLR_77;					inform_L [77][8] <= LLR_78;					inform_L [78][8] <= LLR_79;					inform_L [79][8] <= LLR_80;					inform_L [80][8] <= LLR_81;					inform_L [81][8] <= LLR_82;					inform_L [82][8] <= LLR_83;					inform_L [83][8] <= LLR_84;					inform_L [84][8] <= LLR_85;					inform_L [85][8] <= LLR_86;					inform_L [86][8] <= LLR_87;					inform_L [87][8] <= LLR_88;					inform_L [88][8] <= LLR_89;					inform_L [89][8] <= LLR_90;					inform_L [90][8] <= LLR_91;					inform_L [91][8] <= LLR_92;					inform_L [92][8] <= LLR_93;					inform_L [93][8] <= LLR_94;					inform_L [94][8] <= LLR_95;					inform_L [95][8] <= LLR_96;					inform_L [96][8] <= LLR_97;					inform_L [97][8] <= LLR_98;					inform_L [98][8] <= LLR_99;					inform_L [99][8] <= LLR_100;					inform_L [100][8] <= LLR_101;					inform_L [101][8] <= LLR_102;					inform_L [102][8] <= LLR_103;					inform_L [103][8] <= LLR_104;					inform_L [104][8] <= LLR_105;					inform_L [105][8] <= LLR_106;					inform_L [106][8] <= LLR_107;					inform_L [107][8] <= LLR_108;					inform_L [108][8] <= LLR_109;					inform_L [109][8] <= LLR_110;					inform_L [110][8] <= LLR_111;					inform_L [111][8] <= LLR_112;					inform_L [112][8] <= LLR_113;					inform_L [113][8] <= LLR_114;					inform_L [114][8] <= LLR_115;					inform_L [115][8] <= LLR_116;					inform_L [116][8] <= LLR_117;					inform_L [117][8] <= LLR_118;					inform_L [118][8] <= LLR_119;					inform_L [119][8] <= LLR_120;					inform_L [120][8] <= LLR_121;					inform_L [121][8] <= LLR_122;					inform_L [122][8] <= LLR_123;					inform_L [123][8] <= LLR_124;					inform_L [124][8] <= LLR_125;					inform_L [125][8] <= LLR_126;					inform_L [126][8] <= LLR_127;					inform_L [127][8] <= LLR_128;					inform_L [128][8] <= LLR_129;					inform_L [129][8] <= LLR_130;					inform_L [130][8] <= LLR_131;					inform_L [131][8] <= LLR_132;					inform_L [132][8] <= LLR_133;					inform_L [133][8] <= LLR_134;					inform_L [134][8] <= LLR_135;					inform_L [135][8] <= LLR_136;					inform_L [136][8] <= LLR_137;					inform_L [137][8] <= LLR_138;					inform_L [138][8] <= LLR_139;					inform_L [139][8] <= LLR_140;					inform_L [140][8] <= LLR_141;					inform_L [141][8] <= LLR_142;					inform_L [142][8] <= LLR_143;					inform_L [143][8] <= LLR_144;					inform_L [144][8] <= LLR_145;					inform_L [145][8] <= LLR_146;					inform_L [146][8] <= LLR_147;					inform_L [147][8] <= LLR_148;					inform_L [148][8] <= LLR_149;					inform_L [149][8] <= LLR_150;					inform_L [150][8] <= LLR_151;					inform_L [151][8] <= LLR_152;					inform_L [152][8] <= LLR_153;					inform_L [153][8] <= LLR_154;					inform_L [154][8] <= LLR_155;					inform_L [155][8] <= LLR_156;					inform_L [156][8] <= LLR_157;					inform_L [157][8] <= LLR_158;					inform_L [158][8] <= LLR_159;					inform_L [159][8] <= LLR_160;					inform_L [160][8] <= LLR_161;					inform_L [161][8] <= LLR_162;					inform_L [162][8] <= LLR_163;					inform_L [163][8] <= LLR_164;					inform_L [164][8] <= LLR_165;					inform_L [165][8] <= LLR_166;					inform_L [166][8] <= LLR_167;					inform_L [167][8] <= LLR_168;					inform_L [168][8] <= LLR_169;					inform_L [169][8] <= LLR_170;					inform_L [170][8] <= LLR_171;					inform_L [171][8] <= LLR_172;					inform_L [172][8] <= LLR_173;					inform_L [173][8] <= LLR_174;					inform_L [174][8] <= LLR_175;					inform_L [175][8] <= LLR_176;					inform_L [176][8] <= LLR_177;					inform_L [177][8] <= LLR_178;					inform_L [178][8] <= LLR_179;					inform_L [179][8] <= LLR_180;					inform_L [180][8] <= LLR_181;					inform_L [181][8] <= LLR_182;					inform_L [182][8] <= LLR_183;					inform_L [183][8] <= LLR_184;					inform_L [184][8] <= LLR_185;					inform_L [185][8] <= LLR_186;					inform_L [186][8] <= LLR_187;					inform_L [187][8] <= LLR_188;					inform_L [188][8] <= LLR_189;					inform_L [189][8] <= LLR_190;					inform_L [190][8] <= LLR_191;					inform_L [191][8] <= LLR_192;					inform_L [192][8] <= LLR_193;					inform_L [193][8] <= LLR_194;					inform_L [194][8] <= LLR_195;					inform_L [195][8] <= LLR_196;					inform_L [196][8] <= LLR_197;					inform_L [197][8] <= LLR_198;					inform_L [198][8] <= LLR_199;					inform_L [199][8] <= LLR_200;					inform_L [200][8] <= LLR_201;					inform_L [201][8] <= LLR_202;					inform_L [202][8] <= LLR_203;					inform_L [203][8] <= LLR_204;					inform_L [204][8] <= LLR_205;					inform_L [205][8] <= LLR_206;					inform_L [206][8] <= LLR_207;					inform_L [207][8] <= LLR_208;					inform_L [208][8] <= LLR_209;					inform_L [209][8] <= LLR_210;					inform_L [210][8] <= LLR_211;					inform_L [211][8] <= LLR_212;					inform_L [212][8] <= LLR_213;					inform_L [213][8] <= LLR_214;					inform_L [214][8] <= LLR_215;					inform_L [215][8] <= LLR_216;					inform_L [216][8] <= LLR_217;					inform_L [217][8] <= LLR_218;					inform_L [218][8] <= LLR_219;					inform_L [219][8] <= LLR_220;					inform_L [220][8] <= LLR_221;					inform_L [221][8] <= LLR_222;					inform_L [222][8] <= LLR_223;					inform_L [223][8] <= LLR_224;					inform_L [224][8] <= LLR_225;					inform_L [225][8] <= LLR_226;					inform_L [226][8] <= LLR_227;					inform_L [227][8] <= LLR_228;					inform_L [228][8] <= LLR_229;					inform_L [229][8] <= LLR_230;					inform_L [230][8] <= LLR_231;					inform_L [231][8] <= LLR_232;					inform_L [232][8] <= LLR_233;					inform_L [233][8] <= LLR_234;					inform_L [234][8] <= LLR_235;					inform_L [235][8] <= LLR_236;					inform_L [236][8] <= LLR_237;					inform_L [237][8] <= LLR_238;					inform_L [238][8] <= LLR_239;					inform_L [239][8] <= LLR_240;					inform_L [240][8] <= LLR_241;					inform_L [241][8] <= LLR_242;					inform_L [242][8] <= LLR_243;					inform_L [243][8] <= LLR_244;					inform_L [244][8] <= LLR_245;					inform_L [245][8] <= LLR_246;					inform_L [246][8] <= LLR_247;					inform_L [247][8] <= LLR_248;					inform_L [248][8] <= LLR_249;					inform_L [249][8] <= LLR_250;					inform_L [250][8] <= LLR_251;					inform_L [251][8] <= LLR_252;					inform_L [252][8] <= LLR_253;					inform_L [253][8] <= LLR_254;					inform_L [254][8] <= LLR_255;					inform_L [255][8] <= LLR_256;				end				for (x = 0; x < 256; x = x + 1)					for (y = 0; y < 8; y = y + 1)					begin						inform_R[x][y+1] <= 8'd0;						inform_L[x][y] <= 8'd0;					end			end
		endcase	end
	assign bp_over_flag = (itera_time == `iteration_times + 1) ? 1 : 0;
	always @(*)	begin		case (w2r)			1:			begin				r_cell_reg[0] = inform_R[0][0];				r_cell_reg[1] = inform_R[1][0];				r_cell_reg[2] = inform_R[2][0];				r_cell_reg[3] = inform_R[3][0];				r_cell_reg[4] = inform_R[4][0];				r_cell_reg[5] = inform_R[5][0];				r_cell_reg[6] = inform_R[6][0];				r_cell_reg[7] = inform_R[7][0];				r_cell_reg[8] = inform_R[8][0];				r_cell_reg[9] = inform_R[9][0];				r_cell_reg[10] = inform_R[10][0];				r_cell_reg[11] = inform_R[11][0];				r_cell_reg[12] = inform_R[12][0];				r_cell_reg[13] = inform_R[13][0];				r_cell_reg[14] = inform_R[14][0];				r_cell_reg[15] = inform_R[15][0];				r_cell_reg[16] = inform_R[16][0];				r_cell_reg[17] = inform_R[17][0];				r_cell_reg[18] = inform_R[18][0];				r_cell_reg[19] = inform_R[19][0];				r_cell_reg[20] = inform_R[20][0];				r_cell_reg[21] = inform_R[21][0];				r_cell_reg[22] = inform_R[22][0];				r_cell_reg[23] = inform_R[23][0];				r_cell_reg[24] = inform_R[24][0];				r_cell_reg[25] = inform_R[25][0];				r_cell_reg[26] = inform_R[26][0];				r_cell_reg[27] = inform_R[27][0];				r_cell_reg[28] = inform_R[28][0];				r_cell_reg[29] = inform_R[29][0];				r_cell_reg[30] = inform_R[30][0];				r_cell_reg[31] = inform_R[31][0];				r_cell_reg[32] = inform_R[32][0];				r_cell_reg[33] = inform_R[33][0];				r_cell_reg[34] = inform_R[34][0];				r_cell_reg[35] = inform_R[35][0];				r_cell_reg[36] = inform_R[36][0];				r_cell_reg[37] = inform_R[37][0];				r_cell_reg[38] = inform_R[38][0];				r_cell_reg[39] = inform_R[39][0];				r_cell_reg[40] = inform_R[40][0];				r_cell_reg[41] = inform_R[41][0];				r_cell_reg[42] = inform_R[42][0];				r_cell_reg[43] = inform_R[43][0];				r_cell_reg[44] = inform_R[44][0];				r_cell_reg[45] = inform_R[45][0];				r_cell_reg[46] = inform_R[46][0];				r_cell_reg[47] = inform_R[47][0];				r_cell_reg[48] = inform_R[48][0];				r_cell_reg[49] = inform_R[49][0];				r_cell_reg[50] = inform_R[50][0];				r_cell_reg[51] = inform_R[51][0];				r_cell_reg[52] = inform_R[52][0];				r_cell_reg[53] = inform_R[53][0];				r_cell_reg[54] = inform_R[54][0];				r_cell_reg[55] = inform_R[55][0];				r_cell_reg[56] = inform_R[56][0];				r_cell_reg[57] = inform_R[57][0];				r_cell_reg[58] = inform_R[58][0];				r_cell_reg[59] = inform_R[59][0];				r_cell_reg[60] = inform_R[60][0];				r_cell_reg[61] = inform_R[61][0];				r_cell_reg[62] = inform_R[62][0];				r_cell_reg[63] = inform_R[63][0];				r_cell_reg[64] = inform_R[64][0];				r_cell_reg[65] = inform_R[65][0];				r_cell_reg[66] = inform_R[66][0];				r_cell_reg[67] = inform_R[67][0];				r_cell_reg[68] = inform_R[68][0];				r_cell_reg[69] = inform_R[69][0];				r_cell_reg[70] = inform_R[70][0];				r_cell_reg[71] = inform_R[71][0];				r_cell_reg[72] = inform_R[72][0];				r_cell_reg[73] = inform_R[73][0];				r_cell_reg[74] = inform_R[74][0];				r_cell_reg[75] = inform_R[75][0];				r_cell_reg[76] = inform_R[76][0];				r_cell_reg[77] = inform_R[77][0];				r_cell_reg[78] = inform_R[78][0];				r_cell_reg[79] = inform_R[79][0];				r_cell_reg[80] = inform_R[80][0];				r_cell_reg[81] = inform_R[81][0];				r_cell_reg[82] = inform_R[82][0];				r_cell_reg[83] = inform_R[83][0];				r_cell_reg[84] = inform_R[84][0];				r_cell_reg[85] = inform_R[85][0];				r_cell_reg[86] = inform_R[86][0];				r_cell_reg[87] = inform_R[87][0];				r_cell_reg[88] = inform_R[88][0];				r_cell_reg[89] = inform_R[89][0];				r_cell_reg[90] = inform_R[90][0];				r_cell_reg[91] = inform_R[91][0];				r_cell_reg[92] = inform_R[92][0];				r_cell_reg[93] = inform_R[93][0];				r_cell_reg[94] = inform_R[94][0];				r_cell_reg[95] = inform_R[95][0];				r_cell_reg[96] = inform_R[96][0];				r_cell_reg[97] = inform_R[97][0];				r_cell_reg[98] = inform_R[98][0];				r_cell_reg[99] = inform_R[99][0];				r_cell_reg[100] = inform_R[100][0];				r_cell_reg[101] = inform_R[101][0];				r_cell_reg[102] = inform_R[102][0];				r_cell_reg[103] = inform_R[103][0];				r_cell_reg[104] = inform_R[104][0];				r_cell_reg[105] = inform_R[105][0];				r_cell_reg[106] = inform_R[106][0];				r_cell_reg[107] = inform_R[107][0];				r_cell_reg[108] = inform_R[108][0];				r_cell_reg[109] = inform_R[109][0];				r_cell_reg[110] = inform_R[110][0];				r_cell_reg[111] = inform_R[111][0];				r_cell_reg[112] = inform_R[112][0];				r_cell_reg[113] = inform_R[113][0];				r_cell_reg[114] = inform_R[114][0];				r_cell_reg[115] = inform_R[115][0];				r_cell_reg[116] = inform_R[116][0];				r_cell_reg[117] = inform_R[117][0];				r_cell_reg[118] = inform_R[118][0];				r_cell_reg[119] = inform_R[119][0];				r_cell_reg[120] = inform_R[120][0];				r_cell_reg[121] = inform_R[121][0];				r_cell_reg[122] = inform_R[122][0];				r_cell_reg[123] = inform_R[123][0];				r_cell_reg[124] = inform_R[124][0];				r_cell_reg[125] = inform_R[125][0];				r_cell_reg[126] = inform_R[126][0];				r_cell_reg[127] = inform_R[127][0];				r_cell_reg[128] = inform_R[128][0];				r_cell_reg[129] = inform_R[129][0];				r_cell_reg[130] = inform_R[130][0];				r_cell_reg[131] = inform_R[131][0];				r_cell_reg[132] = inform_R[132][0];				r_cell_reg[133] = inform_R[133][0];				r_cell_reg[134] = inform_R[134][0];				r_cell_reg[135] = inform_R[135][0];				r_cell_reg[136] = inform_R[136][0];				r_cell_reg[137] = inform_R[137][0];				r_cell_reg[138] = inform_R[138][0];				r_cell_reg[139] = inform_R[139][0];				r_cell_reg[140] = inform_R[140][0];				r_cell_reg[141] = inform_R[141][0];				r_cell_reg[142] = inform_R[142][0];				r_cell_reg[143] = inform_R[143][0];				r_cell_reg[144] = inform_R[144][0];				r_cell_reg[145] = inform_R[145][0];				r_cell_reg[146] = inform_R[146][0];				r_cell_reg[147] = inform_R[147][0];				r_cell_reg[148] = inform_R[148][0];				r_cell_reg[149] = inform_R[149][0];				r_cell_reg[150] = inform_R[150][0];				r_cell_reg[151] = inform_R[151][0];				r_cell_reg[152] = inform_R[152][0];				r_cell_reg[153] = inform_R[153][0];				r_cell_reg[154] = inform_R[154][0];				r_cell_reg[155] = inform_R[155][0];				r_cell_reg[156] = inform_R[156][0];				r_cell_reg[157] = inform_R[157][0];				r_cell_reg[158] = inform_R[158][0];				r_cell_reg[159] = inform_R[159][0];				r_cell_reg[160] = inform_R[160][0];				r_cell_reg[161] = inform_R[161][0];				r_cell_reg[162] = inform_R[162][0];				r_cell_reg[163] = inform_R[163][0];				r_cell_reg[164] = inform_R[164][0];				r_cell_reg[165] = inform_R[165][0];				r_cell_reg[166] = inform_R[166][0];				r_cell_reg[167] = inform_R[167][0];				r_cell_reg[168] = inform_R[168][0];				r_cell_reg[169] = inform_R[169][0];				r_cell_reg[170] = inform_R[170][0];				r_cell_reg[171] = inform_R[171][0];				r_cell_reg[172] = inform_R[172][0];				r_cell_reg[173] = inform_R[173][0];				r_cell_reg[174] = inform_R[174][0];				r_cell_reg[175] = inform_R[175][0];				r_cell_reg[176] = inform_R[176][0];				r_cell_reg[177] = inform_R[177][0];				r_cell_reg[178] = inform_R[178][0];				r_cell_reg[179] = inform_R[179][0];				r_cell_reg[180] = inform_R[180][0];				r_cell_reg[181] = inform_R[181][0];				r_cell_reg[182] = inform_R[182][0];				r_cell_reg[183] = inform_R[183][0];				r_cell_reg[184] = inform_R[184][0];				r_cell_reg[185] = inform_R[185][0];				r_cell_reg[186] = inform_R[186][0];				r_cell_reg[187] = inform_R[187][0];				r_cell_reg[188] = inform_R[188][0];				r_cell_reg[189] = inform_R[189][0];				r_cell_reg[190] = inform_R[190][0];				r_cell_reg[191] = inform_R[191][0];				r_cell_reg[192] = inform_R[192][0];				r_cell_reg[193] = inform_R[193][0];				r_cell_reg[194] = inform_R[194][0];				r_cell_reg[195] = inform_R[195][0];				r_cell_reg[196] = inform_R[196][0];				r_cell_reg[197] = inform_R[197][0];				r_cell_reg[198] = inform_R[198][0];				r_cell_reg[199] = inform_R[199][0];				r_cell_reg[200] = inform_R[200][0];				r_cell_reg[201] = inform_R[201][0];				r_cell_reg[202] = inform_R[202][0];				r_cell_reg[203] = inform_R[203][0];				r_cell_reg[204] = inform_R[204][0];				r_cell_reg[205] = inform_R[205][0];				r_cell_reg[206] = inform_R[206][0];				r_cell_reg[207] = inform_R[207][0];				r_cell_reg[208] = inform_R[208][0];				r_cell_reg[209] = inform_R[209][0];				r_cell_reg[210] = inform_R[210][0];				r_cell_reg[211] = inform_R[211][0];				r_cell_reg[212] = inform_R[212][0];				r_cell_reg[213] = inform_R[213][0];				r_cell_reg[214] = inform_R[214][0];				r_cell_reg[215] = inform_R[215][0];				r_cell_reg[216] = inform_R[216][0];				r_cell_reg[217] = inform_R[217][0];				r_cell_reg[218] = inform_R[218][0];				r_cell_reg[219] = inform_R[219][0];				r_cell_reg[220] = inform_R[220][0];				r_cell_reg[221] = inform_R[221][0];				r_cell_reg[222] = inform_R[222][0];				r_cell_reg[223] = inform_R[223][0];				r_cell_reg[224] = inform_R[224][0];				r_cell_reg[225] = inform_R[225][0];				r_cell_reg[226] = inform_R[226][0];				r_cell_reg[227] = inform_R[227][0];				r_cell_reg[228] = inform_R[228][0];				r_cell_reg[229] = inform_R[229][0];				r_cell_reg[230] = inform_R[230][0];				r_cell_reg[231] = inform_R[231][0];				r_cell_reg[232] = inform_R[232][0];				r_cell_reg[233] = inform_R[233][0];				r_cell_reg[234] = inform_R[234][0];				r_cell_reg[235] = inform_R[235][0];				r_cell_reg[236] = inform_R[236][0];				r_cell_reg[237] = inform_R[237][0];				r_cell_reg[238] = inform_R[238][0];				r_cell_reg[239] = inform_R[239][0];				r_cell_reg[240] = inform_R[240][0];				r_cell_reg[241] = inform_R[241][0];				r_cell_reg[242] = inform_R[242][0];				r_cell_reg[243] = inform_R[243][0];				r_cell_reg[244] = inform_R[244][0];				r_cell_reg[245] = inform_R[245][0];				r_cell_reg[246] = inform_R[246][0];				r_cell_reg[247] = inform_R[247][0];				r_cell_reg[248] = inform_R[248][0];				r_cell_reg[249] = inform_R[249][0];				r_cell_reg[250] = inform_R[250][0];				r_cell_reg[251] = inform_R[251][0];				r_cell_reg[252] = inform_R[252][0];				r_cell_reg[253] = inform_R[253][0];				r_cell_reg[254] = inform_R[254][0];				r_cell_reg[255] = inform_R[255][0];				l_cell_reg[0] = inform_L[0][1];				l_cell_reg[1] = inform_L[1][1];				l_cell_reg[2] = inform_L[2][1];				l_cell_reg[3] = inform_L[3][1];				l_cell_reg[4] = inform_L[4][1];				l_cell_reg[5] = inform_L[5][1];				l_cell_reg[6] = inform_L[6][1];				l_cell_reg[7] = inform_L[7][1];				l_cell_reg[8] = inform_L[8][1];				l_cell_reg[9] = inform_L[9][1];				l_cell_reg[10] = inform_L[10][1];				l_cell_reg[11] = inform_L[11][1];				l_cell_reg[12] = inform_L[12][1];				l_cell_reg[13] = inform_L[13][1];				l_cell_reg[14] = inform_L[14][1];				l_cell_reg[15] = inform_L[15][1];				l_cell_reg[16] = inform_L[16][1];				l_cell_reg[17] = inform_L[17][1];				l_cell_reg[18] = inform_L[18][1];				l_cell_reg[19] = inform_L[19][1];				l_cell_reg[20] = inform_L[20][1];				l_cell_reg[21] = inform_L[21][1];				l_cell_reg[22] = inform_L[22][1];				l_cell_reg[23] = inform_L[23][1];				l_cell_reg[24] = inform_L[24][1];				l_cell_reg[25] = inform_L[25][1];				l_cell_reg[26] = inform_L[26][1];				l_cell_reg[27] = inform_L[27][1];				l_cell_reg[28] = inform_L[28][1];				l_cell_reg[29] = inform_L[29][1];				l_cell_reg[30] = inform_L[30][1];				l_cell_reg[31] = inform_L[31][1];				l_cell_reg[32] = inform_L[32][1];				l_cell_reg[33] = inform_L[33][1];				l_cell_reg[34] = inform_L[34][1];				l_cell_reg[35] = inform_L[35][1];				l_cell_reg[36] = inform_L[36][1];				l_cell_reg[37] = inform_L[37][1];				l_cell_reg[38] = inform_L[38][1];				l_cell_reg[39] = inform_L[39][1];				l_cell_reg[40] = inform_L[40][1];				l_cell_reg[41] = inform_L[41][1];				l_cell_reg[42] = inform_L[42][1];				l_cell_reg[43] = inform_L[43][1];				l_cell_reg[44] = inform_L[44][1];				l_cell_reg[45] = inform_L[45][1];				l_cell_reg[46] = inform_L[46][1];				l_cell_reg[47] = inform_L[47][1];				l_cell_reg[48] = inform_L[48][1];				l_cell_reg[49] = inform_L[49][1];				l_cell_reg[50] = inform_L[50][1];				l_cell_reg[51] = inform_L[51][1];				l_cell_reg[52] = inform_L[52][1];				l_cell_reg[53] = inform_L[53][1];				l_cell_reg[54] = inform_L[54][1];				l_cell_reg[55] = inform_L[55][1];				l_cell_reg[56] = inform_L[56][1];				l_cell_reg[57] = inform_L[57][1];				l_cell_reg[58] = inform_L[58][1];				l_cell_reg[59] = inform_L[59][1];				l_cell_reg[60] = inform_L[60][1];				l_cell_reg[61] = inform_L[61][1];				l_cell_reg[62] = inform_L[62][1];				l_cell_reg[63] = inform_L[63][1];				l_cell_reg[64] = inform_L[64][1];				l_cell_reg[65] = inform_L[65][1];				l_cell_reg[66] = inform_L[66][1];				l_cell_reg[67] = inform_L[67][1];				l_cell_reg[68] = inform_L[68][1];				l_cell_reg[69] = inform_L[69][1];				l_cell_reg[70] = inform_L[70][1];				l_cell_reg[71] = inform_L[71][1];				l_cell_reg[72] = inform_L[72][1];				l_cell_reg[73] = inform_L[73][1];				l_cell_reg[74] = inform_L[74][1];				l_cell_reg[75] = inform_L[75][1];				l_cell_reg[76] = inform_L[76][1];				l_cell_reg[77] = inform_L[77][1];				l_cell_reg[78] = inform_L[78][1];				l_cell_reg[79] = inform_L[79][1];				l_cell_reg[80] = inform_L[80][1];				l_cell_reg[81] = inform_L[81][1];				l_cell_reg[82] = inform_L[82][1];				l_cell_reg[83] = inform_L[83][1];				l_cell_reg[84] = inform_L[84][1];				l_cell_reg[85] = inform_L[85][1];				l_cell_reg[86] = inform_L[86][1];				l_cell_reg[87] = inform_L[87][1];				l_cell_reg[88] = inform_L[88][1];				l_cell_reg[89] = inform_L[89][1];				l_cell_reg[90] = inform_L[90][1];				l_cell_reg[91] = inform_L[91][1];				l_cell_reg[92] = inform_L[92][1];				l_cell_reg[93] = inform_L[93][1];				l_cell_reg[94] = inform_L[94][1];				l_cell_reg[95] = inform_L[95][1];				l_cell_reg[96] = inform_L[96][1];				l_cell_reg[97] = inform_L[97][1];				l_cell_reg[98] = inform_L[98][1];				l_cell_reg[99] = inform_L[99][1];				l_cell_reg[100] = inform_L[100][1];				l_cell_reg[101] = inform_L[101][1];				l_cell_reg[102] = inform_L[102][1];				l_cell_reg[103] = inform_L[103][1];				l_cell_reg[104] = inform_L[104][1];				l_cell_reg[105] = inform_L[105][1];				l_cell_reg[106] = inform_L[106][1];				l_cell_reg[107] = inform_L[107][1];				l_cell_reg[108] = inform_L[108][1];				l_cell_reg[109] = inform_L[109][1];				l_cell_reg[110] = inform_L[110][1];				l_cell_reg[111] = inform_L[111][1];				l_cell_reg[112] = inform_L[112][1];				l_cell_reg[113] = inform_L[113][1];				l_cell_reg[114] = inform_L[114][1];				l_cell_reg[115] = inform_L[115][1];				l_cell_reg[116] = inform_L[116][1];				l_cell_reg[117] = inform_L[117][1];				l_cell_reg[118] = inform_L[118][1];				l_cell_reg[119] = inform_L[119][1];				l_cell_reg[120] = inform_L[120][1];				l_cell_reg[121] = inform_L[121][1];				l_cell_reg[122] = inform_L[122][1];				l_cell_reg[123] = inform_L[123][1];				l_cell_reg[124] = inform_L[124][1];				l_cell_reg[125] = inform_L[125][1];				l_cell_reg[126] = inform_L[126][1];				l_cell_reg[127] = inform_L[127][1];				l_cell_reg[128] = inform_L[128][1];				l_cell_reg[129] = inform_L[129][1];				l_cell_reg[130] = inform_L[130][1];				l_cell_reg[131] = inform_L[131][1];				l_cell_reg[132] = inform_L[132][1];				l_cell_reg[133] = inform_L[133][1];				l_cell_reg[134] = inform_L[134][1];				l_cell_reg[135] = inform_L[135][1];				l_cell_reg[136] = inform_L[136][1];				l_cell_reg[137] = inform_L[137][1];				l_cell_reg[138] = inform_L[138][1];				l_cell_reg[139] = inform_L[139][1];				l_cell_reg[140] = inform_L[140][1];				l_cell_reg[141] = inform_L[141][1];				l_cell_reg[142] = inform_L[142][1];				l_cell_reg[143] = inform_L[143][1];				l_cell_reg[144] = inform_L[144][1];				l_cell_reg[145] = inform_L[145][1];				l_cell_reg[146] = inform_L[146][1];				l_cell_reg[147] = inform_L[147][1];				l_cell_reg[148] = inform_L[148][1];				l_cell_reg[149] = inform_L[149][1];				l_cell_reg[150] = inform_L[150][1];				l_cell_reg[151] = inform_L[151][1];				l_cell_reg[152] = inform_L[152][1];				l_cell_reg[153] = inform_L[153][1];				l_cell_reg[154] = inform_L[154][1];				l_cell_reg[155] = inform_L[155][1];				l_cell_reg[156] = inform_L[156][1];				l_cell_reg[157] = inform_L[157][1];				l_cell_reg[158] = inform_L[158][1];				l_cell_reg[159] = inform_L[159][1];				l_cell_reg[160] = inform_L[160][1];				l_cell_reg[161] = inform_L[161][1];				l_cell_reg[162] = inform_L[162][1];				l_cell_reg[163] = inform_L[163][1];				l_cell_reg[164] = inform_L[164][1];				l_cell_reg[165] = inform_L[165][1];				l_cell_reg[166] = inform_L[166][1];				l_cell_reg[167] = inform_L[167][1];				l_cell_reg[168] = inform_L[168][1];				l_cell_reg[169] = inform_L[169][1];				l_cell_reg[170] = inform_L[170][1];				l_cell_reg[171] = inform_L[171][1];				l_cell_reg[172] = inform_L[172][1];				l_cell_reg[173] = inform_L[173][1];				l_cell_reg[174] = inform_L[174][1];				l_cell_reg[175] = inform_L[175][1];				l_cell_reg[176] = inform_L[176][1];				l_cell_reg[177] = inform_L[177][1];				l_cell_reg[178] = inform_L[178][1];				l_cell_reg[179] = inform_L[179][1];				l_cell_reg[180] = inform_L[180][1];				l_cell_reg[181] = inform_L[181][1];				l_cell_reg[182] = inform_L[182][1];				l_cell_reg[183] = inform_L[183][1];				l_cell_reg[184] = inform_L[184][1];				l_cell_reg[185] = inform_L[185][1];				l_cell_reg[186] = inform_L[186][1];				l_cell_reg[187] = inform_L[187][1];				l_cell_reg[188] = inform_L[188][1];				l_cell_reg[189] = inform_L[189][1];				l_cell_reg[190] = inform_L[190][1];				l_cell_reg[191] = inform_L[191][1];				l_cell_reg[192] = inform_L[192][1];				l_cell_reg[193] = inform_L[193][1];				l_cell_reg[194] = inform_L[194][1];				l_cell_reg[195] = inform_L[195][1];				l_cell_reg[196] = inform_L[196][1];				l_cell_reg[197] = inform_L[197][1];				l_cell_reg[198] = inform_L[198][1];				l_cell_reg[199] = inform_L[199][1];				l_cell_reg[200] = inform_L[200][1];				l_cell_reg[201] = inform_L[201][1];				l_cell_reg[202] = inform_L[202][1];				l_cell_reg[203] = inform_L[203][1];				l_cell_reg[204] = inform_L[204][1];				l_cell_reg[205] = inform_L[205][1];				l_cell_reg[206] = inform_L[206][1];				l_cell_reg[207] = inform_L[207][1];				l_cell_reg[208] = inform_L[208][1];				l_cell_reg[209] = inform_L[209][1];				l_cell_reg[210] = inform_L[210][1];				l_cell_reg[211] = inform_L[211][1];				l_cell_reg[212] = inform_L[212][1];				l_cell_reg[213] = inform_L[213][1];				l_cell_reg[214] = inform_L[214][1];				l_cell_reg[215] = inform_L[215][1];				l_cell_reg[216] = inform_L[216][1];				l_cell_reg[217] = inform_L[217][1];				l_cell_reg[218] = inform_L[218][1];				l_cell_reg[219] = inform_L[219][1];				l_cell_reg[220] = inform_L[220][1];				l_cell_reg[221] = inform_L[221][1];				l_cell_reg[222] = inform_L[222][1];				l_cell_reg[223] = inform_L[223][1];				l_cell_reg[224] = inform_L[224][1];				l_cell_reg[225] = inform_L[225][1];				l_cell_reg[226] = inform_L[226][1];				l_cell_reg[227] = inform_L[227][1];				l_cell_reg[228] = inform_L[228][1];				l_cell_reg[229] = inform_L[229][1];				l_cell_reg[230] = inform_L[230][1];				l_cell_reg[231] = inform_L[231][1];				l_cell_reg[232] = inform_L[232][1];				l_cell_reg[233] = inform_L[233][1];				l_cell_reg[234] = inform_L[234][1];				l_cell_reg[235] = inform_L[235][1];				l_cell_reg[236] = inform_L[236][1];				l_cell_reg[237] = inform_L[237][1];				l_cell_reg[238] = inform_L[238][1];				l_cell_reg[239] = inform_L[239][1];				l_cell_reg[240] = inform_L[240][1];				l_cell_reg[241] = inform_L[241][1];				l_cell_reg[242] = inform_L[242][1];				l_cell_reg[243] = inform_L[243][1];				l_cell_reg[244] = inform_L[244][1];				l_cell_reg[245] = inform_L[245][1];				l_cell_reg[246] = inform_L[246][1];				l_cell_reg[247] = inform_L[247][1];				l_cell_reg[248] = inform_L[248][1];				l_cell_reg[249] = inform_L[249][1];				l_cell_reg[250] = inform_L[250][1];				l_cell_reg[251] = inform_L[251][1];				l_cell_reg[252] = inform_L[252][1];				l_cell_reg[253] = inform_L[253][1];				l_cell_reg[254] = inform_L[254][1];				l_cell_reg[255] = inform_L[255][1];			end
			2:			begin				r_cell_reg[0] = inform_R[0][1];				r_cell_reg[1] = inform_R[2][1];				r_cell_reg[2] = inform_R[1][1];				r_cell_reg[3] = inform_R[3][1];				r_cell_reg[4] = inform_R[4][1];				r_cell_reg[5] = inform_R[6][1];				r_cell_reg[6] = inform_R[5][1];				r_cell_reg[7] = inform_R[7][1];				r_cell_reg[8] = inform_R[8][1];				r_cell_reg[9] = inform_R[10][1];				r_cell_reg[10] = inform_R[9][1];				r_cell_reg[11] = inform_R[11][1];				r_cell_reg[12] = inform_R[12][1];				r_cell_reg[13] = inform_R[14][1];				r_cell_reg[14] = inform_R[13][1];				r_cell_reg[15] = inform_R[15][1];				r_cell_reg[16] = inform_R[16][1];				r_cell_reg[17] = inform_R[18][1];				r_cell_reg[18] = inform_R[17][1];				r_cell_reg[19] = inform_R[19][1];				r_cell_reg[20] = inform_R[20][1];				r_cell_reg[21] = inform_R[22][1];				r_cell_reg[22] = inform_R[21][1];				r_cell_reg[23] = inform_R[23][1];				r_cell_reg[24] = inform_R[24][1];				r_cell_reg[25] = inform_R[26][1];				r_cell_reg[26] = inform_R[25][1];				r_cell_reg[27] = inform_R[27][1];				r_cell_reg[28] = inform_R[28][1];				r_cell_reg[29] = inform_R[30][1];				r_cell_reg[30] = inform_R[29][1];				r_cell_reg[31] = inform_R[31][1];				r_cell_reg[32] = inform_R[32][1];				r_cell_reg[33] = inform_R[34][1];				r_cell_reg[34] = inform_R[33][1];				r_cell_reg[35] = inform_R[35][1];				r_cell_reg[36] = inform_R[36][1];				r_cell_reg[37] = inform_R[38][1];				r_cell_reg[38] = inform_R[37][1];				r_cell_reg[39] = inform_R[39][1];				r_cell_reg[40] = inform_R[40][1];				r_cell_reg[41] = inform_R[42][1];				r_cell_reg[42] = inform_R[41][1];				r_cell_reg[43] = inform_R[43][1];				r_cell_reg[44] = inform_R[44][1];				r_cell_reg[45] = inform_R[46][1];				r_cell_reg[46] = inform_R[45][1];				r_cell_reg[47] = inform_R[47][1];				r_cell_reg[48] = inform_R[48][1];				r_cell_reg[49] = inform_R[50][1];				r_cell_reg[50] = inform_R[49][1];				r_cell_reg[51] = inform_R[51][1];				r_cell_reg[52] = inform_R[52][1];				r_cell_reg[53] = inform_R[54][1];				r_cell_reg[54] = inform_R[53][1];				r_cell_reg[55] = inform_R[55][1];				r_cell_reg[56] = inform_R[56][1];				r_cell_reg[57] = inform_R[58][1];				r_cell_reg[58] = inform_R[57][1];				r_cell_reg[59] = inform_R[59][1];				r_cell_reg[60] = inform_R[60][1];				r_cell_reg[61] = inform_R[62][1];				r_cell_reg[62] = inform_R[61][1];				r_cell_reg[63] = inform_R[63][1];				r_cell_reg[64] = inform_R[64][1];				r_cell_reg[65] = inform_R[66][1];				r_cell_reg[66] = inform_R[65][1];				r_cell_reg[67] = inform_R[67][1];				r_cell_reg[68] = inform_R[68][1];				r_cell_reg[69] = inform_R[70][1];				r_cell_reg[70] = inform_R[69][1];				r_cell_reg[71] = inform_R[71][1];				r_cell_reg[72] = inform_R[72][1];				r_cell_reg[73] = inform_R[74][1];				r_cell_reg[74] = inform_R[73][1];				r_cell_reg[75] = inform_R[75][1];				r_cell_reg[76] = inform_R[76][1];				r_cell_reg[77] = inform_R[78][1];				r_cell_reg[78] = inform_R[77][1];				r_cell_reg[79] = inform_R[79][1];				r_cell_reg[80] = inform_R[80][1];				r_cell_reg[81] = inform_R[82][1];				r_cell_reg[82] = inform_R[81][1];				r_cell_reg[83] = inform_R[83][1];				r_cell_reg[84] = inform_R[84][1];				r_cell_reg[85] = inform_R[86][1];				r_cell_reg[86] = inform_R[85][1];				r_cell_reg[87] = inform_R[87][1];				r_cell_reg[88] = inform_R[88][1];				r_cell_reg[89] = inform_R[90][1];				r_cell_reg[90] = inform_R[89][1];				r_cell_reg[91] = inform_R[91][1];				r_cell_reg[92] = inform_R[92][1];				r_cell_reg[93] = inform_R[94][1];				r_cell_reg[94] = inform_R[93][1];				r_cell_reg[95] = inform_R[95][1];				r_cell_reg[96] = inform_R[96][1];				r_cell_reg[97] = inform_R[98][1];				r_cell_reg[98] = inform_R[97][1];				r_cell_reg[99] = inform_R[99][1];				r_cell_reg[100] = inform_R[100][1];				r_cell_reg[101] = inform_R[102][1];				r_cell_reg[102] = inform_R[101][1];				r_cell_reg[103] = inform_R[103][1];				r_cell_reg[104] = inform_R[104][1];				r_cell_reg[105] = inform_R[106][1];				r_cell_reg[106] = inform_R[105][1];				r_cell_reg[107] = inform_R[107][1];				r_cell_reg[108] = inform_R[108][1];				r_cell_reg[109] = inform_R[110][1];				r_cell_reg[110] = inform_R[109][1];				r_cell_reg[111] = inform_R[111][1];				r_cell_reg[112] = inform_R[112][1];				r_cell_reg[113] = inform_R[114][1];				r_cell_reg[114] = inform_R[113][1];				r_cell_reg[115] = inform_R[115][1];				r_cell_reg[116] = inform_R[116][1];				r_cell_reg[117] = inform_R[118][1];				r_cell_reg[118] = inform_R[117][1];				r_cell_reg[119] = inform_R[119][1];				r_cell_reg[120] = inform_R[120][1];				r_cell_reg[121] = inform_R[122][1];				r_cell_reg[122] = inform_R[121][1];				r_cell_reg[123] = inform_R[123][1];				r_cell_reg[124] = inform_R[124][1];				r_cell_reg[125] = inform_R[126][1];				r_cell_reg[126] = inform_R[125][1];				r_cell_reg[127] = inform_R[127][1];				r_cell_reg[128] = inform_R[128][1];				r_cell_reg[129] = inform_R[130][1];				r_cell_reg[130] = inform_R[129][1];				r_cell_reg[131] = inform_R[131][1];				r_cell_reg[132] = inform_R[132][1];				r_cell_reg[133] = inform_R[134][1];				r_cell_reg[134] = inform_R[133][1];				r_cell_reg[135] = inform_R[135][1];				r_cell_reg[136] = inform_R[136][1];				r_cell_reg[137] = inform_R[138][1];				r_cell_reg[138] = inform_R[137][1];				r_cell_reg[139] = inform_R[139][1];				r_cell_reg[140] = inform_R[140][1];				r_cell_reg[141] = inform_R[142][1];				r_cell_reg[142] = inform_R[141][1];				r_cell_reg[143] = inform_R[143][1];				r_cell_reg[144] = inform_R[144][1];				r_cell_reg[145] = inform_R[146][1];				r_cell_reg[146] = inform_R[145][1];				r_cell_reg[147] = inform_R[147][1];				r_cell_reg[148] = inform_R[148][1];				r_cell_reg[149] = inform_R[150][1];				r_cell_reg[150] = inform_R[149][1];				r_cell_reg[151] = inform_R[151][1];				r_cell_reg[152] = inform_R[152][1];				r_cell_reg[153] = inform_R[154][1];				r_cell_reg[154] = inform_R[153][1];				r_cell_reg[155] = inform_R[155][1];				r_cell_reg[156] = inform_R[156][1];				r_cell_reg[157] = inform_R[158][1];				r_cell_reg[158] = inform_R[157][1];				r_cell_reg[159] = inform_R[159][1];				r_cell_reg[160] = inform_R[160][1];				r_cell_reg[161] = inform_R[162][1];				r_cell_reg[162] = inform_R[161][1];				r_cell_reg[163] = inform_R[163][1];				r_cell_reg[164] = inform_R[164][1];				r_cell_reg[165] = inform_R[166][1];				r_cell_reg[166] = inform_R[165][1];				r_cell_reg[167] = inform_R[167][1];				r_cell_reg[168] = inform_R[168][1];				r_cell_reg[169] = inform_R[170][1];				r_cell_reg[170] = inform_R[169][1];				r_cell_reg[171] = inform_R[171][1];				r_cell_reg[172] = inform_R[172][1];				r_cell_reg[173] = inform_R[174][1];				r_cell_reg[174] = inform_R[173][1];				r_cell_reg[175] = inform_R[175][1];				r_cell_reg[176] = inform_R[176][1];				r_cell_reg[177] = inform_R[178][1];				r_cell_reg[178] = inform_R[177][1];				r_cell_reg[179] = inform_R[179][1];				r_cell_reg[180] = inform_R[180][1];				r_cell_reg[181] = inform_R[182][1];				r_cell_reg[182] = inform_R[181][1];				r_cell_reg[183] = inform_R[183][1];				r_cell_reg[184] = inform_R[184][1];				r_cell_reg[185] = inform_R[186][1];				r_cell_reg[186] = inform_R[185][1];				r_cell_reg[187] = inform_R[187][1];				r_cell_reg[188] = inform_R[188][1];				r_cell_reg[189] = inform_R[190][1];				r_cell_reg[190] = inform_R[189][1];				r_cell_reg[191] = inform_R[191][1];				r_cell_reg[192] = inform_R[192][1];				r_cell_reg[193] = inform_R[194][1];				r_cell_reg[194] = inform_R[193][1];				r_cell_reg[195] = inform_R[195][1];				r_cell_reg[196] = inform_R[196][1];				r_cell_reg[197] = inform_R[198][1];				r_cell_reg[198] = inform_R[197][1];				r_cell_reg[199] = inform_R[199][1];				r_cell_reg[200] = inform_R[200][1];				r_cell_reg[201] = inform_R[202][1];				r_cell_reg[202] = inform_R[201][1];				r_cell_reg[203] = inform_R[203][1];				r_cell_reg[204] = inform_R[204][1];				r_cell_reg[205] = inform_R[206][1];				r_cell_reg[206] = inform_R[205][1];				r_cell_reg[207] = inform_R[207][1];				r_cell_reg[208] = inform_R[208][1];				r_cell_reg[209] = inform_R[210][1];				r_cell_reg[210] = inform_R[209][1];				r_cell_reg[211] = inform_R[211][1];				r_cell_reg[212] = inform_R[212][1];				r_cell_reg[213] = inform_R[214][1];				r_cell_reg[214] = inform_R[213][1];				r_cell_reg[215] = inform_R[215][1];				r_cell_reg[216] = inform_R[216][1];				r_cell_reg[217] = inform_R[218][1];				r_cell_reg[218] = inform_R[217][1];				r_cell_reg[219] = inform_R[219][1];				r_cell_reg[220] = inform_R[220][1];				r_cell_reg[221] = inform_R[222][1];				r_cell_reg[222] = inform_R[221][1];				r_cell_reg[223] = inform_R[223][1];				r_cell_reg[224] = inform_R[224][1];				r_cell_reg[225] = inform_R[226][1];				r_cell_reg[226] = inform_R[225][1];				r_cell_reg[227] = inform_R[227][1];				r_cell_reg[228] = inform_R[228][1];				r_cell_reg[229] = inform_R[230][1];				r_cell_reg[230] = inform_R[229][1];				r_cell_reg[231] = inform_R[231][1];				r_cell_reg[232] = inform_R[232][1];				r_cell_reg[233] = inform_R[234][1];				r_cell_reg[234] = inform_R[233][1];				r_cell_reg[235] = inform_R[235][1];				r_cell_reg[236] = inform_R[236][1];				r_cell_reg[237] = inform_R[238][1];				r_cell_reg[238] = inform_R[237][1];				r_cell_reg[239] = inform_R[239][1];				r_cell_reg[240] = inform_R[240][1];				r_cell_reg[241] = inform_R[242][1];				r_cell_reg[242] = inform_R[241][1];				r_cell_reg[243] = inform_R[243][1];				r_cell_reg[244] = inform_R[244][1];				r_cell_reg[245] = inform_R[246][1];				r_cell_reg[246] = inform_R[245][1];				r_cell_reg[247] = inform_R[247][1];				r_cell_reg[248] = inform_R[248][1];				r_cell_reg[249] = inform_R[250][1];				r_cell_reg[250] = inform_R[249][1];				r_cell_reg[251] = inform_R[251][1];				r_cell_reg[252] = inform_R[252][1];				r_cell_reg[253] = inform_R[254][1];				r_cell_reg[254] = inform_R[253][1];				r_cell_reg[255] = inform_R[255][1];				l_cell_reg[0] = inform_L[0][2];				l_cell_reg[1] = inform_L[2][2];				l_cell_reg[2] = inform_L[1][2];				l_cell_reg[3] = inform_L[3][2];				l_cell_reg[4] = inform_L[4][2];				l_cell_reg[5] = inform_L[6][2];				l_cell_reg[6] = inform_L[5][2];				l_cell_reg[7] = inform_L[7][2];				l_cell_reg[8] = inform_L[8][2];				l_cell_reg[9] = inform_L[10][2];				l_cell_reg[10] = inform_L[9][2];				l_cell_reg[11] = inform_L[11][2];				l_cell_reg[12] = inform_L[12][2];				l_cell_reg[13] = inform_L[14][2];				l_cell_reg[14] = inform_L[13][2];				l_cell_reg[15] = inform_L[15][2];				l_cell_reg[16] = inform_L[16][2];				l_cell_reg[17] = inform_L[18][2];				l_cell_reg[18] = inform_L[17][2];				l_cell_reg[19] = inform_L[19][2];				l_cell_reg[20] = inform_L[20][2];				l_cell_reg[21] = inform_L[22][2];				l_cell_reg[22] = inform_L[21][2];				l_cell_reg[23] = inform_L[23][2];				l_cell_reg[24] = inform_L[24][2];				l_cell_reg[25] = inform_L[26][2];				l_cell_reg[26] = inform_L[25][2];				l_cell_reg[27] = inform_L[27][2];				l_cell_reg[28] = inform_L[28][2];				l_cell_reg[29] = inform_L[30][2];				l_cell_reg[30] = inform_L[29][2];				l_cell_reg[31] = inform_L[31][2];				l_cell_reg[32] = inform_L[32][2];				l_cell_reg[33] = inform_L[34][2];				l_cell_reg[34] = inform_L[33][2];				l_cell_reg[35] = inform_L[35][2];				l_cell_reg[36] = inform_L[36][2];				l_cell_reg[37] = inform_L[38][2];				l_cell_reg[38] = inform_L[37][2];				l_cell_reg[39] = inform_L[39][2];				l_cell_reg[40] = inform_L[40][2];				l_cell_reg[41] = inform_L[42][2];				l_cell_reg[42] = inform_L[41][2];				l_cell_reg[43] = inform_L[43][2];				l_cell_reg[44] = inform_L[44][2];				l_cell_reg[45] = inform_L[46][2];				l_cell_reg[46] = inform_L[45][2];				l_cell_reg[47] = inform_L[47][2];				l_cell_reg[48] = inform_L[48][2];				l_cell_reg[49] = inform_L[50][2];				l_cell_reg[50] = inform_L[49][2];				l_cell_reg[51] = inform_L[51][2];				l_cell_reg[52] = inform_L[52][2];				l_cell_reg[53] = inform_L[54][2];				l_cell_reg[54] = inform_L[53][2];				l_cell_reg[55] = inform_L[55][2];				l_cell_reg[56] = inform_L[56][2];				l_cell_reg[57] = inform_L[58][2];				l_cell_reg[58] = inform_L[57][2];				l_cell_reg[59] = inform_L[59][2];				l_cell_reg[60] = inform_L[60][2];				l_cell_reg[61] = inform_L[62][2];				l_cell_reg[62] = inform_L[61][2];				l_cell_reg[63] = inform_L[63][2];				l_cell_reg[64] = inform_L[64][2];				l_cell_reg[65] = inform_L[66][2];				l_cell_reg[66] = inform_L[65][2];				l_cell_reg[67] = inform_L[67][2];				l_cell_reg[68] = inform_L[68][2];				l_cell_reg[69] = inform_L[70][2];				l_cell_reg[70] = inform_L[69][2];				l_cell_reg[71] = inform_L[71][2];				l_cell_reg[72] = inform_L[72][2];				l_cell_reg[73] = inform_L[74][2];				l_cell_reg[74] = inform_L[73][2];				l_cell_reg[75] = inform_L[75][2];				l_cell_reg[76] = inform_L[76][2];				l_cell_reg[77] = inform_L[78][2];				l_cell_reg[78] = inform_L[77][2];				l_cell_reg[79] = inform_L[79][2];				l_cell_reg[80] = inform_L[80][2];				l_cell_reg[81] = inform_L[82][2];				l_cell_reg[82] = inform_L[81][2];				l_cell_reg[83] = inform_L[83][2];				l_cell_reg[84] = inform_L[84][2];				l_cell_reg[85] = inform_L[86][2];				l_cell_reg[86] = inform_L[85][2];				l_cell_reg[87] = inform_L[87][2];				l_cell_reg[88] = inform_L[88][2];				l_cell_reg[89] = inform_L[90][2];				l_cell_reg[90] = inform_L[89][2];				l_cell_reg[91] = inform_L[91][2];				l_cell_reg[92] = inform_L[92][2];				l_cell_reg[93] = inform_L[94][2];				l_cell_reg[94] = inform_L[93][2];				l_cell_reg[95] = inform_L[95][2];				l_cell_reg[96] = inform_L[96][2];				l_cell_reg[97] = inform_L[98][2];				l_cell_reg[98] = inform_L[97][2];				l_cell_reg[99] = inform_L[99][2];				l_cell_reg[100] = inform_L[100][2];				l_cell_reg[101] = inform_L[102][2];				l_cell_reg[102] = inform_L[101][2];				l_cell_reg[103] = inform_L[103][2];				l_cell_reg[104] = inform_L[104][2];				l_cell_reg[105] = inform_L[106][2];				l_cell_reg[106] = inform_L[105][2];				l_cell_reg[107] = inform_L[107][2];				l_cell_reg[108] = inform_L[108][2];				l_cell_reg[109] = inform_L[110][2];				l_cell_reg[110] = inform_L[109][2];				l_cell_reg[111] = inform_L[111][2];				l_cell_reg[112] = inform_L[112][2];				l_cell_reg[113] = inform_L[114][2];				l_cell_reg[114] = inform_L[113][2];				l_cell_reg[115] = inform_L[115][2];				l_cell_reg[116] = inform_L[116][2];				l_cell_reg[117] = inform_L[118][2];				l_cell_reg[118] = inform_L[117][2];				l_cell_reg[119] = inform_L[119][2];				l_cell_reg[120] = inform_L[120][2];				l_cell_reg[121] = inform_L[122][2];				l_cell_reg[122] = inform_L[121][2];				l_cell_reg[123] = inform_L[123][2];				l_cell_reg[124] = inform_L[124][2];				l_cell_reg[125] = inform_L[126][2];				l_cell_reg[126] = inform_L[125][2];				l_cell_reg[127] = inform_L[127][2];				l_cell_reg[128] = inform_L[128][2];				l_cell_reg[129] = inform_L[130][2];				l_cell_reg[130] = inform_L[129][2];				l_cell_reg[131] = inform_L[131][2];				l_cell_reg[132] = inform_L[132][2];				l_cell_reg[133] = inform_L[134][2];				l_cell_reg[134] = inform_L[133][2];				l_cell_reg[135] = inform_L[135][2];				l_cell_reg[136] = inform_L[136][2];				l_cell_reg[137] = inform_L[138][2];				l_cell_reg[138] = inform_L[137][2];				l_cell_reg[139] = inform_L[139][2];				l_cell_reg[140] = inform_L[140][2];				l_cell_reg[141] = inform_L[142][2];				l_cell_reg[142] = inform_L[141][2];				l_cell_reg[143] = inform_L[143][2];				l_cell_reg[144] = inform_L[144][2];				l_cell_reg[145] = inform_L[146][2];				l_cell_reg[146] = inform_L[145][2];				l_cell_reg[147] = inform_L[147][2];				l_cell_reg[148] = inform_L[148][2];				l_cell_reg[149] = inform_L[150][2];				l_cell_reg[150] = inform_L[149][2];				l_cell_reg[151] = inform_L[151][2];				l_cell_reg[152] = inform_L[152][2];				l_cell_reg[153] = inform_L[154][2];				l_cell_reg[154] = inform_L[153][2];				l_cell_reg[155] = inform_L[155][2];				l_cell_reg[156] = inform_L[156][2];				l_cell_reg[157] = inform_L[158][2];				l_cell_reg[158] = inform_L[157][2];				l_cell_reg[159] = inform_L[159][2];				l_cell_reg[160] = inform_L[160][2];				l_cell_reg[161] = inform_L[162][2];				l_cell_reg[162] = inform_L[161][2];				l_cell_reg[163] = inform_L[163][2];				l_cell_reg[164] = inform_L[164][2];				l_cell_reg[165] = inform_L[166][2];				l_cell_reg[166] = inform_L[165][2];				l_cell_reg[167] = inform_L[167][2];				l_cell_reg[168] = inform_L[168][2];				l_cell_reg[169] = inform_L[170][2];				l_cell_reg[170] = inform_L[169][2];				l_cell_reg[171] = inform_L[171][2];				l_cell_reg[172] = inform_L[172][2];				l_cell_reg[173] = inform_L[174][2];				l_cell_reg[174] = inform_L[173][2];				l_cell_reg[175] = inform_L[175][2];				l_cell_reg[176] = inform_L[176][2];				l_cell_reg[177] = inform_L[178][2];				l_cell_reg[178] = inform_L[177][2];				l_cell_reg[179] = inform_L[179][2];				l_cell_reg[180] = inform_L[180][2];				l_cell_reg[181] = inform_L[182][2];				l_cell_reg[182] = inform_L[181][2];				l_cell_reg[183] = inform_L[183][2];				l_cell_reg[184] = inform_L[184][2];				l_cell_reg[185] = inform_L[186][2];				l_cell_reg[186] = inform_L[185][2];				l_cell_reg[187] = inform_L[187][2];				l_cell_reg[188] = inform_L[188][2];				l_cell_reg[189] = inform_L[190][2];				l_cell_reg[190] = inform_L[189][2];				l_cell_reg[191] = inform_L[191][2];				l_cell_reg[192] = inform_L[192][2];				l_cell_reg[193] = inform_L[194][2];				l_cell_reg[194] = inform_L[193][2];				l_cell_reg[195] = inform_L[195][2];				l_cell_reg[196] = inform_L[196][2];				l_cell_reg[197] = inform_L[198][2];				l_cell_reg[198] = inform_L[197][2];				l_cell_reg[199] = inform_L[199][2];				l_cell_reg[200] = inform_L[200][2];				l_cell_reg[201] = inform_L[202][2];				l_cell_reg[202] = inform_L[201][2];				l_cell_reg[203] = inform_L[203][2];				l_cell_reg[204] = inform_L[204][2];				l_cell_reg[205] = inform_L[206][2];				l_cell_reg[206] = inform_L[205][2];				l_cell_reg[207] = inform_L[207][2];				l_cell_reg[208] = inform_L[208][2];				l_cell_reg[209] = inform_L[210][2];				l_cell_reg[210] = inform_L[209][2];				l_cell_reg[211] = inform_L[211][2];				l_cell_reg[212] = inform_L[212][2];				l_cell_reg[213] = inform_L[214][2];				l_cell_reg[214] = inform_L[213][2];				l_cell_reg[215] = inform_L[215][2];				l_cell_reg[216] = inform_L[216][2];				l_cell_reg[217] = inform_L[218][2];				l_cell_reg[218] = inform_L[217][2];				l_cell_reg[219] = inform_L[219][2];				l_cell_reg[220] = inform_L[220][2];				l_cell_reg[221] = inform_L[222][2];				l_cell_reg[222] = inform_L[221][2];				l_cell_reg[223] = inform_L[223][2];				l_cell_reg[224] = inform_L[224][2];				l_cell_reg[225] = inform_L[226][2];				l_cell_reg[226] = inform_L[225][2];				l_cell_reg[227] = inform_L[227][2];				l_cell_reg[228] = inform_L[228][2];				l_cell_reg[229] = inform_L[230][2];				l_cell_reg[230] = inform_L[229][2];				l_cell_reg[231] = inform_L[231][2];				l_cell_reg[232] = inform_L[232][2];				l_cell_reg[233] = inform_L[234][2];				l_cell_reg[234] = inform_L[233][2];				l_cell_reg[235] = inform_L[235][2];				l_cell_reg[236] = inform_L[236][2];				l_cell_reg[237] = inform_L[238][2];				l_cell_reg[238] = inform_L[237][2];				l_cell_reg[239] = inform_L[239][2];				l_cell_reg[240] = inform_L[240][2];				l_cell_reg[241] = inform_L[242][2];				l_cell_reg[242] = inform_L[241][2];				l_cell_reg[243] = inform_L[243][2];				l_cell_reg[244] = inform_L[244][2];				l_cell_reg[245] = inform_L[246][2];				l_cell_reg[246] = inform_L[245][2];				l_cell_reg[247] = inform_L[247][2];				l_cell_reg[248] = inform_L[248][2];				l_cell_reg[249] = inform_L[250][2];				l_cell_reg[250] = inform_L[249][2];				l_cell_reg[251] = inform_L[251][2];				l_cell_reg[252] = inform_L[252][2];				l_cell_reg[253] = inform_L[254][2];				l_cell_reg[254] = inform_L[253][2];				l_cell_reg[255] = inform_L[255][2];			end
			3:			begin				r_cell_reg[0] = inform_R[0][2];				r_cell_reg[1] = inform_R[4][2];				r_cell_reg[2] = inform_R[1][2];				r_cell_reg[3] = inform_R[5][2];				r_cell_reg[4] = inform_R[2][2];				r_cell_reg[5] = inform_R[6][2];				r_cell_reg[6] = inform_R[3][2];				r_cell_reg[7] = inform_R[7][2];				r_cell_reg[8] = inform_R[8][2];				r_cell_reg[9] = inform_R[12][2];				r_cell_reg[10] = inform_R[9][2];				r_cell_reg[11] = inform_R[13][2];				r_cell_reg[12] = inform_R[10][2];				r_cell_reg[13] = inform_R[14][2];				r_cell_reg[14] = inform_R[11][2];				r_cell_reg[15] = inform_R[15][2];				r_cell_reg[16] = inform_R[16][2];				r_cell_reg[17] = inform_R[20][2];				r_cell_reg[18] = inform_R[17][2];				r_cell_reg[19] = inform_R[21][2];				r_cell_reg[20] = inform_R[18][2];				r_cell_reg[21] = inform_R[22][2];				r_cell_reg[22] = inform_R[19][2];				r_cell_reg[23] = inform_R[23][2];				r_cell_reg[24] = inform_R[24][2];				r_cell_reg[25] = inform_R[28][2];				r_cell_reg[26] = inform_R[25][2];				r_cell_reg[27] = inform_R[29][2];				r_cell_reg[28] = inform_R[26][2];				r_cell_reg[29] = inform_R[30][2];				r_cell_reg[30] = inform_R[27][2];				r_cell_reg[31] = inform_R[31][2];				r_cell_reg[32] = inform_R[32][2];				r_cell_reg[33] = inform_R[36][2];				r_cell_reg[34] = inform_R[33][2];				r_cell_reg[35] = inform_R[37][2];				r_cell_reg[36] = inform_R[34][2];				r_cell_reg[37] = inform_R[38][2];				r_cell_reg[38] = inform_R[35][2];				r_cell_reg[39] = inform_R[39][2];				r_cell_reg[40] = inform_R[40][2];				r_cell_reg[41] = inform_R[44][2];				r_cell_reg[42] = inform_R[41][2];				r_cell_reg[43] = inform_R[45][2];				r_cell_reg[44] = inform_R[42][2];				r_cell_reg[45] = inform_R[46][2];				r_cell_reg[46] = inform_R[43][2];				r_cell_reg[47] = inform_R[47][2];				r_cell_reg[48] = inform_R[48][2];				r_cell_reg[49] = inform_R[52][2];				r_cell_reg[50] = inform_R[49][2];				r_cell_reg[51] = inform_R[53][2];				r_cell_reg[52] = inform_R[50][2];				r_cell_reg[53] = inform_R[54][2];				r_cell_reg[54] = inform_R[51][2];				r_cell_reg[55] = inform_R[55][2];				r_cell_reg[56] = inform_R[56][2];				r_cell_reg[57] = inform_R[60][2];				r_cell_reg[58] = inform_R[57][2];				r_cell_reg[59] = inform_R[61][2];				r_cell_reg[60] = inform_R[58][2];				r_cell_reg[61] = inform_R[62][2];				r_cell_reg[62] = inform_R[59][2];				r_cell_reg[63] = inform_R[63][2];				r_cell_reg[64] = inform_R[64][2];				r_cell_reg[65] = inform_R[68][2];				r_cell_reg[66] = inform_R[65][2];				r_cell_reg[67] = inform_R[69][2];				r_cell_reg[68] = inform_R[66][2];				r_cell_reg[69] = inform_R[70][2];				r_cell_reg[70] = inform_R[67][2];				r_cell_reg[71] = inform_R[71][2];				r_cell_reg[72] = inform_R[72][2];				r_cell_reg[73] = inform_R[76][2];				r_cell_reg[74] = inform_R[73][2];				r_cell_reg[75] = inform_R[77][2];				r_cell_reg[76] = inform_R[74][2];				r_cell_reg[77] = inform_R[78][2];				r_cell_reg[78] = inform_R[75][2];				r_cell_reg[79] = inform_R[79][2];				r_cell_reg[80] = inform_R[80][2];				r_cell_reg[81] = inform_R[84][2];				r_cell_reg[82] = inform_R[81][2];				r_cell_reg[83] = inform_R[85][2];				r_cell_reg[84] = inform_R[82][2];				r_cell_reg[85] = inform_R[86][2];				r_cell_reg[86] = inform_R[83][2];				r_cell_reg[87] = inform_R[87][2];				r_cell_reg[88] = inform_R[88][2];				r_cell_reg[89] = inform_R[92][2];				r_cell_reg[90] = inform_R[89][2];				r_cell_reg[91] = inform_R[93][2];				r_cell_reg[92] = inform_R[90][2];				r_cell_reg[93] = inform_R[94][2];				r_cell_reg[94] = inform_R[91][2];				r_cell_reg[95] = inform_R[95][2];				r_cell_reg[96] = inform_R[96][2];				r_cell_reg[97] = inform_R[100][2];				r_cell_reg[98] = inform_R[97][2];				r_cell_reg[99] = inform_R[101][2];				r_cell_reg[100] = inform_R[98][2];				r_cell_reg[101] = inform_R[102][2];				r_cell_reg[102] = inform_R[99][2];				r_cell_reg[103] = inform_R[103][2];				r_cell_reg[104] = inform_R[104][2];				r_cell_reg[105] = inform_R[108][2];				r_cell_reg[106] = inform_R[105][2];				r_cell_reg[107] = inform_R[109][2];				r_cell_reg[108] = inform_R[106][2];				r_cell_reg[109] = inform_R[110][2];				r_cell_reg[110] = inform_R[107][2];				r_cell_reg[111] = inform_R[111][2];				r_cell_reg[112] = inform_R[112][2];				r_cell_reg[113] = inform_R[116][2];				r_cell_reg[114] = inform_R[113][2];				r_cell_reg[115] = inform_R[117][2];				r_cell_reg[116] = inform_R[114][2];				r_cell_reg[117] = inform_R[118][2];				r_cell_reg[118] = inform_R[115][2];				r_cell_reg[119] = inform_R[119][2];				r_cell_reg[120] = inform_R[120][2];				r_cell_reg[121] = inform_R[124][2];				r_cell_reg[122] = inform_R[121][2];				r_cell_reg[123] = inform_R[125][2];				r_cell_reg[124] = inform_R[122][2];				r_cell_reg[125] = inform_R[126][2];				r_cell_reg[126] = inform_R[123][2];				r_cell_reg[127] = inform_R[127][2];				r_cell_reg[128] = inform_R[128][2];				r_cell_reg[129] = inform_R[132][2];				r_cell_reg[130] = inform_R[129][2];				r_cell_reg[131] = inform_R[133][2];				r_cell_reg[132] = inform_R[130][2];				r_cell_reg[133] = inform_R[134][2];				r_cell_reg[134] = inform_R[131][2];				r_cell_reg[135] = inform_R[135][2];				r_cell_reg[136] = inform_R[136][2];				r_cell_reg[137] = inform_R[140][2];				r_cell_reg[138] = inform_R[137][2];				r_cell_reg[139] = inform_R[141][2];				r_cell_reg[140] = inform_R[138][2];				r_cell_reg[141] = inform_R[142][2];				r_cell_reg[142] = inform_R[139][2];				r_cell_reg[143] = inform_R[143][2];				r_cell_reg[144] = inform_R[144][2];				r_cell_reg[145] = inform_R[148][2];				r_cell_reg[146] = inform_R[145][2];				r_cell_reg[147] = inform_R[149][2];				r_cell_reg[148] = inform_R[146][2];				r_cell_reg[149] = inform_R[150][2];				r_cell_reg[150] = inform_R[147][2];				r_cell_reg[151] = inform_R[151][2];				r_cell_reg[152] = inform_R[152][2];				r_cell_reg[153] = inform_R[156][2];				r_cell_reg[154] = inform_R[153][2];				r_cell_reg[155] = inform_R[157][2];				r_cell_reg[156] = inform_R[154][2];				r_cell_reg[157] = inform_R[158][2];				r_cell_reg[158] = inform_R[155][2];				r_cell_reg[159] = inform_R[159][2];				r_cell_reg[160] = inform_R[160][2];				r_cell_reg[161] = inform_R[164][2];				r_cell_reg[162] = inform_R[161][2];				r_cell_reg[163] = inform_R[165][2];				r_cell_reg[164] = inform_R[162][2];				r_cell_reg[165] = inform_R[166][2];				r_cell_reg[166] = inform_R[163][2];				r_cell_reg[167] = inform_R[167][2];				r_cell_reg[168] = inform_R[168][2];				r_cell_reg[169] = inform_R[172][2];				r_cell_reg[170] = inform_R[169][2];				r_cell_reg[171] = inform_R[173][2];				r_cell_reg[172] = inform_R[170][2];				r_cell_reg[173] = inform_R[174][2];				r_cell_reg[174] = inform_R[171][2];				r_cell_reg[175] = inform_R[175][2];				r_cell_reg[176] = inform_R[176][2];				r_cell_reg[177] = inform_R[180][2];				r_cell_reg[178] = inform_R[177][2];				r_cell_reg[179] = inform_R[181][2];				r_cell_reg[180] = inform_R[178][2];				r_cell_reg[181] = inform_R[182][2];				r_cell_reg[182] = inform_R[179][2];				r_cell_reg[183] = inform_R[183][2];				r_cell_reg[184] = inform_R[184][2];				r_cell_reg[185] = inform_R[188][2];				r_cell_reg[186] = inform_R[185][2];				r_cell_reg[187] = inform_R[189][2];				r_cell_reg[188] = inform_R[186][2];				r_cell_reg[189] = inform_R[190][2];				r_cell_reg[190] = inform_R[187][2];				r_cell_reg[191] = inform_R[191][2];				r_cell_reg[192] = inform_R[192][2];				r_cell_reg[193] = inform_R[196][2];				r_cell_reg[194] = inform_R[193][2];				r_cell_reg[195] = inform_R[197][2];				r_cell_reg[196] = inform_R[194][2];				r_cell_reg[197] = inform_R[198][2];				r_cell_reg[198] = inform_R[195][2];				r_cell_reg[199] = inform_R[199][2];				r_cell_reg[200] = inform_R[200][2];				r_cell_reg[201] = inform_R[204][2];				r_cell_reg[202] = inform_R[201][2];				r_cell_reg[203] = inform_R[205][2];				r_cell_reg[204] = inform_R[202][2];				r_cell_reg[205] = inform_R[206][2];				r_cell_reg[206] = inform_R[203][2];				r_cell_reg[207] = inform_R[207][2];				r_cell_reg[208] = inform_R[208][2];				r_cell_reg[209] = inform_R[212][2];				r_cell_reg[210] = inform_R[209][2];				r_cell_reg[211] = inform_R[213][2];				r_cell_reg[212] = inform_R[210][2];				r_cell_reg[213] = inform_R[214][2];				r_cell_reg[214] = inform_R[211][2];				r_cell_reg[215] = inform_R[215][2];				r_cell_reg[216] = inform_R[216][2];				r_cell_reg[217] = inform_R[220][2];				r_cell_reg[218] = inform_R[217][2];				r_cell_reg[219] = inform_R[221][2];				r_cell_reg[220] = inform_R[218][2];				r_cell_reg[221] = inform_R[222][2];				r_cell_reg[222] = inform_R[219][2];				r_cell_reg[223] = inform_R[223][2];				r_cell_reg[224] = inform_R[224][2];				r_cell_reg[225] = inform_R[228][2];				r_cell_reg[226] = inform_R[225][2];				r_cell_reg[227] = inform_R[229][2];				r_cell_reg[228] = inform_R[226][2];				r_cell_reg[229] = inform_R[230][2];				r_cell_reg[230] = inform_R[227][2];				r_cell_reg[231] = inform_R[231][2];				r_cell_reg[232] = inform_R[232][2];				r_cell_reg[233] = inform_R[236][2];				r_cell_reg[234] = inform_R[233][2];				r_cell_reg[235] = inform_R[237][2];				r_cell_reg[236] = inform_R[234][2];				r_cell_reg[237] = inform_R[238][2];				r_cell_reg[238] = inform_R[235][2];				r_cell_reg[239] = inform_R[239][2];				r_cell_reg[240] = inform_R[240][2];				r_cell_reg[241] = inform_R[244][2];				r_cell_reg[242] = inform_R[241][2];				r_cell_reg[243] = inform_R[245][2];				r_cell_reg[244] = inform_R[242][2];				r_cell_reg[245] = inform_R[246][2];				r_cell_reg[246] = inform_R[243][2];				r_cell_reg[247] = inform_R[247][2];				r_cell_reg[248] = inform_R[248][2];				r_cell_reg[249] = inform_R[252][2];				r_cell_reg[250] = inform_R[249][2];				r_cell_reg[251] = inform_R[253][2];				r_cell_reg[252] = inform_R[250][2];				r_cell_reg[253] = inform_R[254][2];				r_cell_reg[254] = inform_R[251][2];				r_cell_reg[255] = inform_R[255][2];				l_cell_reg[0] = inform_L[0][3];				l_cell_reg[1] = inform_L[4][3];				l_cell_reg[2] = inform_L[1][3];				l_cell_reg[3] = inform_L[5][3];				l_cell_reg[4] = inform_L[2][3];				l_cell_reg[5] = inform_L[6][3];				l_cell_reg[6] = inform_L[3][3];				l_cell_reg[7] = inform_L[7][3];				l_cell_reg[8] = inform_L[8][3];				l_cell_reg[9] = inform_L[12][3];				l_cell_reg[10] = inform_L[9][3];				l_cell_reg[11] = inform_L[13][3];				l_cell_reg[12] = inform_L[10][3];				l_cell_reg[13] = inform_L[14][3];				l_cell_reg[14] = inform_L[11][3];				l_cell_reg[15] = inform_L[15][3];				l_cell_reg[16] = inform_L[16][3];				l_cell_reg[17] = inform_L[20][3];				l_cell_reg[18] = inform_L[17][3];				l_cell_reg[19] = inform_L[21][3];				l_cell_reg[20] = inform_L[18][3];				l_cell_reg[21] = inform_L[22][3];				l_cell_reg[22] = inform_L[19][3];				l_cell_reg[23] = inform_L[23][3];				l_cell_reg[24] = inform_L[24][3];				l_cell_reg[25] = inform_L[28][3];				l_cell_reg[26] = inform_L[25][3];				l_cell_reg[27] = inform_L[29][3];				l_cell_reg[28] = inform_L[26][3];				l_cell_reg[29] = inform_L[30][3];				l_cell_reg[30] = inform_L[27][3];				l_cell_reg[31] = inform_L[31][3];				l_cell_reg[32] = inform_L[32][3];				l_cell_reg[33] = inform_L[36][3];				l_cell_reg[34] = inform_L[33][3];				l_cell_reg[35] = inform_L[37][3];				l_cell_reg[36] = inform_L[34][3];				l_cell_reg[37] = inform_L[38][3];				l_cell_reg[38] = inform_L[35][3];				l_cell_reg[39] = inform_L[39][3];				l_cell_reg[40] = inform_L[40][3];				l_cell_reg[41] = inform_L[44][3];				l_cell_reg[42] = inform_L[41][3];				l_cell_reg[43] = inform_L[45][3];				l_cell_reg[44] = inform_L[42][3];				l_cell_reg[45] = inform_L[46][3];				l_cell_reg[46] = inform_L[43][3];				l_cell_reg[47] = inform_L[47][3];				l_cell_reg[48] = inform_L[48][3];				l_cell_reg[49] = inform_L[52][3];				l_cell_reg[50] = inform_L[49][3];				l_cell_reg[51] = inform_L[53][3];				l_cell_reg[52] = inform_L[50][3];				l_cell_reg[53] = inform_L[54][3];				l_cell_reg[54] = inform_L[51][3];				l_cell_reg[55] = inform_L[55][3];				l_cell_reg[56] = inform_L[56][3];				l_cell_reg[57] = inform_L[60][3];				l_cell_reg[58] = inform_L[57][3];				l_cell_reg[59] = inform_L[61][3];				l_cell_reg[60] = inform_L[58][3];				l_cell_reg[61] = inform_L[62][3];				l_cell_reg[62] = inform_L[59][3];				l_cell_reg[63] = inform_L[63][3];				l_cell_reg[64] = inform_L[64][3];				l_cell_reg[65] = inform_L[68][3];				l_cell_reg[66] = inform_L[65][3];				l_cell_reg[67] = inform_L[69][3];				l_cell_reg[68] = inform_L[66][3];				l_cell_reg[69] = inform_L[70][3];				l_cell_reg[70] = inform_L[67][3];				l_cell_reg[71] = inform_L[71][3];				l_cell_reg[72] = inform_L[72][3];				l_cell_reg[73] = inform_L[76][3];				l_cell_reg[74] = inform_L[73][3];				l_cell_reg[75] = inform_L[77][3];				l_cell_reg[76] = inform_L[74][3];				l_cell_reg[77] = inform_L[78][3];				l_cell_reg[78] = inform_L[75][3];				l_cell_reg[79] = inform_L[79][3];				l_cell_reg[80] = inform_L[80][3];				l_cell_reg[81] = inform_L[84][3];				l_cell_reg[82] = inform_L[81][3];				l_cell_reg[83] = inform_L[85][3];				l_cell_reg[84] = inform_L[82][3];				l_cell_reg[85] = inform_L[86][3];				l_cell_reg[86] = inform_L[83][3];				l_cell_reg[87] = inform_L[87][3];				l_cell_reg[88] = inform_L[88][3];				l_cell_reg[89] = inform_L[92][3];				l_cell_reg[90] = inform_L[89][3];				l_cell_reg[91] = inform_L[93][3];				l_cell_reg[92] = inform_L[90][3];				l_cell_reg[93] = inform_L[94][3];				l_cell_reg[94] = inform_L[91][3];				l_cell_reg[95] = inform_L[95][3];				l_cell_reg[96] = inform_L[96][3];				l_cell_reg[97] = inform_L[100][3];				l_cell_reg[98] = inform_L[97][3];				l_cell_reg[99] = inform_L[101][3];				l_cell_reg[100] = inform_L[98][3];				l_cell_reg[101] = inform_L[102][3];				l_cell_reg[102] = inform_L[99][3];				l_cell_reg[103] = inform_L[103][3];				l_cell_reg[104] = inform_L[104][3];				l_cell_reg[105] = inform_L[108][3];				l_cell_reg[106] = inform_L[105][3];				l_cell_reg[107] = inform_L[109][3];				l_cell_reg[108] = inform_L[106][3];				l_cell_reg[109] = inform_L[110][3];				l_cell_reg[110] = inform_L[107][3];				l_cell_reg[111] = inform_L[111][3];				l_cell_reg[112] = inform_L[112][3];				l_cell_reg[113] = inform_L[116][3];				l_cell_reg[114] = inform_L[113][3];				l_cell_reg[115] = inform_L[117][3];				l_cell_reg[116] = inform_L[114][3];				l_cell_reg[117] = inform_L[118][3];				l_cell_reg[118] = inform_L[115][3];				l_cell_reg[119] = inform_L[119][3];				l_cell_reg[120] = inform_L[120][3];				l_cell_reg[121] = inform_L[124][3];				l_cell_reg[122] = inform_L[121][3];				l_cell_reg[123] = inform_L[125][3];				l_cell_reg[124] = inform_L[122][3];				l_cell_reg[125] = inform_L[126][3];				l_cell_reg[126] = inform_L[123][3];				l_cell_reg[127] = inform_L[127][3];				l_cell_reg[128] = inform_L[128][3];				l_cell_reg[129] = inform_L[132][3];				l_cell_reg[130] = inform_L[129][3];				l_cell_reg[131] = inform_L[133][3];				l_cell_reg[132] = inform_L[130][3];				l_cell_reg[133] = inform_L[134][3];				l_cell_reg[134] = inform_L[131][3];				l_cell_reg[135] = inform_L[135][3];				l_cell_reg[136] = inform_L[136][3];				l_cell_reg[137] = inform_L[140][3];				l_cell_reg[138] = inform_L[137][3];				l_cell_reg[139] = inform_L[141][3];				l_cell_reg[140] = inform_L[138][3];				l_cell_reg[141] = inform_L[142][3];				l_cell_reg[142] = inform_L[139][3];				l_cell_reg[143] = inform_L[143][3];				l_cell_reg[144] = inform_L[144][3];				l_cell_reg[145] = inform_L[148][3];				l_cell_reg[146] = inform_L[145][3];				l_cell_reg[147] = inform_L[149][3];				l_cell_reg[148] = inform_L[146][3];				l_cell_reg[149] = inform_L[150][3];				l_cell_reg[150] = inform_L[147][3];				l_cell_reg[151] = inform_L[151][3];				l_cell_reg[152] = inform_L[152][3];				l_cell_reg[153] = inform_L[156][3];				l_cell_reg[154] = inform_L[153][3];				l_cell_reg[155] = inform_L[157][3];				l_cell_reg[156] = inform_L[154][3];				l_cell_reg[157] = inform_L[158][3];				l_cell_reg[158] = inform_L[155][3];				l_cell_reg[159] = inform_L[159][3];				l_cell_reg[160] = inform_L[160][3];				l_cell_reg[161] = inform_L[164][3];				l_cell_reg[162] = inform_L[161][3];				l_cell_reg[163] = inform_L[165][3];				l_cell_reg[164] = inform_L[162][3];				l_cell_reg[165] = inform_L[166][3];				l_cell_reg[166] = inform_L[163][3];				l_cell_reg[167] = inform_L[167][3];				l_cell_reg[168] = inform_L[168][3];				l_cell_reg[169] = inform_L[172][3];				l_cell_reg[170] = inform_L[169][3];				l_cell_reg[171] = inform_L[173][3];				l_cell_reg[172] = inform_L[170][3];				l_cell_reg[173] = inform_L[174][3];				l_cell_reg[174] = inform_L[171][3];				l_cell_reg[175] = inform_L[175][3];				l_cell_reg[176] = inform_L[176][3];				l_cell_reg[177] = inform_L[180][3];				l_cell_reg[178] = inform_L[177][3];				l_cell_reg[179] = inform_L[181][3];				l_cell_reg[180] = inform_L[178][3];				l_cell_reg[181] = inform_L[182][3];				l_cell_reg[182] = inform_L[179][3];				l_cell_reg[183] = inform_L[183][3];				l_cell_reg[184] = inform_L[184][3];				l_cell_reg[185] = inform_L[188][3];				l_cell_reg[186] = inform_L[185][3];				l_cell_reg[187] = inform_L[189][3];				l_cell_reg[188] = inform_L[186][3];				l_cell_reg[189] = inform_L[190][3];				l_cell_reg[190] = inform_L[187][3];				l_cell_reg[191] = inform_L[191][3];				l_cell_reg[192] = inform_L[192][3];				l_cell_reg[193] = inform_L[196][3];				l_cell_reg[194] = inform_L[193][3];				l_cell_reg[195] = inform_L[197][3];				l_cell_reg[196] = inform_L[194][3];				l_cell_reg[197] = inform_L[198][3];				l_cell_reg[198] = inform_L[195][3];				l_cell_reg[199] = inform_L[199][3];				l_cell_reg[200] = inform_L[200][3];				l_cell_reg[201] = inform_L[204][3];				l_cell_reg[202] = inform_L[201][3];				l_cell_reg[203] = inform_L[205][3];				l_cell_reg[204] = inform_L[202][3];				l_cell_reg[205] = inform_L[206][3];				l_cell_reg[206] = inform_L[203][3];				l_cell_reg[207] = inform_L[207][3];				l_cell_reg[208] = inform_L[208][3];				l_cell_reg[209] = inform_L[212][3];				l_cell_reg[210] = inform_L[209][3];				l_cell_reg[211] = inform_L[213][3];				l_cell_reg[212] = inform_L[210][3];				l_cell_reg[213] = inform_L[214][3];				l_cell_reg[214] = inform_L[211][3];				l_cell_reg[215] = inform_L[215][3];				l_cell_reg[216] = inform_L[216][3];				l_cell_reg[217] = inform_L[220][3];				l_cell_reg[218] = inform_L[217][3];				l_cell_reg[219] = inform_L[221][3];				l_cell_reg[220] = inform_L[218][3];				l_cell_reg[221] = inform_L[222][3];				l_cell_reg[222] = inform_L[219][3];				l_cell_reg[223] = inform_L[223][3];				l_cell_reg[224] = inform_L[224][3];				l_cell_reg[225] = inform_L[228][3];				l_cell_reg[226] = inform_L[225][3];				l_cell_reg[227] = inform_L[229][3];				l_cell_reg[228] = inform_L[226][3];				l_cell_reg[229] = inform_L[230][3];				l_cell_reg[230] = inform_L[227][3];				l_cell_reg[231] = inform_L[231][3];				l_cell_reg[232] = inform_L[232][3];				l_cell_reg[233] = inform_L[236][3];				l_cell_reg[234] = inform_L[233][3];				l_cell_reg[235] = inform_L[237][3];				l_cell_reg[236] = inform_L[234][3];				l_cell_reg[237] = inform_L[238][3];				l_cell_reg[238] = inform_L[235][3];				l_cell_reg[239] = inform_L[239][3];				l_cell_reg[240] = inform_L[240][3];				l_cell_reg[241] = inform_L[244][3];				l_cell_reg[242] = inform_L[241][3];				l_cell_reg[243] = inform_L[245][3];				l_cell_reg[244] = inform_L[242][3];				l_cell_reg[245] = inform_L[246][3];				l_cell_reg[246] = inform_L[243][3];				l_cell_reg[247] = inform_L[247][3];				l_cell_reg[248] = inform_L[248][3];				l_cell_reg[249] = inform_L[252][3];				l_cell_reg[250] = inform_L[249][3];				l_cell_reg[251] = inform_L[253][3];				l_cell_reg[252] = inform_L[250][3];				l_cell_reg[253] = inform_L[254][3];				l_cell_reg[254] = inform_L[251][3];				l_cell_reg[255] = inform_L[255][3];			end
			4:			begin				r_cell_reg[0] = inform_R[0][3];				r_cell_reg[1] = inform_R[8][3];				r_cell_reg[2] = inform_R[1][3];				r_cell_reg[3] = inform_R[9][3];				r_cell_reg[4] = inform_R[2][3];				r_cell_reg[5] = inform_R[10][3];				r_cell_reg[6] = inform_R[3][3];				r_cell_reg[7] = inform_R[11][3];				r_cell_reg[8] = inform_R[4][3];				r_cell_reg[9] = inform_R[12][3];				r_cell_reg[10] = inform_R[5][3];				r_cell_reg[11] = inform_R[13][3];				r_cell_reg[12] = inform_R[6][3];				r_cell_reg[13] = inform_R[14][3];				r_cell_reg[14] = inform_R[7][3];				r_cell_reg[15] = inform_R[15][3];				r_cell_reg[16] = inform_R[16][3];				r_cell_reg[17] = inform_R[24][3];				r_cell_reg[18] = inform_R[17][3];				r_cell_reg[19] = inform_R[25][3];				r_cell_reg[20] = inform_R[18][3];				r_cell_reg[21] = inform_R[26][3];				r_cell_reg[22] = inform_R[19][3];				r_cell_reg[23] = inform_R[27][3];				r_cell_reg[24] = inform_R[20][3];				r_cell_reg[25] = inform_R[28][3];				r_cell_reg[26] = inform_R[21][3];				r_cell_reg[27] = inform_R[29][3];				r_cell_reg[28] = inform_R[22][3];				r_cell_reg[29] = inform_R[30][3];				r_cell_reg[30] = inform_R[23][3];				r_cell_reg[31] = inform_R[31][3];				r_cell_reg[32] = inform_R[32][3];				r_cell_reg[33] = inform_R[40][3];				r_cell_reg[34] = inform_R[33][3];				r_cell_reg[35] = inform_R[41][3];				r_cell_reg[36] = inform_R[34][3];				r_cell_reg[37] = inform_R[42][3];				r_cell_reg[38] = inform_R[35][3];				r_cell_reg[39] = inform_R[43][3];				r_cell_reg[40] = inform_R[36][3];				r_cell_reg[41] = inform_R[44][3];				r_cell_reg[42] = inform_R[37][3];				r_cell_reg[43] = inform_R[45][3];				r_cell_reg[44] = inform_R[38][3];				r_cell_reg[45] = inform_R[46][3];				r_cell_reg[46] = inform_R[39][3];				r_cell_reg[47] = inform_R[47][3];				r_cell_reg[48] = inform_R[48][3];				r_cell_reg[49] = inform_R[56][3];				r_cell_reg[50] = inform_R[49][3];				r_cell_reg[51] = inform_R[57][3];				r_cell_reg[52] = inform_R[50][3];				r_cell_reg[53] = inform_R[58][3];				r_cell_reg[54] = inform_R[51][3];				r_cell_reg[55] = inform_R[59][3];				r_cell_reg[56] = inform_R[52][3];				r_cell_reg[57] = inform_R[60][3];				r_cell_reg[58] = inform_R[53][3];				r_cell_reg[59] = inform_R[61][3];				r_cell_reg[60] = inform_R[54][3];				r_cell_reg[61] = inform_R[62][3];				r_cell_reg[62] = inform_R[55][3];				r_cell_reg[63] = inform_R[63][3];				r_cell_reg[64] = inform_R[64][3];				r_cell_reg[65] = inform_R[72][3];				r_cell_reg[66] = inform_R[65][3];				r_cell_reg[67] = inform_R[73][3];				r_cell_reg[68] = inform_R[66][3];				r_cell_reg[69] = inform_R[74][3];				r_cell_reg[70] = inform_R[67][3];				r_cell_reg[71] = inform_R[75][3];				r_cell_reg[72] = inform_R[68][3];				r_cell_reg[73] = inform_R[76][3];				r_cell_reg[74] = inform_R[69][3];				r_cell_reg[75] = inform_R[77][3];				r_cell_reg[76] = inform_R[70][3];				r_cell_reg[77] = inform_R[78][3];				r_cell_reg[78] = inform_R[71][3];				r_cell_reg[79] = inform_R[79][3];				r_cell_reg[80] = inform_R[80][3];				r_cell_reg[81] = inform_R[88][3];				r_cell_reg[82] = inform_R[81][3];				r_cell_reg[83] = inform_R[89][3];				r_cell_reg[84] = inform_R[82][3];				r_cell_reg[85] = inform_R[90][3];				r_cell_reg[86] = inform_R[83][3];				r_cell_reg[87] = inform_R[91][3];				r_cell_reg[88] = inform_R[84][3];				r_cell_reg[89] = inform_R[92][3];				r_cell_reg[90] = inform_R[85][3];				r_cell_reg[91] = inform_R[93][3];				r_cell_reg[92] = inform_R[86][3];				r_cell_reg[93] = inform_R[94][3];				r_cell_reg[94] = inform_R[87][3];				r_cell_reg[95] = inform_R[95][3];				r_cell_reg[96] = inform_R[96][3];				r_cell_reg[97] = inform_R[104][3];				r_cell_reg[98] = inform_R[97][3];				r_cell_reg[99] = inform_R[105][3];				r_cell_reg[100] = inform_R[98][3];				r_cell_reg[101] = inform_R[106][3];				r_cell_reg[102] = inform_R[99][3];				r_cell_reg[103] = inform_R[107][3];				r_cell_reg[104] = inform_R[100][3];				r_cell_reg[105] = inform_R[108][3];				r_cell_reg[106] = inform_R[101][3];				r_cell_reg[107] = inform_R[109][3];				r_cell_reg[108] = inform_R[102][3];				r_cell_reg[109] = inform_R[110][3];				r_cell_reg[110] = inform_R[103][3];				r_cell_reg[111] = inform_R[111][3];				r_cell_reg[112] = inform_R[112][3];				r_cell_reg[113] = inform_R[120][3];				r_cell_reg[114] = inform_R[113][3];				r_cell_reg[115] = inform_R[121][3];				r_cell_reg[116] = inform_R[114][3];				r_cell_reg[117] = inform_R[122][3];				r_cell_reg[118] = inform_R[115][3];				r_cell_reg[119] = inform_R[123][3];				r_cell_reg[120] = inform_R[116][3];				r_cell_reg[121] = inform_R[124][3];				r_cell_reg[122] = inform_R[117][3];				r_cell_reg[123] = inform_R[125][3];				r_cell_reg[124] = inform_R[118][3];				r_cell_reg[125] = inform_R[126][3];				r_cell_reg[126] = inform_R[119][3];				r_cell_reg[127] = inform_R[127][3];				r_cell_reg[128] = inform_R[128][3];				r_cell_reg[129] = inform_R[136][3];				r_cell_reg[130] = inform_R[129][3];				r_cell_reg[131] = inform_R[137][3];				r_cell_reg[132] = inform_R[130][3];				r_cell_reg[133] = inform_R[138][3];				r_cell_reg[134] = inform_R[131][3];				r_cell_reg[135] = inform_R[139][3];				r_cell_reg[136] = inform_R[132][3];				r_cell_reg[137] = inform_R[140][3];				r_cell_reg[138] = inform_R[133][3];				r_cell_reg[139] = inform_R[141][3];				r_cell_reg[140] = inform_R[134][3];				r_cell_reg[141] = inform_R[142][3];				r_cell_reg[142] = inform_R[135][3];				r_cell_reg[143] = inform_R[143][3];				r_cell_reg[144] = inform_R[144][3];				r_cell_reg[145] = inform_R[152][3];				r_cell_reg[146] = inform_R[145][3];				r_cell_reg[147] = inform_R[153][3];				r_cell_reg[148] = inform_R[146][3];				r_cell_reg[149] = inform_R[154][3];				r_cell_reg[150] = inform_R[147][3];				r_cell_reg[151] = inform_R[155][3];				r_cell_reg[152] = inform_R[148][3];				r_cell_reg[153] = inform_R[156][3];				r_cell_reg[154] = inform_R[149][3];				r_cell_reg[155] = inform_R[157][3];				r_cell_reg[156] = inform_R[150][3];				r_cell_reg[157] = inform_R[158][3];				r_cell_reg[158] = inform_R[151][3];				r_cell_reg[159] = inform_R[159][3];				r_cell_reg[160] = inform_R[160][3];				r_cell_reg[161] = inform_R[168][3];				r_cell_reg[162] = inform_R[161][3];				r_cell_reg[163] = inform_R[169][3];				r_cell_reg[164] = inform_R[162][3];				r_cell_reg[165] = inform_R[170][3];				r_cell_reg[166] = inform_R[163][3];				r_cell_reg[167] = inform_R[171][3];				r_cell_reg[168] = inform_R[164][3];				r_cell_reg[169] = inform_R[172][3];				r_cell_reg[170] = inform_R[165][3];				r_cell_reg[171] = inform_R[173][3];				r_cell_reg[172] = inform_R[166][3];				r_cell_reg[173] = inform_R[174][3];				r_cell_reg[174] = inform_R[167][3];				r_cell_reg[175] = inform_R[175][3];				r_cell_reg[176] = inform_R[176][3];				r_cell_reg[177] = inform_R[184][3];				r_cell_reg[178] = inform_R[177][3];				r_cell_reg[179] = inform_R[185][3];				r_cell_reg[180] = inform_R[178][3];				r_cell_reg[181] = inform_R[186][3];				r_cell_reg[182] = inform_R[179][3];				r_cell_reg[183] = inform_R[187][3];				r_cell_reg[184] = inform_R[180][3];				r_cell_reg[185] = inform_R[188][3];				r_cell_reg[186] = inform_R[181][3];				r_cell_reg[187] = inform_R[189][3];				r_cell_reg[188] = inform_R[182][3];				r_cell_reg[189] = inform_R[190][3];				r_cell_reg[190] = inform_R[183][3];				r_cell_reg[191] = inform_R[191][3];				r_cell_reg[192] = inform_R[192][3];				r_cell_reg[193] = inform_R[200][3];				r_cell_reg[194] = inform_R[193][3];				r_cell_reg[195] = inform_R[201][3];				r_cell_reg[196] = inform_R[194][3];				r_cell_reg[197] = inform_R[202][3];				r_cell_reg[198] = inform_R[195][3];				r_cell_reg[199] = inform_R[203][3];				r_cell_reg[200] = inform_R[196][3];				r_cell_reg[201] = inform_R[204][3];				r_cell_reg[202] = inform_R[197][3];				r_cell_reg[203] = inform_R[205][3];				r_cell_reg[204] = inform_R[198][3];				r_cell_reg[205] = inform_R[206][3];				r_cell_reg[206] = inform_R[199][3];				r_cell_reg[207] = inform_R[207][3];				r_cell_reg[208] = inform_R[208][3];				r_cell_reg[209] = inform_R[216][3];				r_cell_reg[210] = inform_R[209][3];				r_cell_reg[211] = inform_R[217][3];				r_cell_reg[212] = inform_R[210][3];				r_cell_reg[213] = inform_R[218][3];				r_cell_reg[214] = inform_R[211][3];				r_cell_reg[215] = inform_R[219][3];				r_cell_reg[216] = inform_R[212][3];				r_cell_reg[217] = inform_R[220][3];				r_cell_reg[218] = inform_R[213][3];				r_cell_reg[219] = inform_R[221][3];				r_cell_reg[220] = inform_R[214][3];				r_cell_reg[221] = inform_R[222][3];				r_cell_reg[222] = inform_R[215][3];				r_cell_reg[223] = inform_R[223][3];				r_cell_reg[224] = inform_R[224][3];				r_cell_reg[225] = inform_R[232][3];				r_cell_reg[226] = inform_R[225][3];				r_cell_reg[227] = inform_R[233][3];				r_cell_reg[228] = inform_R[226][3];				r_cell_reg[229] = inform_R[234][3];				r_cell_reg[230] = inform_R[227][3];				r_cell_reg[231] = inform_R[235][3];				r_cell_reg[232] = inform_R[228][3];				r_cell_reg[233] = inform_R[236][3];				r_cell_reg[234] = inform_R[229][3];				r_cell_reg[235] = inform_R[237][3];				r_cell_reg[236] = inform_R[230][3];				r_cell_reg[237] = inform_R[238][3];				r_cell_reg[238] = inform_R[231][3];				r_cell_reg[239] = inform_R[239][3];				r_cell_reg[240] = inform_R[240][3];				r_cell_reg[241] = inform_R[248][3];				r_cell_reg[242] = inform_R[241][3];				r_cell_reg[243] = inform_R[249][3];				r_cell_reg[244] = inform_R[242][3];				r_cell_reg[245] = inform_R[250][3];				r_cell_reg[246] = inform_R[243][3];				r_cell_reg[247] = inform_R[251][3];				r_cell_reg[248] = inform_R[244][3];				r_cell_reg[249] = inform_R[252][3];				r_cell_reg[250] = inform_R[245][3];				r_cell_reg[251] = inform_R[253][3];				r_cell_reg[252] = inform_R[246][3];				r_cell_reg[253] = inform_R[254][3];				r_cell_reg[254] = inform_R[247][3];				r_cell_reg[255] = inform_R[255][3];				l_cell_reg[0] = inform_L[0][4];				l_cell_reg[1] = inform_L[8][4];				l_cell_reg[2] = inform_L[1][4];				l_cell_reg[3] = inform_L[9][4];				l_cell_reg[4] = inform_L[2][4];				l_cell_reg[5] = inform_L[10][4];				l_cell_reg[6] = inform_L[3][4];				l_cell_reg[7] = inform_L[11][4];				l_cell_reg[8] = inform_L[4][4];				l_cell_reg[9] = inform_L[12][4];				l_cell_reg[10] = inform_L[5][4];				l_cell_reg[11] = inform_L[13][4];				l_cell_reg[12] = inform_L[6][4];				l_cell_reg[13] = inform_L[14][4];				l_cell_reg[14] = inform_L[7][4];				l_cell_reg[15] = inform_L[15][4];				l_cell_reg[16] = inform_L[16][4];				l_cell_reg[17] = inform_L[24][4];				l_cell_reg[18] = inform_L[17][4];				l_cell_reg[19] = inform_L[25][4];				l_cell_reg[20] = inform_L[18][4];				l_cell_reg[21] = inform_L[26][4];				l_cell_reg[22] = inform_L[19][4];				l_cell_reg[23] = inform_L[27][4];				l_cell_reg[24] = inform_L[20][4];				l_cell_reg[25] = inform_L[28][4];				l_cell_reg[26] = inform_L[21][4];				l_cell_reg[27] = inform_L[29][4];				l_cell_reg[28] = inform_L[22][4];				l_cell_reg[29] = inform_L[30][4];				l_cell_reg[30] = inform_L[23][4];				l_cell_reg[31] = inform_L[31][4];				l_cell_reg[32] = inform_L[32][4];				l_cell_reg[33] = inform_L[40][4];				l_cell_reg[34] = inform_L[33][4];				l_cell_reg[35] = inform_L[41][4];				l_cell_reg[36] = inform_L[34][4];				l_cell_reg[37] = inform_L[42][4];				l_cell_reg[38] = inform_L[35][4];				l_cell_reg[39] = inform_L[43][4];				l_cell_reg[40] = inform_L[36][4];				l_cell_reg[41] = inform_L[44][4];				l_cell_reg[42] = inform_L[37][4];				l_cell_reg[43] = inform_L[45][4];				l_cell_reg[44] = inform_L[38][4];				l_cell_reg[45] = inform_L[46][4];				l_cell_reg[46] = inform_L[39][4];				l_cell_reg[47] = inform_L[47][4];				l_cell_reg[48] = inform_L[48][4];				l_cell_reg[49] = inform_L[56][4];				l_cell_reg[50] = inform_L[49][4];				l_cell_reg[51] = inform_L[57][4];				l_cell_reg[52] = inform_L[50][4];				l_cell_reg[53] = inform_L[58][4];				l_cell_reg[54] = inform_L[51][4];				l_cell_reg[55] = inform_L[59][4];				l_cell_reg[56] = inform_L[52][4];				l_cell_reg[57] = inform_L[60][4];				l_cell_reg[58] = inform_L[53][4];				l_cell_reg[59] = inform_L[61][4];				l_cell_reg[60] = inform_L[54][4];				l_cell_reg[61] = inform_L[62][4];				l_cell_reg[62] = inform_L[55][4];				l_cell_reg[63] = inform_L[63][4];				l_cell_reg[64] = inform_L[64][4];				l_cell_reg[65] = inform_L[72][4];				l_cell_reg[66] = inform_L[65][4];				l_cell_reg[67] = inform_L[73][4];				l_cell_reg[68] = inform_L[66][4];				l_cell_reg[69] = inform_L[74][4];				l_cell_reg[70] = inform_L[67][4];				l_cell_reg[71] = inform_L[75][4];				l_cell_reg[72] = inform_L[68][4];				l_cell_reg[73] = inform_L[76][4];				l_cell_reg[74] = inform_L[69][4];				l_cell_reg[75] = inform_L[77][4];				l_cell_reg[76] = inform_L[70][4];				l_cell_reg[77] = inform_L[78][4];				l_cell_reg[78] = inform_L[71][4];				l_cell_reg[79] = inform_L[79][4];				l_cell_reg[80] = inform_L[80][4];				l_cell_reg[81] = inform_L[88][4];				l_cell_reg[82] = inform_L[81][4];				l_cell_reg[83] = inform_L[89][4];				l_cell_reg[84] = inform_L[82][4];				l_cell_reg[85] = inform_L[90][4];				l_cell_reg[86] = inform_L[83][4];				l_cell_reg[87] = inform_L[91][4];				l_cell_reg[88] = inform_L[84][4];				l_cell_reg[89] = inform_L[92][4];				l_cell_reg[90] = inform_L[85][4];				l_cell_reg[91] = inform_L[93][4];				l_cell_reg[92] = inform_L[86][4];				l_cell_reg[93] = inform_L[94][4];				l_cell_reg[94] = inform_L[87][4];				l_cell_reg[95] = inform_L[95][4];				l_cell_reg[96] = inform_L[96][4];				l_cell_reg[97] = inform_L[104][4];				l_cell_reg[98] = inform_L[97][4];				l_cell_reg[99] = inform_L[105][4];				l_cell_reg[100] = inform_L[98][4];				l_cell_reg[101] = inform_L[106][4];				l_cell_reg[102] = inform_L[99][4];				l_cell_reg[103] = inform_L[107][4];				l_cell_reg[104] = inform_L[100][4];				l_cell_reg[105] = inform_L[108][4];				l_cell_reg[106] = inform_L[101][4];				l_cell_reg[107] = inform_L[109][4];				l_cell_reg[108] = inform_L[102][4];				l_cell_reg[109] = inform_L[110][4];				l_cell_reg[110] = inform_L[103][4];				l_cell_reg[111] = inform_L[111][4];				l_cell_reg[112] = inform_L[112][4];				l_cell_reg[113] = inform_L[120][4];				l_cell_reg[114] = inform_L[113][4];				l_cell_reg[115] = inform_L[121][4];				l_cell_reg[116] = inform_L[114][4];				l_cell_reg[117] = inform_L[122][4];				l_cell_reg[118] = inform_L[115][4];				l_cell_reg[119] = inform_L[123][4];				l_cell_reg[120] = inform_L[116][4];				l_cell_reg[121] = inform_L[124][4];				l_cell_reg[122] = inform_L[117][4];				l_cell_reg[123] = inform_L[125][4];				l_cell_reg[124] = inform_L[118][4];				l_cell_reg[125] = inform_L[126][4];				l_cell_reg[126] = inform_L[119][4];				l_cell_reg[127] = inform_L[127][4];				l_cell_reg[128] = inform_L[128][4];				l_cell_reg[129] = inform_L[136][4];				l_cell_reg[130] = inform_L[129][4];				l_cell_reg[131] = inform_L[137][4];				l_cell_reg[132] = inform_L[130][4];				l_cell_reg[133] = inform_L[138][4];				l_cell_reg[134] = inform_L[131][4];				l_cell_reg[135] = inform_L[139][4];				l_cell_reg[136] = inform_L[132][4];				l_cell_reg[137] = inform_L[140][4];				l_cell_reg[138] = inform_L[133][4];				l_cell_reg[139] = inform_L[141][4];				l_cell_reg[140] = inform_L[134][4];				l_cell_reg[141] = inform_L[142][4];				l_cell_reg[142] = inform_L[135][4];				l_cell_reg[143] = inform_L[143][4];				l_cell_reg[144] = inform_L[144][4];				l_cell_reg[145] = inform_L[152][4];				l_cell_reg[146] = inform_L[145][4];				l_cell_reg[147] = inform_L[153][4];				l_cell_reg[148] = inform_L[146][4];				l_cell_reg[149] = inform_L[154][4];				l_cell_reg[150] = inform_L[147][4];				l_cell_reg[151] = inform_L[155][4];				l_cell_reg[152] = inform_L[148][4];				l_cell_reg[153] = inform_L[156][4];				l_cell_reg[154] = inform_L[149][4];				l_cell_reg[155] = inform_L[157][4];				l_cell_reg[156] = inform_L[150][4];				l_cell_reg[157] = inform_L[158][4];				l_cell_reg[158] = inform_L[151][4];				l_cell_reg[159] = inform_L[159][4];				l_cell_reg[160] = inform_L[160][4];				l_cell_reg[161] = inform_L[168][4];				l_cell_reg[162] = inform_L[161][4];				l_cell_reg[163] = inform_L[169][4];				l_cell_reg[164] = inform_L[162][4];				l_cell_reg[165] = inform_L[170][4];				l_cell_reg[166] = inform_L[163][4];				l_cell_reg[167] = inform_L[171][4];				l_cell_reg[168] = inform_L[164][4];				l_cell_reg[169] = inform_L[172][4];				l_cell_reg[170] = inform_L[165][4];				l_cell_reg[171] = inform_L[173][4];				l_cell_reg[172] = inform_L[166][4];				l_cell_reg[173] = inform_L[174][4];				l_cell_reg[174] = inform_L[167][4];				l_cell_reg[175] = inform_L[175][4];				l_cell_reg[176] = inform_L[176][4];				l_cell_reg[177] = inform_L[184][4];				l_cell_reg[178] = inform_L[177][4];				l_cell_reg[179] = inform_L[185][4];				l_cell_reg[180] = inform_L[178][4];				l_cell_reg[181] = inform_L[186][4];				l_cell_reg[182] = inform_L[179][4];				l_cell_reg[183] = inform_L[187][4];				l_cell_reg[184] = inform_L[180][4];				l_cell_reg[185] = inform_L[188][4];				l_cell_reg[186] = inform_L[181][4];				l_cell_reg[187] = inform_L[189][4];				l_cell_reg[188] = inform_L[182][4];				l_cell_reg[189] = inform_L[190][4];				l_cell_reg[190] = inform_L[183][4];				l_cell_reg[191] = inform_L[191][4];				l_cell_reg[192] = inform_L[192][4];				l_cell_reg[193] = inform_L[200][4];				l_cell_reg[194] = inform_L[193][4];				l_cell_reg[195] = inform_L[201][4];				l_cell_reg[196] = inform_L[194][4];				l_cell_reg[197] = inform_L[202][4];				l_cell_reg[198] = inform_L[195][4];				l_cell_reg[199] = inform_L[203][4];				l_cell_reg[200] = inform_L[196][4];				l_cell_reg[201] = inform_L[204][4];				l_cell_reg[202] = inform_L[197][4];				l_cell_reg[203] = inform_L[205][4];				l_cell_reg[204] = inform_L[198][4];				l_cell_reg[205] = inform_L[206][4];				l_cell_reg[206] = inform_L[199][4];				l_cell_reg[207] = inform_L[207][4];				l_cell_reg[208] = inform_L[208][4];				l_cell_reg[209] = inform_L[216][4];				l_cell_reg[210] = inform_L[209][4];				l_cell_reg[211] = inform_L[217][4];				l_cell_reg[212] = inform_L[210][4];				l_cell_reg[213] = inform_L[218][4];				l_cell_reg[214] = inform_L[211][4];				l_cell_reg[215] = inform_L[219][4];				l_cell_reg[216] = inform_L[212][4];				l_cell_reg[217] = inform_L[220][4];				l_cell_reg[218] = inform_L[213][4];				l_cell_reg[219] = inform_L[221][4];				l_cell_reg[220] = inform_L[214][4];				l_cell_reg[221] = inform_L[222][4];				l_cell_reg[222] = inform_L[215][4];				l_cell_reg[223] = inform_L[223][4];				l_cell_reg[224] = inform_L[224][4];				l_cell_reg[225] = inform_L[232][4];				l_cell_reg[226] = inform_L[225][4];				l_cell_reg[227] = inform_L[233][4];				l_cell_reg[228] = inform_L[226][4];				l_cell_reg[229] = inform_L[234][4];				l_cell_reg[230] = inform_L[227][4];				l_cell_reg[231] = inform_L[235][4];				l_cell_reg[232] = inform_L[228][4];				l_cell_reg[233] = inform_L[236][4];				l_cell_reg[234] = inform_L[229][4];				l_cell_reg[235] = inform_L[237][4];				l_cell_reg[236] = inform_L[230][4];				l_cell_reg[237] = inform_L[238][4];				l_cell_reg[238] = inform_L[231][4];				l_cell_reg[239] = inform_L[239][4];				l_cell_reg[240] = inform_L[240][4];				l_cell_reg[241] = inform_L[248][4];				l_cell_reg[242] = inform_L[241][4];				l_cell_reg[243] = inform_L[249][4];				l_cell_reg[244] = inform_L[242][4];				l_cell_reg[245] = inform_L[250][4];				l_cell_reg[246] = inform_L[243][4];				l_cell_reg[247] = inform_L[251][4];				l_cell_reg[248] = inform_L[244][4];				l_cell_reg[249] = inform_L[252][4];				l_cell_reg[250] = inform_L[245][4];				l_cell_reg[251] = inform_L[253][4];				l_cell_reg[252] = inform_L[246][4];				l_cell_reg[253] = inform_L[254][4];				l_cell_reg[254] = inform_L[247][4];				l_cell_reg[255] = inform_L[255][4];			end
			5:			begin				r_cell_reg[0] = inform_R[0][4];				r_cell_reg[1] = inform_R[16][4];				r_cell_reg[2] = inform_R[1][4];				r_cell_reg[3] = inform_R[17][4];				r_cell_reg[4] = inform_R[2][4];				r_cell_reg[5] = inform_R[18][4];				r_cell_reg[6] = inform_R[3][4];				r_cell_reg[7] = inform_R[19][4];				r_cell_reg[8] = inform_R[4][4];				r_cell_reg[9] = inform_R[20][4];				r_cell_reg[10] = inform_R[5][4];				r_cell_reg[11] = inform_R[21][4];				r_cell_reg[12] = inform_R[6][4];				r_cell_reg[13] = inform_R[22][4];				r_cell_reg[14] = inform_R[7][4];				r_cell_reg[15] = inform_R[23][4];				r_cell_reg[16] = inform_R[8][4];				r_cell_reg[17] = inform_R[24][4];				r_cell_reg[18] = inform_R[9][4];				r_cell_reg[19] = inform_R[25][4];				r_cell_reg[20] = inform_R[10][4];				r_cell_reg[21] = inform_R[26][4];				r_cell_reg[22] = inform_R[11][4];				r_cell_reg[23] = inform_R[27][4];				r_cell_reg[24] = inform_R[12][4];				r_cell_reg[25] = inform_R[28][4];				r_cell_reg[26] = inform_R[13][4];				r_cell_reg[27] = inform_R[29][4];				r_cell_reg[28] = inform_R[14][4];				r_cell_reg[29] = inform_R[30][4];				r_cell_reg[30] = inform_R[15][4];				r_cell_reg[31] = inform_R[31][4];				r_cell_reg[32] = inform_R[32][4];				r_cell_reg[33] = inform_R[48][4];				r_cell_reg[34] = inform_R[33][4];				r_cell_reg[35] = inform_R[49][4];				r_cell_reg[36] = inform_R[34][4];				r_cell_reg[37] = inform_R[50][4];				r_cell_reg[38] = inform_R[35][4];				r_cell_reg[39] = inform_R[51][4];				r_cell_reg[40] = inform_R[36][4];				r_cell_reg[41] = inform_R[52][4];				r_cell_reg[42] = inform_R[37][4];				r_cell_reg[43] = inform_R[53][4];				r_cell_reg[44] = inform_R[38][4];				r_cell_reg[45] = inform_R[54][4];				r_cell_reg[46] = inform_R[39][4];				r_cell_reg[47] = inform_R[55][4];				r_cell_reg[48] = inform_R[40][4];				r_cell_reg[49] = inform_R[56][4];				r_cell_reg[50] = inform_R[41][4];				r_cell_reg[51] = inform_R[57][4];				r_cell_reg[52] = inform_R[42][4];				r_cell_reg[53] = inform_R[58][4];				r_cell_reg[54] = inform_R[43][4];				r_cell_reg[55] = inform_R[59][4];				r_cell_reg[56] = inform_R[44][4];				r_cell_reg[57] = inform_R[60][4];				r_cell_reg[58] = inform_R[45][4];				r_cell_reg[59] = inform_R[61][4];				r_cell_reg[60] = inform_R[46][4];				r_cell_reg[61] = inform_R[62][4];				r_cell_reg[62] = inform_R[47][4];				r_cell_reg[63] = inform_R[63][4];				r_cell_reg[64] = inform_R[64][4];				r_cell_reg[65] = inform_R[80][4];				r_cell_reg[66] = inform_R[65][4];				r_cell_reg[67] = inform_R[81][4];				r_cell_reg[68] = inform_R[66][4];				r_cell_reg[69] = inform_R[82][4];				r_cell_reg[70] = inform_R[67][4];				r_cell_reg[71] = inform_R[83][4];				r_cell_reg[72] = inform_R[68][4];				r_cell_reg[73] = inform_R[84][4];				r_cell_reg[74] = inform_R[69][4];				r_cell_reg[75] = inform_R[85][4];				r_cell_reg[76] = inform_R[70][4];				r_cell_reg[77] = inform_R[86][4];				r_cell_reg[78] = inform_R[71][4];				r_cell_reg[79] = inform_R[87][4];				r_cell_reg[80] = inform_R[72][4];				r_cell_reg[81] = inform_R[88][4];				r_cell_reg[82] = inform_R[73][4];				r_cell_reg[83] = inform_R[89][4];				r_cell_reg[84] = inform_R[74][4];				r_cell_reg[85] = inform_R[90][4];				r_cell_reg[86] = inform_R[75][4];				r_cell_reg[87] = inform_R[91][4];				r_cell_reg[88] = inform_R[76][4];				r_cell_reg[89] = inform_R[92][4];				r_cell_reg[90] = inform_R[77][4];				r_cell_reg[91] = inform_R[93][4];				r_cell_reg[92] = inform_R[78][4];				r_cell_reg[93] = inform_R[94][4];				r_cell_reg[94] = inform_R[79][4];				r_cell_reg[95] = inform_R[95][4];				r_cell_reg[96] = inform_R[96][4];				r_cell_reg[97] = inform_R[112][4];				r_cell_reg[98] = inform_R[97][4];				r_cell_reg[99] = inform_R[113][4];				r_cell_reg[100] = inform_R[98][4];				r_cell_reg[101] = inform_R[114][4];				r_cell_reg[102] = inform_R[99][4];				r_cell_reg[103] = inform_R[115][4];				r_cell_reg[104] = inform_R[100][4];				r_cell_reg[105] = inform_R[116][4];				r_cell_reg[106] = inform_R[101][4];				r_cell_reg[107] = inform_R[117][4];				r_cell_reg[108] = inform_R[102][4];				r_cell_reg[109] = inform_R[118][4];				r_cell_reg[110] = inform_R[103][4];				r_cell_reg[111] = inform_R[119][4];				r_cell_reg[112] = inform_R[104][4];				r_cell_reg[113] = inform_R[120][4];				r_cell_reg[114] = inform_R[105][4];				r_cell_reg[115] = inform_R[121][4];				r_cell_reg[116] = inform_R[106][4];				r_cell_reg[117] = inform_R[122][4];				r_cell_reg[118] = inform_R[107][4];				r_cell_reg[119] = inform_R[123][4];				r_cell_reg[120] = inform_R[108][4];				r_cell_reg[121] = inform_R[124][4];				r_cell_reg[122] = inform_R[109][4];				r_cell_reg[123] = inform_R[125][4];				r_cell_reg[124] = inform_R[110][4];				r_cell_reg[125] = inform_R[126][4];				r_cell_reg[126] = inform_R[111][4];				r_cell_reg[127] = inform_R[127][4];				r_cell_reg[128] = inform_R[128][4];				r_cell_reg[129] = inform_R[144][4];				r_cell_reg[130] = inform_R[129][4];				r_cell_reg[131] = inform_R[145][4];				r_cell_reg[132] = inform_R[130][4];				r_cell_reg[133] = inform_R[146][4];				r_cell_reg[134] = inform_R[131][4];				r_cell_reg[135] = inform_R[147][4];				r_cell_reg[136] = inform_R[132][4];				r_cell_reg[137] = inform_R[148][4];				r_cell_reg[138] = inform_R[133][4];				r_cell_reg[139] = inform_R[149][4];				r_cell_reg[140] = inform_R[134][4];				r_cell_reg[141] = inform_R[150][4];				r_cell_reg[142] = inform_R[135][4];				r_cell_reg[143] = inform_R[151][4];				r_cell_reg[144] = inform_R[136][4];				r_cell_reg[145] = inform_R[152][4];				r_cell_reg[146] = inform_R[137][4];				r_cell_reg[147] = inform_R[153][4];				r_cell_reg[148] = inform_R[138][4];				r_cell_reg[149] = inform_R[154][4];				r_cell_reg[150] = inform_R[139][4];				r_cell_reg[151] = inform_R[155][4];				r_cell_reg[152] = inform_R[140][4];				r_cell_reg[153] = inform_R[156][4];				r_cell_reg[154] = inform_R[141][4];				r_cell_reg[155] = inform_R[157][4];				r_cell_reg[156] = inform_R[142][4];				r_cell_reg[157] = inform_R[158][4];				r_cell_reg[158] = inform_R[143][4];				r_cell_reg[159] = inform_R[159][4];				r_cell_reg[160] = inform_R[160][4];				r_cell_reg[161] = inform_R[176][4];				r_cell_reg[162] = inform_R[161][4];				r_cell_reg[163] = inform_R[177][4];				r_cell_reg[164] = inform_R[162][4];				r_cell_reg[165] = inform_R[178][4];				r_cell_reg[166] = inform_R[163][4];				r_cell_reg[167] = inform_R[179][4];				r_cell_reg[168] = inform_R[164][4];				r_cell_reg[169] = inform_R[180][4];				r_cell_reg[170] = inform_R[165][4];				r_cell_reg[171] = inform_R[181][4];				r_cell_reg[172] = inform_R[166][4];				r_cell_reg[173] = inform_R[182][4];				r_cell_reg[174] = inform_R[167][4];				r_cell_reg[175] = inform_R[183][4];				r_cell_reg[176] = inform_R[168][4];				r_cell_reg[177] = inform_R[184][4];				r_cell_reg[178] = inform_R[169][4];				r_cell_reg[179] = inform_R[185][4];				r_cell_reg[180] = inform_R[170][4];				r_cell_reg[181] = inform_R[186][4];				r_cell_reg[182] = inform_R[171][4];				r_cell_reg[183] = inform_R[187][4];				r_cell_reg[184] = inform_R[172][4];				r_cell_reg[185] = inform_R[188][4];				r_cell_reg[186] = inform_R[173][4];				r_cell_reg[187] = inform_R[189][4];				r_cell_reg[188] = inform_R[174][4];				r_cell_reg[189] = inform_R[190][4];				r_cell_reg[190] = inform_R[175][4];				r_cell_reg[191] = inform_R[191][4];				r_cell_reg[192] = inform_R[192][4];				r_cell_reg[193] = inform_R[208][4];				r_cell_reg[194] = inform_R[193][4];				r_cell_reg[195] = inform_R[209][4];				r_cell_reg[196] = inform_R[194][4];				r_cell_reg[197] = inform_R[210][4];				r_cell_reg[198] = inform_R[195][4];				r_cell_reg[199] = inform_R[211][4];				r_cell_reg[200] = inform_R[196][4];				r_cell_reg[201] = inform_R[212][4];				r_cell_reg[202] = inform_R[197][4];				r_cell_reg[203] = inform_R[213][4];				r_cell_reg[204] = inform_R[198][4];				r_cell_reg[205] = inform_R[214][4];				r_cell_reg[206] = inform_R[199][4];				r_cell_reg[207] = inform_R[215][4];				r_cell_reg[208] = inform_R[200][4];				r_cell_reg[209] = inform_R[216][4];				r_cell_reg[210] = inform_R[201][4];				r_cell_reg[211] = inform_R[217][4];				r_cell_reg[212] = inform_R[202][4];				r_cell_reg[213] = inform_R[218][4];				r_cell_reg[214] = inform_R[203][4];				r_cell_reg[215] = inform_R[219][4];				r_cell_reg[216] = inform_R[204][4];				r_cell_reg[217] = inform_R[220][4];				r_cell_reg[218] = inform_R[205][4];				r_cell_reg[219] = inform_R[221][4];				r_cell_reg[220] = inform_R[206][4];				r_cell_reg[221] = inform_R[222][4];				r_cell_reg[222] = inform_R[207][4];				r_cell_reg[223] = inform_R[223][4];				r_cell_reg[224] = inform_R[224][4];				r_cell_reg[225] = inform_R[240][4];				r_cell_reg[226] = inform_R[225][4];				r_cell_reg[227] = inform_R[241][4];				r_cell_reg[228] = inform_R[226][4];				r_cell_reg[229] = inform_R[242][4];				r_cell_reg[230] = inform_R[227][4];				r_cell_reg[231] = inform_R[243][4];				r_cell_reg[232] = inform_R[228][4];				r_cell_reg[233] = inform_R[244][4];				r_cell_reg[234] = inform_R[229][4];				r_cell_reg[235] = inform_R[245][4];				r_cell_reg[236] = inform_R[230][4];				r_cell_reg[237] = inform_R[246][4];				r_cell_reg[238] = inform_R[231][4];				r_cell_reg[239] = inform_R[247][4];				r_cell_reg[240] = inform_R[232][4];				r_cell_reg[241] = inform_R[248][4];				r_cell_reg[242] = inform_R[233][4];				r_cell_reg[243] = inform_R[249][4];				r_cell_reg[244] = inform_R[234][4];				r_cell_reg[245] = inform_R[250][4];				r_cell_reg[246] = inform_R[235][4];				r_cell_reg[247] = inform_R[251][4];				r_cell_reg[248] = inform_R[236][4];				r_cell_reg[249] = inform_R[252][4];				r_cell_reg[250] = inform_R[237][4];				r_cell_reg[251] = inform_R[253][4];				r_cell_reg[252] = inform_R[238][4];				r_cell_reg[253] = inform_R[254][4];				r_cell_reg[254] = inform_R[239][4];				r_cell_reg[255] = inform_R[255][4];				l_cell_reg[0] = inform_L[0][5];				l_cell_reg[1] = inform_L[16][5];				l_cell_reg[2] = inform_L[1][5];				l_cell_reg[3] = inform_L[17][5];				l_cell_reg[4] = inform_L[2][5];				l_cell_reg[5] = inform_L[18][5];				l_cell_reg[6] = inform_L[3][5];				l_cell_reg[7] = inform_L[19][5];				l_cell_reg[8] = inform_L[4][5];				l_cell_reg[9] = inform_L[20][5];				l_cell_reg[10] = inform_L[5][5];				l_cell_reg[11] = inform_L[21][5];				l_cell_reg[12] = inform_L[6][5];				l_cell_reg[13] = inform_L[22][5];				l_cell_reg[14] = inform_L[7][5];				l_cell_reg[15] = inform_L[23][5];				l_cell_reg[16] = inform_L[8][5];				l_cell_reg[17] = inform_L[24][5];				l_cell_reg[18] = inform_L[9][5];				l_cell_reg[19] = inform_L[25][5];				l_cell_reg[20] = inform_L[10][5];				l_cell_reg[21] = inform_L[26][5];				l_cell_reg[22] = inform_L[11][5];				l_cell_reg[23] = inform_L[27][5];				l_cell_reg[24] = inform_L[12][5];				l_cell_reg[25] = inform_L[28][5];				l_cell_reg[26] = inform_L[13][5];				l_cell_reg[27] = inform_L[29][5];				l_cell_reg[28] = inform_L[14][5];				l_cell_reg[29] = inform_L[30][5];				l_cell_reg[30] = inform_L[15][5];				l_cell_reg[31] = inform_L[31][5];				l_cell_reg[32] = inform_L[32][5];				l_cell_reg[33] = inform_L[48][5];				l_cell_reg[34] = inform_L[33][5];				l_cell_reg[35] = inform_L[49][5];				l_cell_reg[36] = inform_L[34][5];				l_cell_reg[37] = inform_L[50][5];				l_cell_reg[38] = inform_L[35][5];				l_cell_reg[39] = inform_L[51][5];				l_cell_reg[40] = inform_L[36][5];				l_cell_reg[41] = inform_L[52][5];				l_cell_reg[42] = inform_L[37][5];				l_cell_reg[43] = inform_L[53][5];				l_cell_reg[44] = inform_L[38][5];				l_cell_reg[45] = inform_L[54][5];				l_cell_reg[46] = inform_L[39][5];				l_cell_reg[47] = inform_L[55][5];				l_cell_reg[48] = inform_L[40][5];				l_cell_reg[49] = inform_L[56][5];				l_cell_reg[50] = inform_L[41][5];				l_cell_reg[51] = inform_L[57][5];				l_cell_reg[52] = inform_L[42][5];				l_cell_reg[53] = inform_L[58][5];				l_cell_reg[54] = inform_L[43][5];				l_cell_reg[55] = inform_L[59][5];				l_cell_reg[56] = inform_L[44][5];				l_cell_reg[57] = inform_L[60][5];				l_cell_reg[58] = inform_L[45][5];				l_cell_reg[59] = inform_L[61][5];				l_cell_reg[60] = inform_L[46][5];				l_cell_reg[61] = inform_L[62][5];				l_cell_reg[62] = inform_L[47][5];				l_cell_reg[63] = inform_L[63][5];				l_cell_reg[64] = inform_L[64][5];				l_cell_reg[65] = inform_L[80][5];				l_cell_reg[66] = inform_L[65][5];				l_cell_reg[67] = inform_L[81][5];				l_cell_reg[68] = inform_L[66][5];				l_cell_reg[69] = inform_L[82][5];				l_cell_reg[70] = inform_L[67][5];				l_cell_reg[71] = inform_L[83][5];				l_cell_reg[72] = inform_L[68][5];				l_cell_reg[73] = inform_L[84][5];				l_cell_reg[74] = inform_L[69][5];				l_cell_reg[75] = inform_L[85][5];				l_cell_reg[76] = inform_L[70][5];				l_cell_reg[77] = inform_L[86][5];				l_cell_reg[78] = inform_L[71][5];				l_cell_reg[79] = inform_L[87][5];				l_cell_reg[80] = inform_L[72][5];				l_cell_reg[81] = inform_L[88][5];				l_cell_reg[82] = inform_L[73][5];				l_cell_reg[83] = inform_L[89][5];				l_cell_reg[84] = inform_L[74][5];				l_cell_reg[85] = inform_L[90][5];				l_cell_reg[86] = inform_L[75][5];				l_cell_reg[87] = inform_L[91][5];				l_cell_reg[88] = inform_L[76][5];				l_cell_reg[89] = inform_L[92][5];				l_cell_reg[90] = inform_L[77][5];				l_cell_reg[91] = inform_L[93][5];				l_cell_reg[92] = inform_L[78][5];				l_cell_reg[93] = inform_L[94][5];				l_cell_reg[94] = inform_L[79][5];				l_cell_reg[95] = inform_L[95][5];				l_cell_reg[96] = inform_L[96][5];				l_cell_reg[97] = inform_L[112][5];				l_cell_reg[98] = inform_L[97][5];				l_cell_reg[99] = inform_L[113][5];				l_cell_reg[100] = inform_L[98][5];				l_cell_reg[101] = inform_L[114][5];				l_cell_reg[102] = inform_L[99][5];				l_cell_reg[103] = inform_L[115][5];				l_cell_reg[104] = inform_L[100][5];				l_cell_reg[105] = inform_L[116][5];				l_cell_reg[106] = inform_L[101][5];				l_cell_reg[107] = inform_L[117][5];				l_cell_reg[108] = inform_L[102][5];				l_cell_reg[109] = inform_L[118][5];				l_cell_reg[110] = inform_L[103][5];				l_cell_reg[111] = inform_L[119][5];				l_cell_reg[112] = inform_L[104][5];				l_cell_reg[113] = inform_L[120][5];				l_cell_reg[114] = inform_L[105][5];				l_cell_reg[115] = inform_L[121][5];				l_cell_reg[116] = inform_L[106][5];				l_cell_reg[117] = inform_L[122][5];				l_cell_reg[118] = inform_L[107][5];				l_cell_reg[119] = inform_L[123][5];				l_cell_reg[120] = inform_L[108][5];				l_cell_reg[121] = inform_L[124][5];				l_cell_reg[122] = inform_L[109][5];				l_cell_reg[123] = inform_L[125][5];				l_cell_reg[124] = inform_L[110][5];				l_cell_reg[125] = inform_L[126][5];				l_cell_reg[126] = inform_L[111][5];				l_cell_reg[127] = inform_L[127][5];				l_cell_reg[128] = inform_L[128][5];				l_cell_reg[129] = inform_L[144][5];				l_cell_reg[130] = inform_L[129][5];				l_cell_reg[131] = inform_L[145][5];				l_cell_reg[132] = inform_L[130][5];				l_cell_reg[133] = inform_L[146][5];				l_cell_reg[134] = inform_L[131][5];				l_cell_reg[135] = inform_L[147][5];				l_cell_reg[136] = inform_L[132][5];				l_cell_reg[137] = inform_L[148][5];				l_cell_reg[138] = inform_L[133][5];				l_cell_reg[139] = inform_L[149][5];				l_cell_reg[140] = inform_L[134][5];				l_cell_reg[141] = inform_L[150][5];				l_cell_reg[142] = inform_L[135][5];				l_cell_reg[143] = inform_L[151][5];				l_cell_reg[144] = inform_L[136][5];				l_cell_reg[145] = inform_L[152][5];				l_cell_reg[146] = inform_L[137][5];				l_cell_reg[147] = inform_L[153][5];				l_cell_reg[148] = inform_L[138][5];				l_cell_reg[149] = inform_L[154][5];				l_cell_reg[150] = inform_L[139][5];				l_cell_reg[151] = inform_L[155][5];				l_cell_reg[152] = inform_L[140][5];				l_cell_reg[153] = inform_L[156][5];				l_cell_reg[154] = inform_L[141][5];				l_cell_reg[155] = inform_L[157][5];				l_cell_reg[156] = inform_L[142][5];				l_cell_reg[157] = inform_L[158][5];				l_cell_reg[158] = inform_L[143][5];				l_cell_reg[159] = inform_L[159][5];				l_cell_reg[160] = inform_L[160][5];				l_cell_reg[161] = inform_L[176][5];				l_cell_reg[162] = inform_L[161][5];				l_cell_reg[163] = inform_L[177][5];				l_cell_reg[164] = inform_L[162][5];				l_cell_reg[165] = inform_L[178][5];				l_cell_reg[166] = inform_L[163][5];				l_cell_reg[167] = inform_L[179][5];				l_cell_reg[168] = inform_L[164][5];				l_cell_reg[169] = inform_L[180][5];				l_cell_reg[170] = inform_L[165][5];				l_cell_reg[171] = inform_L[181][5];				l_cell_reg[172] = inform_L[166][5];				l_cell_reg[173] = inform_L[182][5];				l_cell_reg[174] = inform_L[167][5];				l_cell_reg[175] = inform_L[183][5];				l_cell_reg[176] = inform_L[168][5];				l_cell_reg[177] = inform_L[184][5];				l_cell_reg[178] = inform_L[169][5];				l_cell_reg[179] = inform_L[185][5];				l_cell_reg[180] = inform_L[170][5];				l_cell_reg[181] = inform_L[186][5];				l_cell_reg[182] = inform_L[171][5];				l_cell_reg[183] = inform_L[187][5];				l_cell_reg[184] = inform_L[172][5];				l_cell_reg[185] = inform_L[188][5];				l_cell_reg[186] = inform_L[173][5];				l_cell_reg[187] = inform_L[189][5];				l_cell_reg[188] = inform_L[174][5];				l_cell_reg[189] = inform_L[190][5];				l_cell_reg[190] = inform_L[175][5];				l_cell_reg[191] = inform_L[191][5];				l_cell_reg[192] = inform_L[192][5];				l_cell_reg[193] = inform_L[208][5];				l_cell_reg[194] = inform_L[193][5];				l_cell_reg[195] = inform_L[209][5];				l_cell_reg[196] = inform_L[194][5];				l_cell_reg[197] = inform_L[210][5];				l_cell_reg[198] = inform_L[195][5];				l_cell_reg[199] = inform_L[211][5];				l_cell_reg[200] = inform_L[196][5];				l_cell_reg[201] = inform_L[212][5];				l_cell_reg[202] = inform_L[197][5];				l_cell_reg[203] = inform_L[213][5];				l_cell_reg[204] = inform_L[198][5];				l_cell_reg[205] = inform_L[214][5];				l_cell_reg[206] = inform_L[199][5];				l_cell_reg[207] = inform_L[215][5];				l_cell_reg[208] = inform_L[200][5];				l_cell_reg[209] = inform_L[216][5];				l_cell_reg[210] = inform_L[201][5];				l_cell_reg[211] = inform_L[217][5];				l_cell_reg[212] = inform_L[202][5];				l_cell_reg[213] = inform_L[218][5];				l_cell_reg[214] = inform_L[203][5];				l_cell_reg[215] = inform_L[219][5];				l_cell_reg[216] = inform_L[204][5];				l_cell_reg[217] = inform_L[220][5];				l_cell_reg[218] = inform_L[205][5];				l_cell_reg[219] = inform_L[221][5];				l_cell_reg[220] = inform_L[206][5];				l_cell_reg[221] = inform_L[222][5];				l_cell_reg[222] = inform_L[207][5];				l_cell_reg[223] = inform_L[223][5];				l_cell_reg[224] = inform_L[224][5];				l_cell_reg[225] = inform_L[240][5];				l_cell_reg[226] = inform_L[225][5];				l_cell_reg[227] = inform_L[241][5];				l_cell_reg[228] = inform_L[226][5];				l_cell_reg[229] = inform_L[242][5];				l_cell_reg[230] = inform_L[227][5];				l_cell_reg[231] = inform_L[243][5];				l_cell_reg[232] = inform_L[228][5];				l_cell_reg[233] = inform_L[244][5];				l_cell_reg[234] = inform_L[229][5];				l_cell_reg[235] = inform_L[245][5];				l_cell_reg[236] = inform_L[230][5];				l_cell_reg[237] = inform_L[246][5];				l_cell_reg[238] = inform_L[231][5];				l_cell_reg[239] = inform_L[247][5];				l_cell_reg[240] = inform_L[232][5];				l_cell_reg[241] = inform_L[248][5];				l_cell_reg[242] = inform_L[233][5];				l_cell_reg[243] = inform_L[249][5];				l_cell_reg[244] = inform_L[234][5];				l_cell_reg[245] = inform_L[250][5];				l_cell_reg[246] = inform_L[235][5];				l_cell_reg[247] = inform_L[251][5];				l_cell_reg[248] = inform_L[236][5];				l_cell_reg[249] = inform_L[252][5];				l_cell_reg[250] = inform_L[237][5];				l_cell_reg[251] = inform_L[253][5];				l_cell_reg[252] = inform_L[238][5];				l_cell_reg[253] = inform_L[254][5];				l_cell_reg[254] = inform_L[239][5];				l_cell_reg[255] = inform_L[255][5];			end
			6:			begin				r_cell_reg[0] = inform_R[0][5];				r_cell_reg[1] = inform_R[32][5];				r_cell_reg[2] = inform_R[1][5];				r_cell_reg[3] = inform_R[33][5];				r_cell_reg[4] = inform_R[2][5];				r_cell_reg[5] = inform_R[34][5];				r_cell_reg[6] = inform_R[3][5];				r_cell_reg[7] = inform_R[35][5];				r_cell_reg[8] = inform_R[4][5];				r_cell_reg[9] = inform_R[36][5];				r_cell_reg[10] = inform_R[5][5];				r_cell_reg[11] = inform_R[37][5];				r_cell_reg[12] = inform_R[6][5];				r_cell_reg[13] = inform_R[38][5];				r_cell_reg[14] = inform_R[7][5];				r_cell_reg[15] = inform_R[39][5];				r_cell_reg[16] = inform_R[8][5];				r_cell_reg[17] = inform_R[40][5];				r_cell_reg[18] = inform_R[9][5];				r_cell_reg[19] = inform_R[41][5];				r_cell_reg[20] = inform_R[10][5];				r_cell_reg[21] = inform_R[42][5];				r_cell_reg[22] = inform_R[11][5];				r_cell_reg[23] = inform_R[43][5];				r_cell_reg[24] = inform_R[12][5];				r_cell_reg[25] = inform_R[44][5];				r_cell_reg[26] = inform_R[13][5];				r_cell_reg[27] = inform_R[45][5];				r_cell_reg[28] = inform_R[14][5];				r_cell_reg[29] = inform_R[46][5];				r_cell_reg[30] = inform_R[15][5];				r_cell_reg[31] = inform_R[47][5];				r_cell_reg[32] = inform_R[16][5];				r_cell_reg[33] = inform_R[48][5];				r_cell_reg[34] = inform_R[17][5];				r_cell_reg[35] = inform_R[49][5];				r_cell_reg[36] = inform_R[18][5];				r_cell_reg[37] = inform_R[50][5];				r_cell_reg[38] = inform_R[19][5];				r_cell_reg[39] = inform_R[51][5];				r_cell_reg[40] = inform_R[20][5];				r_cell_reg[41] = inform_R[52][5];				r_cell_reg[42] = inform_R[21][5];				r_cell_reg[43] = inform_R[53][5];				r_cell_reg[44] = inform_R[22][5];				r_cell_reg[45] = inform_R[54][5];				r_cell_reg[46] = inform_R[23][5];				r_cell_reg[47] = inform_R[55][5];				r_cell_reg[48] = inform_R[24][5];				r_cell_reg[49] = inform_R[56][5];				r_cell_reg[50] = inform_R[25][5];				r_cell_reg[51] = inform_R[57][5];				r_cell_reg[52] = inform_R[26][5];				r_cell_reg[53] = inform_R[58][5];				r_cell_reg[54] = inform_R[27][5];				r_cell_reg[55] = inform_R[59][5];				r_cell_reg[56] = inform_R[28][5];				r_cell_reg[57] = inform_R[60][5];				r_cell_reg[58] = inform_R[29][5];				r_cell_reg[59] = inform_R[61][5];				r_cell_reg[60] = inform_R[30][5];				r_cell_reg[61] = inform_R[62][5];				r_cell_reg[62] = inform_R[31][5];				r_cell_reg[63] = inform_R[63][5];				r_cell_reg[64] = inform_R[64][5];				r_cell_reg[65] = inform_R[96][5];				r_cell_reg[66] = inform_R[65][5];				r_cell_reg[67] = inform_R[97][5];				r_cell_reg[68] = inform_R[66][5];				r_cell_reg[69] = inform_R[98][5];				r_cell_reg[70] = inform_R[67][5];				r_cell_reg[71] = inform_R[99][5];				r_cell_reg[72] = inform_R[68][5];				r_cell_reg[73] = inform_R[100][5];				r_cell_reg[74] = inform_R[69][5];				r_cell_reg[75] = inform_R[101][5];				r_cell_reg[76] = inform_R[70][5];				r_cell_reg[77] = inform_R[102][5];				r_cell_reg[78] = inform_R[71][5];				r_cell_reg[79] = inform_R[103][5];				r_cell_reg[80] = inform_R[72][5];				r_cell_reg[81] = inform_R[104][5];				r_cell_reg[82] = inform_R[73][5];				r_cell_reg[83] = inform_R[105][5];				r_cell_reg[84] = inform_R[74][5];				r_cell_reg[85] = inform_R[106][5];				r_cell_reg[86] = inform_R[75][5];				r_cell_reg[87] = inform_R[107][5];				r_cell_reg[88] = inform_R[76][5];				r_cell_reg[89] = inform_R[108][5];				r_cell_reg[90] = inform_R[77][5];				r_cell_reg[91] = inform_R[109][5];				r_cell_reg[92] = inform_R[78][5];				r_cell_reg[93] = inform_R[110][5];				r_cell_reg[94] = inform_R[79][5];				r_cell_reg[95] = inform_R[111][5];				r_cell_reg[96] = inform_R[80][5];				r_cell_reg[97] = inform_R[112][5];				r_cell_reg[98] = inform_R[81][5];				r_cell_reg[99] = inform_R[113][5];				r_cell_reg[100] = inform_R[82][5];				r_cell_reg[101] = inform_R[114][5];				r_cell_reg[102] = inform_R[83][5];				r_cell_reg[103] = inform_R[115][5];				r_cell_reg[104] = inform_R[84][5];				r_cell_reg[105] = inform_R[116][5];				r_cell_reg[106] = inform_R[85][5];				r_cell_reg[107] = inform_R[117][5];				r_cell_reg[108] = inform_R[86][5];				r_cell_reg[109] = inform_R[118][5];				r_cell_reg[110] = inform_R[87][5];				r_cell_reg[111] = inform_R[119][5];				r_cell_reg[112] = inform_R[88][5];				r_cell_reg[113] = inform_R[120][5];				r_cell_reg[114] = inform_R[89][5];				r_cell_reg[115] = inform_R[121][5];				r_cell_reg[116] = inform_R[90][5];				r_cell_reg[117] = inform_R[122][5];				r_cell_reg[118] = inform_R[91][5];				r_cell_reg[119] = inform_R[123][5];				r_cell_reg[120] = inform_R[92][5];				r_cell_reg[121] = inform_R[124][5];				r_cell_reg[122] = inform_R[93][5];				r_cell_reg[123] = inform_R[125][5];				r_cell_reg[124] = inform_R[94][5];				r_cell_reg[125] = inform_R[126][5];				r_cell_reg[126] = inform_R[95][5];				r_cell_reg[127] = inform_R[127][5];				r_cell_reg[128] = inform_R[128][5];				r_cell_reg[129] = inform_R[160][5];				r_cell_reg[130] = inform_R[129][5];				r_cell_reg[131] = inform_R[161][5];				r_cell_reg[132] = inform_R[130][5];				r_cell_reg[133] = inform_R[162][5];				r_cell_reg[134] = inform_R[131][5];				r_cell_reg[135] = inform_R[163][5];				r_cell_reg[136] = inform_R[132][5];				r_cell_reg[137] = inform_R[164][5];				r_cell_reg[138] = inform_R[133][5];				r_cell_reg[139] = inform_R[165][5];				r_cell_reg[140] = inform_R[134][5];				r_cell_reg[141] = inform_R[166][5];				r_cell_reg[142] = inform_R[135][5];				r_cell_reg[143] = inform_R[167][5];				r_cell_reg[144] = inform_R[136][5];				r_cell_reg[145] = inform_R[168][5];				r_cell_reg[146] = inform_R[137][5];				r_cell_reg[147] = inform_R[169][5];				r_cell_reg[148] = inform_R[138][5];				r_cell_reg[149] = inform_R[170][5];				r_cell_reg[150] = inform_R[139][5];				r_cell_reg[151] = inform_R[171][5];				r_cell_reg[152] = inform_R[140][5];				r_cell_reg[153] = inform_R[172][5];				r_cell_reg[154] = inform_R[141][5];				r_cell_reg[155] = inform_R[173][5];				r_cell_reg[156] = inform_R[142][5];				r_cell_reg[157] = inform_R[174][5];				r_cell_reg[158] = inform_R[143][5];				r_cell_reg[159] = inform_R[175][5];				r_cell_reg[160] = inform_R[144][5];				r_cell_reg[161] = inform_R[176][5];				r_cell_reg[162] = inform_R[145][5];				r_cell_reg[163] = inform_R[177][5];				r_cell_reg[164] = inform_R[146][5];				r_cell_reg[165] = inform_R[178][5];				r_cell_reg[166] = inform_R[147][5];				r_cell_reg[167] = inform_R[179][5];				r_cell_reg[168] = inform_R[148][5];				r_cell_reg[169] = inform_R[180][5];				r_cell_reg[170] = inform_R[149][5];				r_cell_reg[171] = inform_R[181][5];				r_cell_reg[172] = inform_R[150][5];				r_cell_reg[173] = inform_R[182][5];				r_cell_reg[174] = inform_R[151][5];				r_cell_reg[175] = inform_R[183][5];				r_cell_reg[176] = inform_R[152][5];				r_cell_reg[177] = inform_R[184][5];				r_cell_reg[178] = inform_R[153][5];				r_cell_reg[179] = inform_R[185][5];				r_cell_reg[180] = inform_R[154][5];				r_cell_reg[181] = inform_R[186][5];				r_cell_reg[182] = inform_R[155][5];				r_cell_reg[183] = inform_R[187][5];				r_cell_reg[184] = inform_R[156][5];				r_cell_reg[185] = inform_R[188][5];				r_cell_reg[186] = inform_R[157][5];				r_cell_reg[187] = inform_R[189][5];				r_cell_reg[188] = inform_R[158][5];				r_cell_reg[189] = inform_R[190][5];				r_cell_reg[190] = inform_R[159][5];				r_cell_reg[191] = inform_R[191][5];				r_cell_reg[192] = inform_R[192][5];				r_cell_reg[193] = inform_R[224][5];				r_cell_reg[194] = inform_R[193][5];				r_cell_reg[195] = inform_R[225][5];				r_cell_reg[196] = inform_R[194][5];				r_cell_reg[197] = inform_R[226][5];				r_cell_reg[198] = inform_R[195][5];				r_cell_reg[199] = inform_R[227][5];				r_cell_reg[200] = inform_R[196][5];				r_cell_reg[201] = inform_R[228][5];				r_cell_reg[202] = inform_R[197][5];				r_cell_reg[203] = inform_R[229][5];				r_cell_reg[204] = inform_R[198][5];				r_cell_reg[205] = inform_R[230][5];				r_cell_reg[206] = inform_R[199][5];				r_cell_reg[207] = inform_R[231][5];				r_cell_reg[208] = inform_R[200][5];				r_cell_reg[209] = inform_R[232][5];				r_cell_reg[210] = inform_R[201][5];				r_cell_reg[211] = inform_R[233][5];				r_cell_reg[212] = inform_R[202][5];				r_cell_reg[213] = inform_R[234][5];				r_cell_reg[214] = inform_R[203][5];				r_cell_reg[215] = inform_R[235][5];				r_cell_reg[216] = inform_R[204][5];				r_cell_reg[217] = inform_R[236][5];				r_cell_reg[218] = inform_R[205][5];				r_cell_reg[219] = inform_R[237][5];				r_cell_reg[220] = inform_R[206][5];				r_cell_reg[221] = inform_R[238][5];				r_cell_reg[222] = inform_R[207][5];				r_cell_reg[223] = inform_R[239][5];				r_cell_reg[224] = inform_R[208][5];				r_cell_reg[225] = inform_R[240][5];				r_cell_reg[226] = inform_R[209][5];				r_cell_reg[227] = inform_R[241][5];				r_cell_reg[228] = inform_R[210][5];				r_cell_reg[229] = inform_R[242][5];				r_cell_reg[230] = inform_R[211][5];				r_cell_reg[231] = inform_R[243][5];				r_cell_reg[232] = inform_R[212][5];				r_cell_reg[233] = inform_R[244][5];				r_cell_reg[234] = inform_R[213][5];				r_cell_reg[235] = inform_R[245][5];				r_cell_reg[236] = inform_R[214][5];				r_cell_reg[237] = inform_R[246][5];				r_cell_reg[238] = inform_R[215][5];				r_cell_reg[239] = inform_R[247][5];				r_cell_reg[240] = inform_R[216][5];				r_cell_reg[241] = inform_R[248][5];				r_cell_reg[242] = inform_R[217][5];				r_cell_reg[243] = inform_R[249][5];				r_cell_reg[244] = inform_R[218][5];				r_cell_reg[245] = inform_R[250][5];				r_cell_reg[246] = inform_R[219][5];				r_cell_reg[247] = inform_R[251][5];				r_cell_reg[248] = inform_R[220][5];				r_cell_reg[249] = inform_R[252][5];				r_cell_reg[250] = inform_R[221][5];				r_cell_reg[251] = inform_R[253][5];				r_cell_reg[252] = inform_R[222][5];				r_cell_reg[253] = inform_R[254][5];				r_cell_reg[254] = inform_R[223][5];				r_cell_reg[255] = inform_R[255][5];				l_cell_reg[0] = inform_L[0][6];				l_cell_reg[1] = inform_L[32][6];				l_cell_reg[2] = inform_L[1][6];				l_cell_reg[3] = inform_L[33][6];				l_cell_reg[4] = inform_L[2][6];				l_cell_reg[5] = inform_L[34][6];				l_cell_reg[6] = inform_L[3][6];				l_cell_reg[7] = inform_L[35][6];				l_cell_reg[8] = inform_L[4][6];				l_cell_reg[9] = inform_L[36][6];				l_cell_reg[10] = inform_L[5][6];				l_cell_reg[11] = inform_L[37][6];				l_cell_reg[12] = inform_L[6][6];				l_cell_reg[13] = inform_L[38][6];				l_cell_reg[14] = inform_L[7][6];				l_cell_reg[15] = inform_L[39][6];				l_cell_reg[16] = inform_L[8][6];				l_cell_reg[17] = inform_L[40][6];				l_cell_reg[18] = inform_L[9][6];				l_cell_reg[19] = inform_L[41][6];				l_cell_reg[20] = inform_L[10][6];				l_cell_reg[21] = inform_L[42][6];				l_cell_reg[22] = inform_L[11][6];				l_cell_reg[23] = inform_L[43][6];				l_cell_reg[24] = inform_L[12][6];				l_cell_reg[25] = inform_L[44][6];				l_cell_reg[26] = inform_L[13][6];				l_cell_reg[27] = inform_L[45][6];				l_cell_reg[28] = inform_L[14][6];				l_cell_reg[29] = inform_L[46][6];				l_cell_reg[30] = inform_L[15][6];				l_cell_reg[31] = inform_L[47][6];				l_cell_reg[32] = inform_L[16][6];				l_cell_reg[33] = inform_L[48][6];				l_cell_reg[34] = inform_L[17][6];				l_cell_reg[35] = inform_L[49][6];				l_cell_reg[36] = inform_L[18][6];				l_cell_reg[37] = inform_L[50][6];				l_cell_reg[38] = inform_L[19][6];				l_cell_reg[39] = inform_L[51][6];				l_cell_reg[40] = inform_L[20][6];				l_cell_reg[41] = inform_L[52][6];				l_cell_reg[42] = inform_L[21][6];				l_cell_reg[43] = inform_L[53][6];				l_cell_reg[44] = inform_L[22][6];				l_cell_reg[45] = inform_L[54][6];				l_cell_reg[46] = inform_L[23][6];				l_cell_reg[47] = inform_L[55][6];				l_cell_reg[48] = inform_L[24][6];				l_cell_reg[49] = inform_L[56][6];				l_cell_reg[50] = inform_L[25][6];				l_cell_reg[51] = inform_L[57][6];				l_cell_reg[52] = inform_L[26][6];				l_cell_reg[53] = inform_L[58][6];				l_cell_reg[54] = inform_L[27][6];				l_cell_reg[55] = inform_L[59][6];				l_cell_reg[56] = inform_L[28][6];				l_cell_reg[57] = inform_L[60][6];				l_cell_reg[58] = inform_L[29][6];				l_cell_reg[59] = inform_L[61][6];				l_cell_reg[60] = inform_L[30][6];				l_cell_reg[61] = inform_L[62][6];				l_cell_reg[62] = inform_L[31][6];				l_cell_reg[63] = inform_L[63][6];				l_cell_reg[64] = inform_L[64][6];				l_cell_reg[65] = inform_L[96][6];				l_cell_reg[66] = inform_L[65][6];				l_cell_reg[67] = inform_L[97][6];				l_cell_reg[68] = inform_L[66][6];				l_cell_reg[69] = inform_L[98][6];				l_cell_reg[70] = inform_L[67][6];				l_cell_reg[71] = inform_L[99][6];				l_cell_reg[72] = inform_L[68][6];				l_cell_reg[73] = inform_L[100][6];				l_cell_reg[74] = inform_L[69][6];				l_cell_reg[75] = inform_L[101][6];				l_cell_reg[76] = inform_L[70][6];				l_cell_reg[77] = inform_L[102][6];				l_cell_reg[78] = inform_L[71][6];				l_cell_reg[79] = inform_L[103][6];				l_cell_reg[80] = inform_L[72][6];				l_cell_reg[81] = inform_L[104][6];				l_cell_reg[82] = inform_L[73][6];				l_cell_reg[83] = inform_L[105][6];				l_cell_reg[84] = inform_L[74][6];				l_cell_reg[85] = inform_L[106][6];				l_cell_reg[86] = inform_L[75][6];				l_cell_reg[87] = inform_L[107][6];				l_cell_reg[88] = inform_L[76][6];				l_cell_reg[89] = inform_L[108][6];				l_cell_reg[90] = inform_L[77][6];				l_cell_reg[91] = inform_L[109][6];				l_cell_reg[92] = inform_L[78][6];				l_cell_reg[93] = inform_L[110][6];				l_cell_reg[94] = inform_L[79][6];				l_cell_reg[95] = inform_L[111][6];				l_cell_reg[96] = inform_L[80][6];				l_cell_reg[97] = inform_L[112][6];				l_cell_reg[98] = inform_L[81][6];				l_cell_reg[99] = inform_L[113][6];				l_cell_reg[100] = inform_L[82][6];				l_cell_reg[101] = inform_L[114][6];				l_cell_reg[102] = inform_L[83][6];				l_cell_reg[103] = inform_L[115][6];				l_cell_reg[104] = inform_L[84][6];				l_cell_reg[105] = inform_L[116][6];				l_cell_reg[106] = inform_L[85][6];				l_cell_reg[107] = inform_L[117][6];				l_cell_reg[108] = inform_L[86][6];				l_cell_reg[109] = inform_L[118][6];				l_cell_reg[110] = inform_L[87][6];				l_cell_reg[111] = inform_L[119][6];				l_cell_reg[112] = inform_L[88][6];				l_cell_reg[113] = inform_L[120][6];				l_cell_reg[114] = inform_L[89][6];				l_cell_reg[115] = inform_L[121][6];				l_cell_reg[116] = inform_L[90][6];				l_cell_reg[117] = inform_L[122][6];				l_cell_reg[118] = inform_L[91][6];				l_cell_reg[119] = inform_L[123][6];				l_cell_reg[120] = inform_L[92][6];				l_cell_reg[121] = inform_L[124][6];				l_cell_reg[122] = inform_L[93][6];				l_cell_reg[123] = inform_L[125][6];				l_cell_reg[124] = inform_L[94][6];				l_cell_reg[125] = inform_L[126][6];				l_cell_reg[126] = inform_L[95][6];				l_cell_reg[127] = inform_L[127][6];				l_cell_reg[128] = inform_L[128][6];				l_cell_reg[129] = inform_L[160][6];				l_cell_reg[130] = inform_L[129][6];				l_cell_reg[131] = inform_L[161][6];				l_cell_reg[132] = inform_L[130][6];				l_cell_reg[133] = inform_L[162][6];				l_cell_reg[134] = inform_L[131][6];				l_cell_reg[135] = inform_L[163][6];				l_cell_reg[136] = inform_L[132][6];				l_cell_reg[137] = inform_L[164][6];				l_cell_reg[138] = inform_L[133][6];				l_cell_reg[139] = inform_L[165][6];				l_cell_reg[140] = inform_L[134][6];				l_cell_reg[141] = inform_L[166][6];				l_cell_reg[142] = inform_L[135][6];				l_cell_reg[143] = inform_L[167][6];				l_cell_reg[144] = inform_L[136][6];				l_cell_reg[145] = inform_L[168][6];				l_cell_reg[146] = inform_L[137][6];				l_cell_reg[147] = inform_L[169][6];				l_cell_reg[148] = inform_L[138][6];				l_cell_reg[149] = inform_L[170][6];				l_cell_reg[150] = inform_L[139][6];				l_cell_reg[151] = inform_L[171][6];				l_cell_reg[152] = inform_L[140][6];				l_cell_reg[153] = inform_L[172][6];				l_cell_reg[154] = inform_L[141][6];				l_cell_reg[155] = inform_L[173][6];				l_cell_reg[156] = inform_L[142][6];				l_cell_reg[157] = inform_L[174][6];				l_cell_reg[158] = inform_L[143][6];				l_cell_reg[159] = inform_L[175][6];				l_cell_reg[160] = inform_L[144][6];				l_cell_reg[161] = inform_L[176][6];				l_cell_reg[162] = inform_L[145][6];				l_cell_reg[163] = inform_L[177][6];				l_cell_reg[164] = inform_L[146][6];				l_cell_reg[165] = inform_L[178][6];				l_cell_reg[166] = inform_L[147][6];				l_cell_reg[167] = inform_L[179][6];				l_cell_reg[168] = inform_L[148][6];				l_cell_reg[169] = inform_L[180][6];				l_cell_reg[170] = inform_L[149][6];				l_cell_reg[171] = inform_L[181][6];				l_cell_reg[172] = inform_L[150][6];				l_cell_reg[173] = inform_L[182][6];				l_cell_reg[174] = inform_L[151][6];				l_cell_reg[175] = inform_L[183][6];				l_cell_reg[176] = inform_L[152][6];				l_cell_reg[177] = inform_L[184][6];				l_cell_reg[178] = inform_L[153][6];				l_cell_reg[179] = inform_L[185][6];				l_cell_reg[180] = inform_L[154][6];				l_cell_reg[181] = inform_L[186][6];				l_cell_reg[182] = inform_L[155][6];				l_cell_reg[183] = inform_L[187][6];				l_cell_reg[184] = inform_L[156][6];				l_cell_reg[185] = inform_L[188][6];				l_cell_reg[186] = inform_L[157][6];				l_cell_reg[187] = inform_L[189][6];				l_cell_reg[188] = inform_L[158][6];				l_cell_reg[189] = inform_L[190][6];				l_cell_reg[190] = inform_L[159][6];				l_cell_reg[191] = inform_L[191][6];				l_cell_reg[192] = inform_L[192][6];				l_cell_reg[193] = inform_L[224][6];				l_cell_reg[194] = inform_L[193][6];				l_cell_reg[195] = inform_L[225][6];				l_cell_reg[196] = inform_L[194][6];				l_cell_reg[197] = inform_L[226][6];				l_cell_reg[198] = inform_L[195][6];				l_cell_reg[199] = inform_L[227][6];				l_cell_reg[200] = inform_L[196][6];				l_cell_reg[201] = inform_L[228][6];				l_cell_reg[202] = inform_L[197][6];				l_cell_reg[203] = inform_L[229][6];				l_cell_reg[204] = inform_L[198][6];				l_cell_reg[205] = inform_L[230][6];				l_cell_reg[206] = inform_L[199][6];				l_cell_reg[207] = inform_L[231][6];				l_cell_reg[208] = inform_L[200][6];				l_cell_reg[209] = inform_L[232][6];				l_cell_reg[210] = inform_L[201][6];				l_cell_reg[211] = inform_L[233][6];				l_cell_reg[212] = inform_L[202][6];				l_cell_reg[213] = inform_L[234][6];				l_cell_reg[214] = inform_L[203][6];				l_cell_reg[215] = inform_L[235][6];				l_cell_reg[216] = inform_L[204][6];				l_cell_reg[217] = inform_L[236][6];				l_cell_reg[218] = inform_L[205][6];				l_cell_reg[219] = inform_L[237][6];				l_cell_reg[220] = inform_L[206][6];				l_cell_reg[221] = inform_L[238][6];				l_cell_reg[222] = inform_L[207][6];				l_cell_reg[223] = inform_L[239][6];				l_cell_reg[224] = inform_L[208][6];				l_cell_reg[225] = inform_L[240][6];				l_cell_reg[226] = inform_L[209][6];				l_cell_reg[227] = inform_L[241][6];				l_cell_reg[228] = inform_L[210][6];				l_cell_reg[229] = inform_L[242][6];				l_cell_reg[230] = inform_L[211][6];				l_cell_reg[231] = inform_L[243][6];				l_cell_reg[232] = inform_L[212][6];				l_cell_reg[233] = inform_L[244][6];				l_cell_reg[234] = inform_L[213][6];				l_cell_reg[235] = inform_L[245][6];				l_cell_reg[236] = inform_L[214][6];				l_cell_reg[237] = inform_L[246][6];				l_cell_reg[238] = inform_L[215][6];				l_cell_reg[239] = inform_L[247][6];				l_cell_reg[240] = inform_L[216][6];				l_cell_reg[241] = inform_L[248][6];				l_cell_reg[242] = inform_L[217][6];				l_cell_reg[243] = inform_L[249][6];				l_cell_reg[244] = inform_L[218][6];				l_cell_reg[245] = inform_L[250][6];				l_cell_reg[246] = inform_L[219][6];				l_cell_reg[247] = inform_L[251][6];				l_cell_reg[248] = inform_L[220][6];				l_cell_reg[249] = inform_L[252][6];				l_cell_reg[250] = inform_L[221][6];				l_cell_reg[251] = inform_L[253][6];				l_cell_reg[252] = inform_L[222][6];				l_cell_reg[253] = inform_L[254][6];				l_cell_reg[254] = inform_L[223][6];				l_cell_reg[255] = inform_L[255][6];			end
			7:			begin				r_cell_reg[0] = inform_R[0][6];				r_cell_reg[1] = inform_R[64][6];				r_cell_reg[2] = inform_R[1][6];				r_cell_reg[3] = inform_R[65][6];				r_cell_reg[4] = inform_R[2][6];				r_cell_reg[5] = inform_R[66][6];				r_cell_reg[6] = inform_R[3][6];				r_cell_reg[7] = inform_R[67][6];				r_cell_reg[8] = inform_R[4][6];				r_cell_reg[9] = inform_R[68][6];				r_cell_reg[10] = inform_R[5][6];				r_cell_reg[11] = inform_R[69][6];				r_cell_reg[12] = inform_R[6][6];				r_cell_reg[13] = inform_R[70][6];				r_cell_reg[14] = inform_R[7][6];				r_cell_reg[15] = inform_R[71][6];				r_cell_reg[16] = inform_R[8][6];				r_cell_reg[17] = inform_R[72][6];				r_cell_reg[18] = inform_R[9][6];				r_cell_reg[19] = inform_R[73][6];				r_cell_reg[20] = inform_R[10][6];				r_cell_reg[21] = inform_R[74][6];				r_cell_reg[22] = inform_R[11][6];				r_cell_reg[23] = inform_R[75][6];				r_cell_reg[24] = inform_R[12][6];				r_cell_reg[25] = inform_R[76][6];				r_cell_reg[26] = inform_R[13][6];				r_cell_reg[27] = inform_R[77][6];				r_cell_reg[28] = inform_R[14][6];				r_cell_reg[29] = inform_R[78][6];				r_cell_reg[30] = inform_R[15][6];				r_cell_reg[31] = inform_R[79][6];				r_cell_reg[32] = inform_R[16][6];				r_cell_reg[33] = inform_R[80][6];				r_cell_reg[34] = inform_R[17][6];				r_cell_reg[35] = inform_R[81][6];				r_cell_reg[36] = inform_R[18][6];				r_cell_reg[37] = inform_R[82][6];				r_cell_reg[38] = inform_R[19][6];				r_cell_reg[39] = inform_R[83][6];				r_cell_reg[40] = inform_R[20][6];				r_cell_reg[41] = inform_R[84][6];				r_cell_reg[42] = inform_R[21][6];				r_cell_reg[43] = inform_R[85][6];				r_cell_reg[44] = inform_R[22][6];				r_cell_reg[45] = inform_R[86][6];				r_cell_reg[46] = inform_R[23][6];				r_cell_reg[47] = inform_R[87][6];				r_cell_reg[48] = inform_R[24][6];				r_cell_reg[49] = inform_R[88][6];				r_cell_reg[50] = inform_R[25][6];				r_cell_reg[51] = inform_R[89][6];				r_cell_reg[52] = inform_R[26][6];				r_cell_reg[53] = inform_R[90][6];				r_cell_reg[54] = inform_R[27][6];				r_cell_reg[55] = inform_R[91][6];				r_cell_reg[56] = inform_R[28][6];				r_cell_reg[57] = inform_R[92][6];				r_cell_reg[58] = inform_R[29][6];				r_cell_reg[59] = inform_R[93][6];				r_cell_reg[60] = inform_R[30][6];				r_cell_reg[61] = inform_R[94][6];				r_cell_reg[62] = inform_R[31][6];				r_cell_reg[63] = inform_R[95][6];				r_cell_reg[64] = inform_R[32][6];				r_cell_reg[65] = inform_R[96][6];				r_cell_reg[66] = inform_R[33][6];				r_cell_reg[67] = inform_R[97][6];				r_cell_reg[68] = inform_R[34][6];				r_cell_reg[69] = inform_R[98][6];				r_cell_reg[70] = inform_R[35][6];				r_cell_reg[71] = inform_R[99][6];				r_cell_reg[72] = inform_R[36][6];				r_cell_reg[73] = inform_R[100][6];				r_cell_reg[74] = inform_R[37][6];				r_cell_reg[75] = inform_R[101][6];				r_cell_reg[76] = inform_R[38][6];				r_cell_reg[77] = inform_R[102][6];				r_cell_reg[78] = inform_R[39][6];				r_cell_reg[79] = inform_R[103][6];				r_cell_reg[80] = inform_R[40][6];				r_cell_reg[81] = inform_R[104][6];				r_cell_reg[82] = inform_R[41][6];				r_cell_reg[83] = inform_R[105][6];				r_cell_reg[84] = inform_R[42][6];				r_cell_reg[85] = inform_R[106][6];				r_cell_reg[86] = inform_R[43][6];				r_cell_reg[87] = inform_R[107][6];				r_cell_reg[88] = inform_R[44][6];				r_cell_reg[89] = inform_R[108][6];				r_cell_reg[90] = inform_R[45][6];				r_cell_reg[91] = inform_R[109][6];				r_cell_reg[92] = inform_R[46][6];				r_cell_reg[93] = inform_R[110][6];				r_cell_reg[94] = inform_R[47][6];				r_cell_reg[95] = inform_R[111][6];				r_cell_reg[96] = inform_R[48][6];				r_cell_reg[97] = inform_R[112][6];				r_cell_reg[98] = inform_R[49][6];				r_cell_reg[99] = inform_R[113][6];				r_cell_reg[100] = inform_R[50][6];				r_cell_reg[101] = inform_R[114][6];				r_cell_reg[102] = inform_R[51][6];				r_cell_reg[103] = inform_R[115][6];				r_cell_reg[104] = inform_R[52][6];				r_cell_reg[105] = inform_R[116][6];				r_cell_reg[106] = inform_R[53][6];				r_cell_reg[107] = inform_R[117][6];				r_cell_reg[108] = inform_R[54][6];				r_cell_reg[109] = inform_R[118][6];				r_cell_reg[110] = inform_R[55][6];				r_cell_reg[111] = inform_R[119][6];				r_cell_reg[112] = inform_R[56][6];				r_cell_reg[113] = inform_R[120][6];				r_cell_reg[114] = inform_R[57][6];				r_cell_reg[115] = inform_R[121][6];				r_cell_reg[116] = inform_R[58][6];				r_cell_reg[117] = inform_R[122][6];				r_cell_reg[118] = inform_R[59][6];				r_cell_reg[119] = inform_R[123][6];				r_cell_reg[120] = inform_R[60][6];				r_cell_reg[121] = inform_R[124][6];				r_cell_reg[122] = inform_R[61][6];				r_cell_reg[123] = inform_R[125][6];				r_cell_reg[124] = inform_R[62][6];				r_cell_reg[125] = inform_R[126][6];				r_cell_reg[126] = inform_R[63][6];				r_cell_reg[127] = inform_R[127][6];				r_cell_reg[128] = inform_R[128][6];				r_cell_reg[129] = inform_R[192][6];				r_cell_reg[130] = inform_R[129][6];				r_cell_reg[131] = inform_R[193][6];				r_cell_reg[132] = inform_R[130][6];				r_cell_reg[133] = inform_R[194][6];				r_cell_reg[134] = inform_R[131][6];				r_cell_reg[135] = inform_R[195][6];				r_cell_reg[136] = inform_R[132][6];				r_cell_reg[137] = inform_R[196][6];				r_cell_reg[138] = inform_R[133][6];				r_cell_reg[139] = inform_R[197][6];				r_cell_reg[140] = inform_R[134][6];				r_cell_reg[141] = inform_R[198][6];				r_cell_reg[142] = inform_R[135][6];				r_cell_reg[143] = inform_R[199][6];				r_cell_reg[144] = inform_R[136][6];				r_cell_reg[145] = inform_R[200][6];				r_cell_reg[146] = inform_R[137][6];				r_cell_reg[147] = inform_R[201][6];				r_cell_reg[148] = inform_R[138][6];				r_cell_reg[149] = inform_R[202][6];				r_cell_reg[150] = inform_R[139][6];				r_cell_reg[151] = inform_R[203][6];				r_cell_reg[152] = inform_R[140][6];				r_cell_reg[153] = inform_R[204][6];				r_cell_reg[154] = inform_R[141][6];				r_cell_reg[155] = inform_R[205][6];				r_cell_reg[156] = inform_R[142][6];				r_cell_reg[157] = inform_R[206][6];				r_cell_reg[158] = inform_R[143][6];				r_cell_reg[159] = inform_R[207][6];				r_cell_reg[160] = inform_R[144][6];				r_cell_reg[161] = inform_R[208][6];				r_cell_reg[162] = inform_R[145][6];				r_cell_reg[163] = inform_R[209][6];				r_cell_reg[164] = inform_R[146][6];				r_cell_reg[165] = inform_R[210][6];				r_cell_reg[166] = inform_R[147][6];				r_cell_reg[167] = inform_R[211][6];				r_cell_reg[168] = inform_R[148][6];				r_cell_reg[169] = inform_R[212][6];				r_cell_reg[170] = inform_R[149][6];				r_cell_reg[171] = inform_R[213][6];				r_cell_reg[172] = inform_R[150][6];				r_cell_reg[173] = inform_R[214][6];				r_cell_reg[174] = inform_R[151][6];				r_cell_reg[175] = inform_R[215][6];				r_cell_reg[176] = inform_R[152][6];				r_cell_reg[177] = inform_R[216][6];				r_cell_reg[178] = inform_R[153][6];				r_cell_reg[179] = inform_R[217][6];				r_cell_reg[180] = inform_R[154][6];				r_cell_reg[181] = inform_R[218][6];				r_cell_reg[182] = inform_R[155][6];				r_cell_reg[183] = inform_R[219][6];				r_cell_reg[184] = inform_R[156][6];				r_cell_reg[185] = inform_R[220][6];				r_cell_reg[186] = inform_R[157][6];				r_cell_reg[187] = inform_R[221][6];				r_cell_reg[188] = inform_R[158][6];				r_cell_reg[189] = inform_R[222][6];				r_cell_reg[190] = inform_R[159][6];				r_cell_reg[191] = inform_R[223][6];				r_cell_reg[192] = inform_R[160][6];				r_cell_reg[193] = inform_R[224][6];				r_cell_reg[194] = inform_R[161][6];				r_cell_reg[195] = inform_R[225][6];				r_cell_reg[196] = inform_R[162][6];				r_cell_reg[197] = inform_R[226][6];				r_cell_reg[198] = inform_R[163][6];				r_cell_reg[199] = inform_R[227][6];				r_cell_reg[200] = inform_R[164][6];				r_cell_reg[201] = inform_R[228][6];				r_cell_reg[202] = inform_R[165][6];				r_cell_reg[203] = inform_R[229][6];				r_cell_reg[204] = inform_R[166][6];				r_cell_reg[205] = inform_R[230][6];				r_cell_reg[206] = inform_R[167][6];				r_cell_reg[207] = inform_R[231][6];				r_cell_reg[208] = inform_R[168][6];				r_cell_reg[209] = inform_R[232][6];				r_cell_reg[210] = inform_R[169][6];				r_cell_reg[211] = inform_R[233][6];				r_cell_reg[212] = inform_R[170][6];				r_cell_reg[213] = inform_R[234][6];				r_cell_reg[214] = inform_R[171][6];				r_cell_reg[215] = inform_R[235][6];				r_cell_reg[216] = inform_R[172][6];				r_cell_reg[217] = inform_R[236][6];				r_cell_reg[218] = inform_R[173][6];				r_cell_reg[219] = inform_R[237][6];				r_cell_reg[220] = inform_R[174][6];				r_cell_reg[221] = inform_R[238][6];				r_cell_reg[222] = inform_R[175][6];				r_cell_reg[223] = inform_R[239][6];				r_cell_reg[224] = inform_R[176][6];				r_cell_reg[225] = inform_R[240][6];				r_cell_reg[226] = inform_R[177][6];				r_cell_reg[227] = inform_R[241][6];				r_cell_reg[228] = inform_R[178][6];				r_cell_reg[229] = inform_R[242][6];				r_cell_reg[230] = inform_R[179][6];				r_cell_reg[231] = inform_R[243][6];				r_cell_reg[232] = inform_R[180][6];				r_cell_reg[233] = inform_R[244][6];				r_cell_reg[234] = inform_R[181][6];				r_cell_reg[235] = inform_R[245][6];				r_cell_reg[236] = inform_R[182][6];				r_cell_reg[237] = inform_R[246][6];				r_cell_reg[238] = inform_R[183][6];				r_cell_reg[239] = inform_R[247][6];				r_cell_reg[240] = inform_R[184][6];				r_cell_reg[241] = inform_R[248][6];				r_cell_reg[242] = inform_R[185][6];				r_cell_reg[243] = inform_R[249][6];				r_cell_reg[244] = inform_R[186][6];				r_cell_reg[245] = inform_R[250][6];				r_cell_reg[246] = inform_R[187][6];				r_cell_reg[247] = inform_R[251][6];				r_cell_reg[248] = inform_R[188][6];				r_cell_reg[249] = inform_R[252][6];				r_cell_reg[250] = inform_R[189][6];				r_cell_reg[251] = inform_R[253][6];				r_cell_reg[252] = inform_R[190][6];				r_cell_reg[253] = inform_R[254][6];				r_cell_reg[254] = inform_R[191][6];				r_cell_reg[255] = inform_R[255][6];				l_cell_reg[0] = inform_L[0][7];				l_cell_reg[1] = inform_L[64][7];				l_cell_reg[2] = inform_L[1][7];				l_cell_reg[3] = inform_L[65][7];				l_cell_reg[4] = inform_L[2][7];				l_cell_reg[5] = inform_L[66][7];				l_cell_reg[6] = inform_L[3][7];				l_cell_reg[7] = inform_L[67][7];				l_cell_reg[8] = inform_L[4][7];				l_cell_reg[9] = inform_L[68][7];				l_cell_reg[10] = inform_L[5][7];				l_cell_reg[11] = inform_L[69][7];				l_cell_reg[12] = inform_L[6][7];				l_cell_reg[13] = inform_L[70][7];				l_cell_reg[14] = inform_L[7][7];				l_cell_reg[15] = inform_L[71][7];				l_cell_reg[16] = inform_L[8][7];				l_cell_reg[17] = inform_L[72][7];				l_cell_reg[18] = inform_L[9][7];				l_cell_reg[19] = inform_L[73][7];				l_cell_reg[20] = inform_L[10][7];				l_cell_reg[21] = inform_L[74][7];				l_cell_reg[22] = inform_L[11][7];				l_cell_reg[23] = inform_L[75][7];				l_cell_reg[24] = inform_L[12][7];				l_cell_reg[25] = inform_L[76][7];				l_cell_reg[26] = inform_L[13][7];				l_cell_reg[27] = inform_L[77][7];				l_cell_reg[28] = inform_L[14][7];				l_cell_reg[29] = inform_L[78][7];				l_cell_reg[30] = inform_L[15][7];				l_cell_reg[31] = inform_L[79][7];				l_cell_reg[32] = inform_L[16][7];				l_cell_reg[33] = inform_L[80][7];				l_cell_reg[34] = inform_L[17][7];				l_cell_reg[35] = inform_L[81][7];				l_cell_reg[36] = inform_L[18][7];				l_cell_reg[37] = inform_L[82][7];				l_cell_reg[38] = inform_L[19][7];				l_cell_reg[39] = inform_L[83][7];				l_cell_reg[40] = inform_L[20][7];				l_cell_reg[41] = inform_L[84][7];				l_cell_reg[42] = inform_L[21][7];				l_cell_reg[43] = inform_L[85][7];				l_cell_reg[44] = inform_L[22][7];				l_cell_reg[45] = inform_L[86][7];				l_cell_reg[46] = inform_L[23][7];				l_cell_reg[47] = inform_L[87][7];				l_cell_reg[48] = inform_L[24][7];				l_cell_reg[49] = inform_L[88][7];				l_cell_reg[50] = inform_L[25][7];				l_cell_reg[51] = inform_L[89][7];				l_cell_reg[52] = inform_L[26][7];				l_cell_reg[53] = inform_L[90][7];				l_cell_reg[54] = inform_L[27][7];				l_cell_reg[55] = inform_L[91][7];				l_cell_reg[56] = inform_L[28][7];				l_cell_reg[57] = inform_L[92][7];				l_cell_reg[58] = inform_L[29][7];				l_cell_reg[59] = inform_L[93][7];				l_cell_reg[60] = inform_L[30][7];				l_cell_reg[61] = inform_L[94][7];				l_cell_reg[62] = inform_L[31][7];				l_cell_reg[63] = inform_L[95][7];				l_cell_reg[64] = inform_L[32][7];				l_cell_reg[65] = inform_L[96][7];				l_cell_reg[66] = inform_L[33][7];				l_cell_reg[67] = inform_L[97][7];				l_cell_reg[68] = inform_L[34][7];				l_cell_reg[69] = inform_L[98][7];				l_cell_reg[70] = inform_L[35][7];				l_cell_reg[71] = inform_L[99][7];				l_cell_reg[72] = inform_L[36][7];				l_cell_reg[73] = inform_L[100][7];				l_cell_reg[74] = inform_L[37][7];				l_cell_reg[75] = inform_L[101][7];				l_cell_reg[76] = inform_L[38][7];				l_cell_reg[77] = inform_L[102][7];				l_cell_reg[78] = inform_L[39][7];				l_cell_reg[79] = inform_L[103][7];				l_cell_reg[80] = inform_L[40][7];				l_cell_reg[81] = inform_L[104][7];				l_cell_reg[82] = inform_L[41][7];				l_cell_reg[83] = inform_L[105][7];				l_cell_reg[84] = inform_L[42][7];				l_cell_reg[85] = inform_L[106][7];				l_cell_reg[86] = inform_L[43][7];				l_cell_reg[87] = inform_L[107][7];				l_cell_reg[88] = inform_L[44][7];				l_cell_reg[89] = inform_L[108][7];				l_cell_reg[90] = inform_L[45][7];				l_cell_reg[91] = inform_L[109][7];				l_cell_reg[92] = inform_L[46][7];				l_cell_reg[93] = inform_L[110][7];				l_cell_reg[94] = inform_L[47][7];				l_cell_reg[95] = inform_L[111][7];				l_cell_reg[96] = inform_L[48][7];				l_cell_reg[97] = inform_L[112][7];				l_cell_reg[98] = inform_L[49][7];				l_cell_reg[99] = inform_L[113][7];				l_cell_reg[100] = inform_L[50][7];				l_cell_reg[101] = inform_L[114][7];				l_cell_reg[102] = inform_L[51][7];				l_cell_reg[103] = inform_L[115][7];				l_cell_reg[104] = inform_L[52][7];				l_cell_reg[105] = inform_L[116][7];				l_cell_reg[106] = inform_L[53][7];				l_cell_reg[107] = inform_L[117][7];				l_cell_reg[108] = inform_L[54][7];				l_cell_reg[109] = inform_L[118][7];				l_cell_reg[110] = inform_L[55][7];				l_cell_reg[111] = inform_L[119][7];				l_cell_reg[112] = inform_L[56][7];				l_cell_reg[113] = inform_L[120][7];				l_cell_reg[114] = inform_L[57][7];				l_cell_reg[115] = inform_L[121][7];				l_cell_reg[116] = inform_L[58][7];				l_cell_reg[117] = inform_L[122][7];				l_cell_reg[118] = inform_L[59][7];				l_cell_reg[119] = inform_L[123][7];				l_cell_reg[120] = inform_L[60][7];				l_cell_reg[121] = inform_L[124][7];				l_cell_reg[122] = inform_L[61][7];				l_cell_reg[123] = inform_L[125][7];				l_cell_reg[124] = inform_L[62][7];				l_cell_reg[125] = inform_L[126][7];				l_cell_reg[126] = inform_L[63][7];				l_cell_reg[127] = inform_L[127][7];				l_cell_reg[128] = inform_L[128][7];				l_cell_reg[129] = inform_L[192][7];				l_cell_reg[130] = inform_L[129][7];				l_cell_reg[131] = inform_L[193][7];				l_cell_reg[132] = inform_L[130][7];				l_cell_reg[133] = inform_L[194][7];				l_cell_reg[134] = inform_L[131][7];				l_cell_reg[135] = inform_L[195][7];				l_cell_reg[136] = inform_L[132][7];				l_cell_reg[137] = inform_L[196][7];				l_cell_reg[138] = inform_L[133][7];				l_cell_reg[139] = inform_L[197][7];				l_cell_reg[140] = inform_L[134][7];				l_cell_reg[141] = inform_L[198][7];				l_cell_reg[142] = inform_L[135][7];				l_cell_reg[143] = inform_L[199][7];				l_cell_reg[144] = inform_L[136][7];				l_cell_reg[145] = inform_L[200][7];				l_cell_reg[146] = inform_L[137][7];				l_cell_reg[147] = inform_L[201][7];				l_cell_reg[148] = inform_L[138][7];				l_cell_reg[149] = inform_L[202][7];				l_cell_reg[150] = inform_L[139][7];				l_cell_reg[151] = inform_L[203][7];				l_cell_reg[152] = inform_L[140][7];				l_cell_reg[153] = inform_L[204][7];				l_cell_reg[154] = inform_L[141][7];				l_cell_reg[155] = inform_L[205][7];				l_cell_reg[156] = inform_L[142][7];				l_cell_reg[157] = inform_L[206][7];				l_cell_reg[158] = inform_L[143][7];				l_cell_reg[159] = inform_L[207][7];				l_cell_reg[160] = inform_L[144][7];				l_cell_reg[161] = inform_L[208][7];				l_cell_reg[162] = inform_L[145][7];				l_cell_reg[163] = inform_L[209][7];				l_cell_reg[164] = inform_L[146][7];				l_cell_reg[165] = inform_L[210][7];				l_cell_reg[166] = inform_L[147][7];				l_cell_reg[167] = inform_L[211][7];				l_cell_reg[168] = inform_L[148][7];				l_cell_reg[169] = inform_L[212][7];				l_cell_reg[170] = inform_L[149][7];				l_cell_reg[171] = inform_L[213][7];				l_cell_reg[172] = inform_L[150][7];				l_cell_reg[173] = inform_L[214][7];				l_cell_reg[174] = inform_L[151][7];				l_cell_reg[175] = inform_L[215][7];				l_cell_reg[176] = inform_L[152][7];				l_cell_reg[177] = inform_L[216][7];				l_cell_reg[178] = inform_L[153][7];				l_cell_reg[179] = inform_L[217][7];				l_cell_reg[180] = inform_L[154][7];				l_cell_reg[181] = inform_L[218][7];				l_cell_reg[182] = inform_L[155][7];				l_cell_reg[183] = inform_L[219][7];				l_cell_reg[184] = inform_L[156][7];				l_cell_reg[185] = inform_L[220][7];				l_cell_reg[186] = inform_L[157][7];				l_cell_reg[187] = inform_L[221][7];				l_cell_reg[188] = inform_L[158][7];				l_cell_reg[189] = inform_L[222][7];				l_cell_reg[190] = inform_L[159][7];				l_cell_reg[191] = inform_L[223][7];				l_cell_reg[192] = inform_L[160][7];				l_cell_reg[193] = inform_L[224][7];				l_cell_reg[194] = inform_L[161][7];				l_cell_reg[195] = inform_L[225][7];				l_cell_reg[196] = inform_L[162][7];				l_cell_reg[197] = inform_L[226][7];				l_cell_reg[198] = inform_L[163][7];				l_cell_reg[199] = inform_L[227][7];				l_cell_reg[200] = inform_L[164][7];				l_cell_reg[201] = inform_L[228][7];				l_cell_reg[202] = inform_L[165][7];				l_cell_reg[203] = inform_L[229][7];				l_cell_reg[204] = inform_L[166][7];				l_cell_reg[205] = inform_L[230][7];				l_cell_reg[206] = inform_L[167][7];				l_cell_reg[207] = inform_L[231][7];				l_cell_reg[208] = inform_L[168][7];				l_cell_reg[209] = inform_L[232][7];				l_cell_reg[210] = inform_L[169][7];				l_cell_reg[211] = inform_L[233][7];				l_cell_reg[212] = inform_L[170][7];				l_cell_reg[213] = inform_L[234][7];				l_cell_reg[214] = inform_L[171][7];				l_cell_reg[215] = inform_L[235][7];				l_cell_reg[216] = inform_L[172][7];				l_cell_reg[217] = inform_L[236][7];				l_cell_reg[218] = inform_L[173][7];				l_cell_reg[219] = inform_L[237][7];				l_cell_reg[220] = inform_L[174][7];				l_cell_reg[221] = inform_L[238][7];				l_cell_reg[222] = inform_L[175][7];				l_cell_reg[223] = inform_L[239][7];				l_cell_reg[224] = inform_L[176][7];				l_cell_reg[225] = inform_L[240][7];				l_cell_reg[226] = inform_L[177][7];				l_cell_reg[227] = inform_L[241][7];				l_cell_reg[228] = inform_L[178][7];				l_cell_reg[229] = inform_L[242][7];				l_cell_reg[230] = inform_L[179][7];				l_cell_reg[231] = inform_L[243][7];				l_cell_reg[232] = inform_L[180][7];				l_cell_reg[233] = inform_L[244][7];				l_cell_reg[234] = inform_L[181][7];				l_cell_reg[235] = inform_L[245][7];				l_cell_reg[236] = inform_L[182][7];				l_cell_reg[237] = inform_L[246][7];				l_cell_reg[238] = inform_L[183][7];				l_cell_reg[239] = inform_L[247][7];				l_cell_reg[240] = inform_L[184][7];				l_cell_reg[241] = inform_L[248][7];				l_cell_reg[242] = inform_L[185][7];				l_cell_reg[243] = inform_L[249][7];				l_cell_reg[244] = inform_L[186][7];				l_cell_reg[245] = inform_L[250][7];				l_cell_reg[246] = inform_L[187][7];				l_cell_reg[247] = inform_L[251][7];				l_cell_reg[248] = inform_L[188][7];				l_cell_reg[249] = inform_L[252][7];				l_cell_reg[250] = inform_L[189][7];				l_cell_reg[251] = inform_L[253][7];				l_cell_reg[252] = inform_L[190][7];				l_cell_reg[253] = inform_L[254][7];				l_cell_reg[254] = inform_L[191][7];				l_cell_reg[255] = inform_L[255][7];			end
			8:			begin				r_cell_reg[0] = inform_R[0][7];				r_cell_reg[1] = inform_R[128][7];				r_cell_reg[2] = inform_R[1][7];				r_cell_reg[3] = inform_R[129][7];				r_cell_reg[4] = inform_R[2][7];				r_cell_reg[5] = inform_R[130][7];				r_cell_reg[6] = inform_R[3][7];				r_cell_reg[7] = inform_R[131][7];				r_cell_reg[8] = inform_R[4][7];				r_cell_reg[9] = inform_R[132][7];				r_cell_reg[10] = inform_R[5][7];				r_cell_reg[11] = inform_R[133][7];				r_cell_reg[12] = inform_R[6][7];				r_cell_reg[13] = inform_R[134][7];				r_cell_reg[14] = inform_R[7][7];				r_cell_reg[15] = inform_R[135][7];				r_cell_reg[16] = inform_R[8][7];				r_cell_reg[17] = inform_R[136][7];				r_cell_reg[18] = inform_R[9][7];				r_cell_reg[19] = inform_R[137][7];				r_cell_reg[20] = inform_R[10][7];				r_cell_reg[21] = inform_R[138][7];				r_cell_reg[22] = inform_R[11][7];				r_cell_reg[23] = inform_R[139][7];				r_cell_reg[24] = inform_R[12][7];				r_cell_reg[25] = inform_R[140][7];				r_cell_reg[26] = inform_R[13][7];				r_cell_reg[27] = inform_R[141][7];				r_cell_reg[28] = inform_R[14][7];				r_cell_reg[29] = inform_R[142][7];				r_cell_reg[30] = inform_R[15][7];				r_cell_reg[31] = inform_R[143][7];				r_cell_reg[32] = inform_R[16][7];				r_cell_reg[33] = inform_R[144][7];				r_cell_reg[34] = inform_R[17][7];				r_cell_reg[35] = inform_R[145][7];				r_cell_reg[36] = inform_R[18][7];				r_cell_reg[37] = inform_R[146][7];				r_cell_reg[38] = inform_R[19][7];				r_cell_reg[39] = inform_R[147][7];				r_cell_reg[40] = inform_R[20][7];				r_cell_reg[41] = inform_R[148][7];				r_cell_reg[42] = inform_R[21][7];				r_cell_reg[43] = inform_R[149][7];				r_cell_reg[44] = inform_R[22][7];				r_cell_reg[45] = inform_R[150][7];				r_cell_reg[46] = inform_R[23][7];				r_cell_reg[47] = inform_R[151][7];				r_cell_reg[48] = inform_R[24][7];				r_cell_reg[49] = inform_R[152][7];				r_cell_reg[50] = inform_R[25][7];				r_cell_reg[51] = inform_R[153][7];				r_cell_reg[52] = inform_R[26][7];				r_cell_reg[53] = inform_R[154][7];				r_cell_reg[54] = inform_R[27][7];				r_cell_reg[55] = inform_R[155][7];				r_cell_reg[56] = inform_R[28][7];				r_cell_reg[57] = inform_R[156][7];				r_cell_reg[58] = inform_R[29][7];				r_cell_reg[59] = inform_R[157][7];				r_cell_reg[60] = inform_R[30][7];				r_cell_reg[61] = inform_R[158][7];				r_cell_reg[62] = inform_R[31][7];				r_cell_reg[63] = inform_R[159][7];				r_cell_reg[64] = inform_R[32][7];				r_cell_reg[65] = inform_R[160][7];				r_cell_reg[66] = inform_R[33][7];				r_cell_reg[67] = inform_R[161][7];				r_cell_reg[68] = inform_R[34][7];				r_cell_reg[69] = inform_R[162][7];				r_cell_reg[70] = inform_R[35][7];				r_cell_reg[71] = inform_R[163][7];				r_cell_reg[72] = inform_R[36][7];				r_cell_reg[73] = inform_R[164][7];				r_cell_reg[74] = inform_R[37][7];				r_cell_reg[75] = inform_R[165][7];				r_cell_reg[76] = inform_R[38][7];				r_cell_reg[77] = inform_R[166][7];				r_cell_reg[78] = inform_R[39][7];				r_cell_reg[79] = inform_R[167][7];				r_cell_reg[80] = inform_R[40][7];				r_cell_reg[81] = inform_R[168][7];				r_cell_reg[82] = inform_R[41][7];				r_cell_reg[83] = inform_R[169][7];				r_cell_reg[84] = inform_R[42][7];				r_cell_reg[85] = inform_R[170][7];				r_cell_reg[86] = inform_R[43][7];				r_cell_reg[87] = inform_R[171][7];				r_cell_reg[88] = inform_R[44][7];				r_cell_reg[89] = inform_R[172][7];				r_cell_reg[90] = inform_R[45][7];				r_cell_reg[91] = inform_R[173][7];				r_cell_reg[92] = inform_R[46][7];				r_cell_reg[93] = inform_R[174][7];				r_cell_reg[94] = inform_R[47][7];				r_cell_reg[95] = inform_R[175][7];				r_cell_reg[96] = inform_R[48][7];				r_cell_reg[97] = inform_R[176][7];				r_cell_reg[98] = inform_R[49][7];				r_cell_reg[99] = inform_R[177][7];				r_cell_reg[100] = inform_R[50][7];				r_cell_reg[101] = inform_R[178][7];				r_cell_reg[102] = inform_R[51][7];				r_cell_reg[103] = inform_R[179][7];				r_cell_reg[104] = inform_R[52][7];				r_cell_reg[105] = inform_R[180][7];				r_cell_reg[106] = inform_R[53][7];				r_cell_reg[107] = inform_R[181][7];				r_cell_reg[108] = inform_R[54][7];				r_cell_reg[109] = inform_R[182][7];				r_cell_reg[110] = inform_R[55][7];				r_cell_reg[111] = inform_R[183][7];				r_cell_reg[112] = inform_R[56][7];				r_cell_reg[113] = inform_R[184][7];				r_cell_reg[114] = inform_R[57][7];				r_cell_reg[115] = inform_R[185][7];				r_cell_reg[116] = inform_R[58][7];				r_cell_reg[117] = inform_R[186][7];				r_cell_reg[118] = inform_R[59][7];				r_cell_reg[119] = inform_R[187][7];				r_cell_reg[120] = inform_R[60][7];				r_cell_reg[121] = inform_R[188][7];				r_cell_reg[122] = inform_R[61][7];				r_cell_reg[123] = inform_R[189][7];				r_cell_reg[124] = inform_R[62][7];				r_cell_reg[125] = inform_R[190][7];				r_cell_reg[126] = inform_R[63][7];				r_cell_reg[127] = inform_R[191][7];				r_cell_reg[128] = inform_R[64][7];				r_cell_reg[129] = inform_R[192][7];				r_cell_reg[130] = inform_R[65][7];				r_cell_reg[131] = inform_R[193][7];				r_cell_reg[132] = inform_R[66][7];				r_cell_reg[133] = inform_R[194][7];				r_cell_reg[134] = inform_R[67][7];				r_cell_reg[135] = inform_R[195][7];				r_cell_reg[136] = inform_R[68][7];				r_cell_reg[137] = inform_R[196][7];				r_cell_reg[138] = inform_R[69][7];				r_cell_reg[139] = inform_R[197][7];				r_cell_reg[140] = inform_R[70][7];				r_cell_reg[141] = inform_R[198][7];				r_cell_reg[142] = inform_R[71][7];				r_cell_reg[143] = inform_R[199][7];				r_cell_reg[144] = inform_R[72][7];				r_cell_reg[145] = inform_R[200][7];				r_cell_reg[146] = inform_R[73][7];				r_cell_reg[147] = inform_R[201][7];				r_cell_reg[148] = inform_R[74][7];				r_cell_reg[149] = inform_R[202][7];				r_cell_reg[150] = inform_R[75][7];				r_cell_reg[151] = inform_R[203][7];				r_cell_reg[152] = inform_R[76][7];				r_cell_reg[153] = inform_R[204][7];				r_cell_reg[154] = inform_R[77][7];				r_cell_reg[155] = inform_R[205][7];				r_cell_reg[156] = inform_R[78][7];				r_cell_reg[157] = inform_R[206][7];				r_cell_reg[158] = inform_R[79][7];				r_cell_reg[159] = inform_R[207][7];				r_cell_reg[160] = inform_R[80][7];				r_cell_reg[161] = inform_R[208][7];				r_cell_reg[162] = inform_R[81][7];				r_cell_reg[163] = inform_R[209][7];				r_cell_reg[164] = inform_R[82][7];				r_cell_reg[165] = inform_R[210][7];				r_cell_reg[166] = inform_R[83][7];				r_cell_reg[167] = inform_R[211][7];				r_cell_reg[168] = inform_R[84][7];				r_cell_reg[169] = inform_R[212][7];				r_cell_reg[170] = inform_R[85][7];				r_cell_reg[171] = inform_R[213][7];				r_cell_reg[172] = inform_R[86][7];				r_cell_reg[173] = inform_R[214][7];				r_cell_reg[174] = inform_R[87][7];				r_cell_reg[175] = inform_R[215][7];				r_cell_reg[176] = inform_R[88][7];				r_cell_reg[177] = inform_R[216][7];				r_cell_reg[178] = inform_R[89][7];				r_cell_reg[179] = inform_R[217][7];				r_cell_reg[180] = inform_R[90][7];				r_cell_reg[181] = inform_R[218][7];				r_cell_reg[182] = inform_R[91][7];				r_cell_reg[183] = inform_R[219][7];				r_cell_reg[184] = inform_R[92][7];				r_cell_reg[185] = inform_R[220][7];				r_cell_reg[186] = inform_R[93][7];				r_cell_reg[187] = inform_R[221][7];				r_cell_reg[188] = inform_R[94][7];				r_cell_reg[189] = inform_R[222][7];				r_cell_reg[190] = inform_R[95][7];				r_cell_reg[191] = inform_R[223][7];				r_cell_reg[192] = inform_R[96][7];				r_cell_reg[193] = inform_R[224][7];				r_cell_reg[194] = inform_R[97][7];				r_cell_reg[195] = inform_R[225][7];				r_cell_reg[196] = inform_R[98][7];				r_cell_reg[197] = inform_R[226][7];				r_cell_reg[198] = inform_R[99][7];				r_cell_reg[199] = inform_R[227][7];				r_cell_reg[200] = inform_R[100][7];				r_cell_reg[201] = inform_R[228][7];				r_cell_reg[202] = inform_R[101][7];				r_cell_reg[203] = inform_R[229][7];				r_cell_reg[204] = inform_R[102][7];				r_cell_reg[205] = inform_R[230][7];				r_cell_reg[206] = inform_R[103][7];				r_cell_reg[207] = inform_R[231][7];				r_cell_reg[208] = inform_R[104][7];				r_cell_reg[209] = inform_R[232][7];				r_cell_reg[210] = inform_R[105][7];				r_cell_reg[211] = inform_R[233][7];				r_cell_reg[212] = inform_R[106][7];				r_cell_reg[213] = inform_R[234][7];				r_cell_reg[214] = inform_R[107][7];				r_cell_reg[215] = inform_R[235][7];				r_cell_reg[216] = inform_R[108][7];				r_cell_reg[217] = inform_R[236][7];				r_cell_reg[218] = inform_R[109][7];				r_cell_reg[219] = inform_R[237][7];				r_cell_reg[220] = inform_R[110][7];				r_cell_reg[221] = inform_R[238][7];				r_cell_reg[222] = inform_R[111][7];				r_cell_reg[223] = inform_R[239][7];				r_cell_reg[224] = inform_R[112][7];				r_cell_reg[225] = inform_R[240][7];				r_cell_reg[226] = inform_R[113][7];				r_cell_reg[227] = inform_R[241][7];				r_cell_reg[228] = inform_R[114][7];				r_cell_reg[229] = inform_R[242][7];				r_cell_reg[230] = inform_R[115][7];				r_cell_reg[231] = inform_R[243][7];				r_cell_reg[232] = inform_R[116][7];				r_cell_reg[233] = inform_R[244][7];				r_cell_reg[234] = inform_R[117][7];				r_cell_reg[235] = inform_R[245][7];				r_cell_reg[236] = inform_R[118][7];				r_cell_reg[237] = inform_R[246][7];				r_cell_reg[238] = inform_R[119][7];				r_cell_reg[239] = inform_R[247][7];				r_cell_reg[240] = inform_R[120][7];				r_cell_reg[241] = inform_R[248][7];				r_cell_reg[242] = inform_R[121][7];				r_cell_reg[243] = inform_R[249][7];				r_cell_reg[244] = inform_R[122][7];				r_cell_reg[245] = inform_R[250][7];				r_cell_reg[246] = inform_R[123][7];				r_cell_reg[247] = inform_R[251][7];				r_cell_reg[248] = inform_R[124][7];				r_cell_reg[249] = inform_R[252][7];				r_cell_reg[250] = inform_R[125][7];				r_cell_reg[251] = inform_R[253][7];				r_cell_reg[252] = inform_R[126][7];				r_cell_reg[253] = inform_R[254][7];				r_cell_reg[254] = inform_R[127][7];				r_cell_reg[255] = inform_R[255][7];				l_cell_reg[0] = inform_L[0][8];				l_cell_reg[1] = inform_L[128][8];				l_cell_reg[2] = inform_L[1][8];				l_cell_reg[3] = inform_L[129][8];				l_cell_reg[4] = inform_L[2][8];				l_cell_reg[5] = inform_L[130][8];				l_cell_reg[6] = inform_L[3][8];				l_cell_reg[7] = inform_L[131][8];				l_cell_reg[8] = inform_L[4][8];				l_cell_reg[9] = inform_L[132][8];				l_cell_reg[10] = inform_L[5][8];				l_cell_reg[11] = inform_L[133][8];				l_cell_reg[12] = inform_L[6][8];				l_cell_reg[13] = inform_L[134][8];				l_cell_reg[14] = inform_L[7][8];				l_cell_reg[15] = inform_L[135][8];				l_cell_reg[16] = inform_L[8][8];				l_cell_reg[17] = inform_L[136][8];				l_cell_reg[18] = inform_L[9][8];				l_cell_reg[19] = inform_L[137][8];				l_cell_reg[20] = inform_L[10][8];				l_cell_reg[21] = inform_L[138][8];				l_cell_reg[22] = inform_L[11][8];				l_cell_reg[23] = inform_L[139][8];				l_cell_reg[24] = inform_L[12][8];				l_cell_reg[25] = inform_L[140][8];				l_cell_reg[26] = inform_L[13][8];				l_cell_reg[27] = inform_L[141][8];				l_cell_reg[28] = inform_L[14][8];				l_cell_reg[29] = inform_L[142][8];				l_cell_reg[30] = inform_L[15][8];				l_cell_reg[31] = inform_L[143][8];				l_cell_reg[32] = inform_L[16][8];				l_cell_reg[33] = inform_L[144][8];				l_cell_reg[34] = inform_L[17][8];				l_cell_reg[35] = inform_L[145][8];				l_cell_reg[36] = inform_L[18][8];				l_cell_reg[37] = inform_L[146][8];				l_cell_reg[38] = inform_L[19][8];				l_cell_reg[39] = inform_L[147][8];				l_cell_reg[40] = inform_L[20][8];				l_cell_reg[41] = inform_L[148][8];				l_cell_reg[42] = inform_L[21][8];				l_cell_reg[43] = inform_L[149][8];				l_cell_reg[44] = inform_L[22][8];				l_cell_reg[45] = inform_L[150][8];				l_cell_reg[46] = inform_L[23][8];				l_cell_reg[47] = inform_L[151][8];				l_cell_reg[48] = inform_L[24][8];				l_cell_reg[49] = inform_L[152][8];				l_cell_reg[50] = inform_L[25][8];				l_cell_reg[51] = inform_L[153][8];				l_cell_reg[52] = inform_L[26][8];				l_cell_reg[53] = inform_L[154][8];				l_cell_reg[54] = inform_L[27][8];				l_cell_reg[55] = inform_L[155][8];				l_cell_reg[56] = inform_L[28][8];				l_cell_reg[57] = inform_L[156][8];				l_cell_reg[58] = inform_L[29][8];				l_cell_reg[59] = inform_L[157][8];				l_cell_reg[60] = inform_L[30][8];				l_cell_reg[61] = inform_L[158][8];				l_cell_reg[62] = inform_L[31][8];				l_cell_reg[63] = inform_L[159][8];				l_cell_reg[64] = inform_L[32][8];				l_cell_reg[65] = inform_L[160][8];				l_cell_reg[66] = inform_L[33][8];				l_cell_reg[67] = inform_L[161][8];				l_cell_reg[68] = inform_L[34][8];				l_cell_reg[69] = inform_L[162][8];				l_cell_reg[70] = inform_L[35][8];				l_cell_reg[71] = inform_L[163][8];				l_cell_reg[72] = inform_L[36][8];				l_cell_reg[73] = inform_L[164][8];				l_cell_reg[74] = inform_L[37][8];				l_cell_reg[75] = inform_L[165][8];				l_cell_reg[76] = inform_L[38][8];				l_cell_reg[77] = inform_L[166][8];				l_cell_reg[78] = inform_L[39][8];				l_cell_reg[79] = inform_L[167][8];				l_cell_reg[80] = inform_L[40][8];				l_cell_reg[81] = inform_L[168][8];				l_cell_reg[82] = inform_L[41][8];				l_cell_reg[83] = inform_L[169][8];				l_cell_reg[84] = inform_L[42][8];				l_cell_reg[85] = inform_L[170][8];				l_cell_reg[86] = inform_L[43][8];				l_cell_reg[87] = inform_L[171][8];				l_cell_reg[88] = inform_L[44][8];				l_cell_reg[89] = inform_L[172][8];				l_cell_reg[90] = inform_L[45][8];				l_cell_reg[91] = inform_L[173][8];				l_cell_reg[92] = inform_L[46][8];				l_cell_reg[93] = inform_L[174][8];				l_cell_reg[94] = inform_L[47][8];				l_cell_reg[95] = inform_L[175][8];				l_cell_reg[96] = inform_L[48][8];				l_cell_reg[97] = inform_L[176][8];				l_cell_reg[98] = inform_L[49][8];				l_cell_reg[99] = inform_L[177][8];				l_cell_reg[100] = inform_L[50][8];				l_cell_reg[101] = inform_L[178][8];				l_cell_reg[102] = inform_L[51][8];				l_cell_reg[103] = inform_L[179][8];				l_cell_reg[104] = inform_L[52][8];				l_cell_reg[105] = inform_L[180][8];				l_cell_reg[106] = inform_L[53][8];				l_cell_reg[107] = inform_L[181][8];				l_cell_reg[108] = inform_L[54][8];				l_cell_reg[109] = inform_L[182][8];				l_cell_reg[110] = inform_L[55][8];				l_cell_reg[111] = inform_L[183][8];				l_cell_reg[112] = inform_L[56][8];				l_cell_reg[113] = inform_L[184][8];				l_cell_reg[114] = inform_L[57][8];				l_cell_reg[115] = inform_L[185][8];				l_cell_reg[116] = inform_L[58][8];				l_cell_reg[117] = inform_L[186][8];				l_cell_reg[118] = inform_L[59][8];				l_cell_reg[119] = inform_L[187][8];				l_cell_reg[120] = inform_L[60][8];				l_cell_reg[121] = inform_L[188][8];				l_cell_reg[122] = inform_L[61][8];				l_cell_reg[123] = inform_L[189][8];				l_cell_reg[124] = inform_L[62][8];				l_cell_reg[125] = inform_L[190][8];				l_cell_reg[126] = inform_L[63][8];				l_cell_reg[127] = inform_L[191][8];				l_cell_reg[128] = inform_L[64][8];				l_cell_reg[129] = inform_L[192][8];				l_cell_reg[130] = inform_L[65][8];				l_cell_reg[131] = inform_L[193][8];				l_cell_reg[132] = inform_L[66][8];				l_cell_reg[133] = inform_L[194][8];				l_cell_reg[134] = inform_L[67][8];				l_cell_reg[135] = inform_L[195][8];				l_cell_reg[136] = inform_L[68][8];				l_cell_reg[137] = inform_L[196][8];				l_cell_reg[138] = inform_L[69][8];				l_cell_reg[139] = inform_L[197][8];				l_cell_reg[140] = inform_L[70][8];				l_cell_reg[141] = inform_L[198][8];				l_cell_reg[142] = inform_L[71][8];				l_cell_reg[143] = inform_L[199][8];				l_cell_reg[144] = inform_L[72][8];				l_cell_reg[145] = inform_L[200][8];				l_cell_reg[146] = inform_L[73][8];				l_cell_reg[147] = inform_L[201][8];				l_cell_reg[148] = inform_L[74][8];				l_cell_reg[149] = inform_L[202][8];				l_cell_reg[150] = inform_L[75][8];				l_cell_reg[151] = inform_L[203][8];				l_cell_reg[152] = inform_L[76][8];				l_cell_reg[153] = inform_L[204][8];				l_cell_reg[154] = inform_L[77][8];				l_cell_reg[155] = inform_L[205][8];				l_cell_reg[156] = inform_L[78][8];				l_cell_reg[157] = inform_L[206][8];				l_cell_reg[158] = inform_L[79][8];				l_cell_reg[159] = inform_L[207][8];				l_cell_reg[160] = inform_L[80][8];				l_cell_reg[161] = inform_L[208][8];				l_cell_reg[162] = inform_L[81][8];				l_cell_reg[163] = inform_L[209][8];				l_cell_reg[164] = inform_L[82][8];				l_cell_reg[165] = inform_L[210][8];				l_cell_reg[166] = inform_L[83][8];				l_cell_reg[167] = inform_L[211][8];				l_cell_reg[168] = inform_L[84][8];				l_cell_reg[169] = inform_L[212][8];				l_cell_reg[170] = inform_L[85][8];				l_cell_reg[171] = inform_L[213][8];				l_cell_reg[172] = inform_L[86][8];				l_cell_reg[173] = inform_L[214][8];				l_cell_reg[174] = inform_L[87][8];				l_cell_reg[175] = inform_L[215][8];				l_cell_reg[176] = inform_L[88][8];				l_cell_reg[177] = inform_L[216][8];				l_cell_reg[178] = inform_L[89][8];				l_cell_reg[179] = inform_L[217][8];				l_cell_reg[180] = inform_L[90][8];				l_cell_reg[181] = inform_L[218][8];				l_cell_reg[182] = inform_L[91][8];				l_cell_reg[183] = inform_L[219][8];				l_cell_reg[184] = inform_L[92][8];				l_cell_reg[185] = inform_L[220][8];				l_cell_reg[186] = inform_L[93][8];				l_cell_reg[187] = inform_L[221][8];				l_cell_reg[188] = inform_L[94][8];				l_cell_reg[189] = inform_L[222][8];				l_cell_reg[190] = inform_L[95][8];				l_cell_reg[191] = inform_L[223][8];				l_cell_reg[192] = inform_L[96][8];				l_cell_reg[193] = inform_L[224][8];				l_cell_reg[194] = inform_L[97][8];				l_cell_reg[195] = inform_L[225][8];				l_cell_reg[196] = inform_L[98][8];				l_cell_reg[197] = inform_L[226][8];				l_cell_reg[198] = inform_L[99][8];				l_cell_reg[199] = inform_L[227][8];				l_cell_reg[200] = inform_L[100][8];				l_cell_reg[201] = inform_L[228][8];				l_cell_reg[202] = inform_L[101][8];				l_cell_reg[203] = inform_L[229][8];				l_cell_reg[204] = inform_L[102][8];				l_cell_reg[205] = inform_L[230][8];				l_cell_reg[206] = inform_L[103][8];				l_cell_reg[207] = inform_L[231][8];				l_cell_reg[208] = inform_L[104][8];				l_cell_reg[209] = inform_L[232][8];				l_cell_reg[210] = inform_L[105][8];				l_cell_reg[211] = inform_L[233][8];				l_cell_reg[212] = inform_L[106][8];				l_cell_reg[213] = inform_L[234][8];				l_cell_reg[214] = inform_L[107][8];				l_cell_reg[215] = inform_L[235][8];				l_cell_reg[216] = inform_L[108][8];				l_cell_reg[217] = inform_L[236][8];				l_cell_reg[218] = inform_L[109][8];				l_cell_reg[219] = inform_L[237][8];				l_cell_reg[220] = inform_L[110][8];				l_cell_reg[221] = inform_L[238][8];				l_cell_reg[222] = inform_L[111][8];				l_cell_reg[223] = inform_L[239][8];				l_cell_reg[224] = inform_L[112][8];				l_cell_reg[225] = inform_L[240][8];				l_cell_reg[226] = inform_L[113][8];				l_cell_reg[227] = inform_L[241][8];				l_cell_reg[228] = inform_L[114][8];				l_cell_reg[229] = inform_L[242][8];				l_cell_reg[230] = inform_L[115][8];				l_cell_reg[231] = inform_L[243][8];				l_cell_reg[232] = inform_L[116][8];				l_cell_reg[233] = inform_L[244][8];				l_cell_reg[234] = inform_L[117][8];				l_cell_reg[235] = inform_L[245][8];				l_cell_reg[236] = inform_L[118][8];				l_cell_reg[237] = inform_L[246][8];				l_cell_reg[238] = inform_L[119][8];				l_cell_reg[239] = inform_L[247][8];				l_cell_reg[240] = inform_L[120][8];				l_cell_reg[241] = inform_L[248][8];				l_cell_reg[242] = inform_L[121][8];				l_cell_reg[243] = inform_L[249][8];				l_cell_reg[244] = inform_L[122][8];				l_cell_reg[245] = inform_L[250][8];				l_cell_reg[246] = inform_L[123][8];				l_cell_reg[247] = inform_L[251][8];				l_cell_reg[248] = inform_L[124][8];				l_cell_reg[249] = inform_L[252][8];				l_cell_reg[250] = inform_L[125][8];				l_cell_reg[251] = inform_L[253][8];				l_cell_reg[252] = inform_L[126][8];				l_cell_reg[253] = inform_L[254][8];				l_cell_reg[254] = inform_L[127][8];				l_cell_reg[255] = inform_L[255][8];			end
			default:			begin					r_cell_reg[0] <= 0;					r_cell_reg[1] <= 0;					r_cell_reg[2] <= 0;					r_cell_reg[3] <= 0;					r_cell_reg[4] <= 0;					r_cell_reg[5] <= 0;					r_cell_reg[6] <= 0;					r_cell_reg[7] <= 0;					r_cell_reg[8] <= 0;					r_cell_reg[9] <= 0;					r_cell_reg[10] <= 0;					r_cell_reg[11] <= 0;					r_cell_reg[12] <= 0;					r_cell_reg[13] <= 0;					r_cell_reg[14] <= 0;					r_cell_reg[15] <= 0;					r_cell_reg[16] <= 0;					r_cell_reg[17] <= 0;					r_cell_reg[18] <= 0;					r_cell_reg[19] <= 0;					r_cell_reg[20] <= 0;					r_cell_reg[21] <= 0;					r_cell_reg[22] <= 0;					r_cell_reg[23] <= 0;					r_cell_reg[24] <= 0;					r_cell_reg[25] <= 0;					r_cell_reg[26] <= 0;					r_cell_reg[27] <= 0;					r_cell_reg[28] <= 0;					r_cell_reg[29] <= 0;					r_cell_reg[30] <= 0;					r_cell_reg[31] <= 0;					r_cell_reg[32] <= 0;					r_cell_reg[33] <= 0;					r_cell_reg[34] <= 0;					r_cell_reg[35] <= 0;					r_cell_reg[36] <= 0;					r_cell_reg[37] <= 0;					r_cell_reg[38] <= 0;					r_cell_reg[39] <= 0;					r_cell_reg[40] <= 0;					r_cell_reg[41] <= 0;					r_cell_reg[42] <= 0;					r_cell_reg[43] <= 0;					r_cell_reg[44] <= 0;					r_cell_reg[45] <= 0;					r_cell_reg[46] <= 0;					r_cell_reg[47] <= 0;					r_cell_reg[48] <= 0;					r_cell_reg[49] <= 0;					r_cell_reg[50] <= 0;					r_cell_reg[51] <= 0;					r_cell_reg[52] <= 0;					r_cell_reg[53] <= 0;					r_cell_reg[54] <= 0;					r_cell_reg[55] <= 0;					r_cell_reg[56] <= 0;					r_cell_reg[57] <= 0;					r_cell_reg[58] <= 0;					r_cell_reg[59] <= 0;					r_cell_reg[60] <= 0;					r_cell_reg[61] <= 0;					r_cell_reg[62] <= 0;					r_cell_reg[63] <= 0;					r_cell_reg[64] <= 0;					r_cell_reg[65] <= 0;					r_cell_reg[66] <= 0;					r_cell_reg[67] <= 0;					r_cell_reg[68] <= 0;					r_cell_reg[69] <= 0;					r_cell_reg[70] <= 0;					r_cell_reg[71] <= 0;					r_cell_reg[72] <= 0;					r_cell_reg[73] <= 0;					r_cell_reg[74] <= 0;					r_cell_reg[75] <= 0;					r_cell_reg[76] <= 0;					r_cell_reg[77] <= 0;					r_cell_reg[78] <= 0;					r_cell_reg[79] <= 0;					r_cell_reg[80] <= 0;					r_cell_reg[81] <= 0;					r_cell_reg[82] <= 0;					r_cell_reg[83] <= 0;					r_cell_reg[84] <= 0;					r_cell_reg[85] <= 0;					r_cell_reg[86] <= 0;					r_cell_reg[87] <= 0;					r_cell_reg[88] <= 0;					r_cell_reg[89] <= 0;					r_cell_reg[90] <= 0;					r_cell_reg[91] <= 0;					r_cell_reg[92] <= 0;					r_cell_reg[93] <= 0;					r_cell_reg[94] <= 0;					r_cell_reg[95] <= 0;					r_cell_reg[96] <= 0;					r_cell_reg[97] <= 0;					r_cell_reg[98] <= 0;					r_cell_reg[99] <= 0;					r_cell_reg[100] <= 0;					r_cell_reg[101] <= 0;					r_cell_reg[102] <= 0;					r_cell_reg[103] <= 0;					r_cell_reg[104] <= 0;					r_cell_reg[105] <= 0;					r_cell_reg[106] <= 0;					r_cell_reg[107] <= 0;					r_cell_reg[108] <= 0;					r_cell_reg[109] <= 0;					r_cell_reg[110] <= 0;					r_cell_reg[111] <= 0;					r_cell_reg[112] <= 0;					r_cell_reg[113] <= 0;					r_cell_reg[114] <= 0;					r_cell_reg[115] <= 0;					r_cell_reg[116] <= 0;					r_cell_reg[117] <= 0;					r_cell_reg[118] <= 0;					r_cell_reg[119] <= 0;					r_cell_reg[120] <= 0;					r_cell_reg[121] <= 0;					r_cell_reg[122] <= 0;					r_cell_reg[123] <= 0;					r_cell_reg[124] <= 0;					r_cell_reg[125] <= 0;					r_cell_reg[126] <= 0;					r_cell_reg[127] <= 0;					r_cell_reg[128] <= 0;					r_cell_reg[129] <= 0;					r_cell_reg[130] <= 0;					r_cell_reg[131] <= 0;					r_cell_reg[132] <= 0;					r_cell_reg[133] <= 0;					r_cell_reg[134] <= 0;					r_cell_reg[135] <= 0;					r_cell_reg[136] <= 0;					r_cell_reg[137] <= 0;					r_cell_reg[138] <= 0;					r_cell_reg[139] <= 0;					r_cell_reg[140] <= 0;					r_cell_reg[141] <= 0;					r_cell_reg[142] <= 0;					r_cell_reg[143] <= 0;					r_cell_reg[144] <= 0;					r_cell_reg[145] <= 0;					r_cell_reg[146] <= 0;					r_cell_reg[147] <= 0;					r_cell_reg[148] <= 0;					r_cell_reg[149] <= 0;					r_cell_reg[150] <= 0;					r_cell_reg[151] <= 0;					r_cell_reg[152] <= 0;					r_cell_reg[153] <= 0;					r_cell_reg[154] <= 0;					r_cell_reg[155] <= 0;					r_cell_reg[156] <= 0;					r_cell_reg[157] <= 0;					r_cell_reg[158] <= 0;					r_cell_reg[159] <= 0;					r_cell_reg[160] <= 0;					r_cell_reg[161] <= 0;					r_cell_reg[162] <= 0;					r_cell_reg[163] <= 0;					r_cell_reg[164] <= 0;					r_cell_reg[165] <= 0;					r_cell_reg[166] <= 0;					r_cell_reg[167] <= 0;					r_cell_reg[168] <= 0;					r_cell_reg[169] <= 0;					r_cell_reg[170] <= 0;					r_cell_reg[171] <= 0;					r_cell_reg[172] <= 0;					r_cell_reg[173] <= 0;					r_cell_reg[174] <= 0;					r_cell_reg[175] <= 0;					r_cell_reg[176] <= 0;					r_cell_reg[177] <= 0;					r_cell_reg[178] <= 0;					r_cell_reg[179] <= 0;					r_cell_reg[180] <= 0;					r_cell_reg[181] <= 0;					r_cell_reg[182] <= 0;					r_cell_reg[183] <= 0;					r_cell_reg[184] <= 0;					r_cell_reg[185] <= 0;					r_cell_reg[186] <= 0;					r_cell_reg[187] <= 0;					r_cell_reg[188] <= 0;					r_cell_reg[189] <= 0;					r_cell_reg[190] <= 0;					r_cell_reg[191] <= 0;					r_cell_reg[192] <= 0;					r_cell_reg[193] <= 0;					r_cell_reg[194] <= 0;					r_cell_reg[195] <= 0;					r_cell_reg[196] <= 0;					r_cell_reg[197] <= 0;					r_cell_reg[198] <= 0;					r_cell_reg[199] <= 0;					r_cell_reg[200] <= 0;					r_cell_reg[201] <= 0;					r_cell_reg[202] <= 0;					r_cell_reg[203] <= 0;					r_cell_reg[204] <= 0;					r_cell_reg[205] <= 0;					r_cell_reg[206] <= 0;					r_cell_reg[207] <= 0;					r_cell_reg[208] <= 0;					r_cell_reg[209] <= 0;					r_cell_reg[210] <= 0;					r_cell_reg[211] <= 0;					r_cell_reg[212] <= 0;					r_cell_reg[213] <= 0;					r_cell_reg[214] <= 0;					r_cell_reg[215] <= 0;					r_cell_reg[216] <= 0;					r_cell_reg[217] <= 0;					r_cell_reg[218] <= 0;					r_cell_reg[219] <= 0;					r_cell_reg[220] <= 0;					r_cell_reg[221] <= 0;					r_cell_reg[222] <= 0;					r_cell_reg[223] <= 0;					r_cell_reg[224] <= 0;					r_cell_reg[225] <= 0;					r_cell_reg[226] <= 0;					r_cell_reg[227] <= 0;					r_cell_reg[228] <= 0;					r_cell_reg[229] <= 0;					r_cell_reg[230] <= 0;					r_cell_reg[231] <= 0;					r_cell_reg[232] <= 0;					r_cell_reg[233] <= 0;					r_cell_reg[234] <= 0;					r_cell_reg[235] <= 0;					r_cell_reg[236] <= 0;					r_cell_reg[237] <= 0;					r_cell_reg[238] <= 0;					r_cell_reg[239] <= 0;					r_cell_reg[240] <= 0;					r_cell_reg[241] <= 0;					r_cell_reg[242] <= 0;					r_cell_reg[243] <= 0;					r_cell_reg[244] <= 0;					r_cell_reg[245] <= 0;					r_cell_reg[246] <= 0;					r_cell_reg[247] <= 0;					r_cell_reg[248] <= 0;					r_cell_reg[249] <= 0;					r_cell_reg[250] <= 0;					r_cell_reg[251] <= 0;					r_cell_reg[252] <= 0;					r_cell_reg[253] <= 0;					r_cell_reg[254] <= 0;					r_cell_reg[255] <= 0;					l_cell_reg[0] <= 0;					l_cell_reg[1] <= 0;					l_cell_reg[2] <= 0;					l_cell_reg[3] <= 0;					l_cell_reg[4] <= 0;					l_cell_reg[5] <= 0;					l_cell_reg[6] <= 0;					l_cell_reg[7] <= 0;					l_cell_reg[8] <= 0;					l_cell_reg[9] <= 0;					l_cell_reg[10] <= 0;					l_cell_reg[11] <= 0;					l_cell_reg[12] <= 0;					l_cell_reg[13] <= 0;					l_cell_reg[14] <= 0;					l_cell_reg[15] <= 0;					l_cell_reg[16] <= 0;					l_cell_reg[17] <= 0;					l_cell_reg[18] <= 0;					l_cell_reg[19] <= 0;					l_cell_reg[20] <= 0;					l_cell_reg[21] <= 0;					l_cell_reg[22] <= 0;					l_cell_reg[23] <= 0;					l_cell_reg[24] <= 0;					l_cell_reg[25] <= 0;					l_cell_reg[26] <= 0;					l_cell_reg[27] <= 0;					l_cell_reg[28] <= 0;					l_cell_reg[29] <= 0;					l_cell_reg[30] <= 0;					l_cell_reg[31] <= 0;					l_cell_reg[32] <= 0;					l_cell_reg[33] <= 0;					l_cell_reg[34] <= 0;					l_cell_reg[35] <= 0;					l_cell_reg[36] <= 0;					l_cell_reg[37] <= 0;					l_cell_reg[38] <= 0;					l_cell_reg[39] <= 0;					l_cell_reg[40] <= 0;					l_cell_reg[41] <= 0;					l_cell_reg[42] <= 0;					l_cell_reg[43] <= 0;					l_cell_reg[44] <= 0;					l_cell_reg[45] <= 0;					l_cell_reg[46] <= 0;					l_cell_reg[47] <= 0;					l_cell_reg[48] <= 0;					l_cell_reg[49] <= 0;					l_cell_reg[50] <= 0;					l_cell_reg[51] <= 0;					l_cell_reg[52] <= 0;					l_cell_reg[53] <= 0;					l_cell_reg[54] <= 0;					l_cell_reg[55] <= 0;					l_cell_reg[56] <= 0;					l_cell_reg[57] <= 0;					l_cell_reg[58] <= 0;					l_cell_reg[59] <= 0;					l_cell_reg[60] <= 0;					l_cell_reg[61] <= 0;					l_cell_reg[62] <= 0;					l_cell_reg[63] <= 0;					l_cell_reg[64] <= 0;					l_cell_reg[65] <= 0;					l_cell_reg[66] <= 0;					l_cell_reg[67] <= 0;					l_cell_reg[68] <= 0;					l_cell_reg[69] <= 0;					l_cell_reg[70] <= 0;					l_cell_reg[71] <= 0;					l_cell_reg[72] <= 0;					l_cell_reg[73] <= 0;					l_cell_reg[74] <= 0;					l_cell_reg[75] <= 0;					l_cell_reg[76] <= 0;					l_cell_reg[77] <= 0;					l_cell_reg[78] <= 0;					l_cell_reg[79] <= 0;					l_cell_reg[80] <= 0;					l_cell_reg[81] <= 0;					l_cell_reg[82] <= 0;					l_cell_reg[83] <= 0;					l_cell_reg[84] <= 0;					l_cell_reg[85] <= 0;					l_cell_reg[86] <= 0;					l_cell_reg[87] <= 0;					l_cell_reg[88] <= 0;					l_cell_reg[89] <= 0;					l_cell_reg[90] <= 0;					l_cell_reg[91] <= 0;					l_cell_reg[92] <= 0;					l_cell_reg[93] <= 0;					l_cell_reg[94] <= 0;					l_cell_reg[95] <= 0;					l_cell_reg[96] <= 0;					l_cell_reg[97] <= 0;					l_cell_reg[98] <= 0;					l_cell_reg[99] <= 0;					l_cell_reg[100] <= 0;					l_cell_reg[101] <= 0;					l_cell_reg[102] <= 0;					l_cell_reg[103] <= 0;					l_cell_reg[104] <= 0;					l_cell_reg[105] <= 0;					l_cell_reg[106] <= 0;					l_cell_reg[107] <= 0;					l_cell_reg[108] <= 0;					l_cell_reg[109] <= 0;					l_cell_reg[110] <= 0;					l_cell_reg[111] <= 0;					l_cell_reg[112] <= 0;					l_cell_reg[113] <= 0;					l_cell_reg[114] <= 0;					l_cell_reg[115] <= 0;					l_cell_reg[116] <= 0;					l_cell_reg[117] <= 0;					l_cell_reg[118] <= 0;					l_cell_reg[119] <= 0;					l_cell_reg[120] <= 0;					l_cell_reg[121] <= 0;					l_cell_reg[122] <= 0;					l_cell_reg[123] <= 0;					l_cell_reg[124] <= 0;					l_cell_reg[125] <= 0;					l_cell_reg[126] <= 0;					l_cell_reg[127] <= 0;					l_cell_reg[128] <= 0;					l_cell_reg[129] <= 0;					l_cell_reg[130] <= 0;					l_cell_reg[131] <= 0;					l_cell_reg[132] <= 0;					l_cell_reg[133] <= 0;					l_cell_reg[134] <= 0;					l_cell_reg[135] <= 0;					l_cell_reg[136] <= 0;					l_cell_reg[137] <= 0;					l_cell_reg[138] <= 0;					l_cell_reg[139] <= 0;					l_cell_reg[140] <= 0;					l_cell_reg[141] <= 0;					l_cell_reg[142] <= 0;					l_cell_reg[143] <= 0;					l_cell_reg[144] <= 0;					l_cell_reg[145] <= 0;					l_cell_reg[146] <= 0;					l_cell_reg[147] <= 0;					l_cell_reg[148] <= 0;					l_cell_reg[149] <= 0;					l_cell_reg[150] <= 0;					l_cell_reg[151] <= 0;					l_cell_reg[152] <= 0;					l_cell_reg[153] <= 0;					l_cell_reg[154] <= 0;					l_cell_reg[155] <= 0;					l_cell_reg[156] <= 0;					l_cell_reg[157] <= 0;					l_cell_reg[158] <= 0;					l_cell_reg[159] <= 0;					l_cell_reg[160] <= 0;					l_cell_reg[161] <= 0;					l_cell_reg[162] <= 0;					l_cell_reg[163] <= 0;					l_cell_reg[164] <= 0;					l_cell_reg[165] <= 0;					l_cell_reg[166] <= 0;					l_cell_reg[167] <= 0;					l_cell_reg[168] <= 0;					l_cell_reg[169] <= 0;					l_cell_reg[170] <= 0;					l_cell_reg[171] <= 0;					l_cell_reg[172] <= 0;					l_cell_reg[173] <= 0;					l_cell_reg[174] <= 0;					l_cell_reg[175] <= 0;					l_cell_reg[176] <= 0;					l_cell_reg[177] <= 0;					l_cell_reg[178] <= 0;					l_cell_reg[179] <= 0;					l_cell_reg[180] <= 0;					l_cell_reg[181] <= 0;					l_cell_reg[182] <= 0;					l_cell_reg[183] <= 0;					l_cell_reg[184] <= 0;					l_cell_reg[185] <= 0;					l_cell_reg[186] <= 0;					l_cell_reg[187] <= 0;					l_cell_reg[188] <= 0;					l_cell_reg[189] <= 0;					l_cell_reg[190] <= 0;					l_cell_reg[191] <= 0;					l_cell_reg[192] <= 0;					l_cell_reg[193] <= 0;					l_cell_reg[194] <= 0;					l_cell_reg[195] <= 0;					l_cell_reg[196] <= 0;					l_cell_reg[197] <= 0;					l_cell_reg[198] <= 0;					l_cell_reg[199] <= 0;					l_cell_reg[200] <= 0;					l_cell_reg[201] <= 0;					l_cell_reg[202] <= 0;					l_cell_reg[203] <= 0;					l_cell_reg[204] <= 0;					l_cell_reg[205] <= 0;					l_cell_reg[206] <= 0;					l_cell_reg[207] <= 0;					l_cell_reg[208] <= 0;					l_cell_reg[209] <= 0;					l_cell_reg[210] <= 0;					l_cell_reg[211] <= 0;					l_cell_reg[212] <= 0;					l_cell_reg[213] <= 0;					l_cell_reg[214] <= 0;					l_cell_reg[215] <= 0;					l_cell_reg[216] <= 0;					l_cell_reg[217] <= 0;					l_cell_reg[218] <= 0;					l_cell_reg[219] <= 0;					l_cell_reg[220] <= 0;					l_cell_reg[221] <= 0;					l_cell_reg[222] <= 0;					l_cell_reg[223] <= 0;					l_cell_reg[224] <= 0;					l_cell_reg[225] <= 0;					l_cell_reg[226] <= 0;					l_cell_reg[227] <= 0;					l_cell_reg[228] <= 0;					l_cell_reg[229] <= 0;					l_cell_reg[230] <= 0;					l_cell_reg[231] <= 0;					l_cell_reg[232] <= 0;					l_cell_reg[233] <= 0;					l_cell_reg[234] <= 0;					l_cell_reg[235] <= 0;					l_cell_reg[236] <= 0;					l_cell_reg[237] <= 0;					l_cell_reg[238] <= 0;					l_cell_reg[239] <= 0;					l_cell_reg[240] <= 0;					l_cell_reg[241] <= 0;					l_cell_reg[242] <= 0;					l_cell_reg[243] <= 0;					l_cell_reg[244] <= 0;					l_cell_reg[245] <= 0;					l_cell_reg[246] <= 0;					l_cell_reg[247] <= 0;					l_cell_reg[248] <= 0;					l_cell_reg[249] <= 0;					l_cell_reg[250] <= 0;					l_cell_reg[251] <= 0;					l_cell_reg[252] <= 0;					l_cell_reg[253] <= 0;					l_cell_reg[254] <= 0;					l_cell_reg[255] <= 0;			end
		endcase	end
	genvar i;	generate		for (i = 0; i < 256 ; i = i+2)			begin :bp_2				bp_2_cell fun(					.clk(clk),					.en(1),					.R_IN1(r_cell_reg[i]),					.R_IN2(r_cell_reg[i+1]),					.L_IN1(l_cell_reg[i]),					.L_IN2(l_cell_reg[i+1]),					.R_OUT1(r_cell_wire[i]),					.R_OUT2(r_cell_wire[i+1]),					.L_OUT1(l_cell_wire[i]),					.L_OUT2(l_cell_wire[i+1])				);			end	endgenerate
	always @(posedge clk) begin		if (bp_over_flag) begin			OUT_1 <= inform_L [0][0] ;			OUT_2 <= inform_L [1][0] ;			OUT_3 <= inform_L [2][0] ;			OUT_4 <= inform_L [3][0] ;			OUT_5 <= inform_L [4][0] ;			OUT_6 <= inform_L [5][0] ;			OUT_7 <= inform_L [6][0] ;			OUT_8 <= inform_L [7][0] ;			OUT_9 <= inform_L [8][0] ;			OUT_10 <= inform_L [9][0] ;			OUT_11 <= inform_L [10][0] ;			OUT_12 <= inform_L [11][0] ;			OUT_13 <= inform_L [12][0] ;			OUT_14 <= inform_L [13][0] ;			OUT_15 <= inform_L [14][0] ;			OUT_16 <= inform_L [15][0] ;			OUT_17 <= inform_L [16][0] ;			OUT_18 <= inform_L [17][0] ;			OUT_19 <= inform_L [18][0] ;			OUT_20 <= inform_L [19][0] ;			OUT_21 <= inform_L [20][0] ;			OUT_22 <= inform_L [21][0] ;			OUT_23 <= inform_L [22][0] ;			OUT_24 <= inform_L [23][0] ;			OUT_25 <= inform_L [24][0] ;			OUT_26 <= inform_L [25][0] ;			OUT_27 <= inform_L [26][0] ;			OUT_28 <= inform_L [27][0] ;			OUT_29 <= inform_L [28][0] ;			OUT_30 <= inform_L [29][0] ;			OUT_31 <= inform_L [30][0] ;			OUT_32 <= inform_L [31][0] ;			OUT_33 <= inform_L [32][0] ;			OUT_34 <= inform_L [33][0] ;			OUT_35 <= inform_L [34][0] ;			OUT_36 <= inform_L [35][0] ;			OUT_37 <= inform_L [36][0] ;			OUT_38 <= inform_L [37][0] ;			OUT_39 <= inform_L [38][0] ;			OUT_40 <= inform_L [39][0] ;			OUT_41 <= inform_L [40][0] ;			OUT_42 <= inform_L [41][0] ;			OUT_43 <= inform_L [42][0] ;			OUT_44 <= inform_L [43][0] ;			OUT_45 <= inform_L [44][0] ;			OUT_46 <= inform_L [45][0] ;			OUT_47 <= inform_L [46][0] ;			OUT_48 <= inform_L [47][0] ;			OUT_49 <= inform_L [48][0] ;			OUT_50 <= inform_L [49][0] ;			OUT_51 <= inform_L [50][0] ;			OUT_52 <= inform_L [51][0] ;			OUT_53 <= inform_L [52][0] ;			OUT_54 <= inform_L [53][0] ;			OUT_55 <= inform_L [54][0] ;			OUT_56 <= inform_L [55][0] ;			OUT_57 <= inform_L [56][0] ;			OUT_58 <= inform_L [57][0] ;			OUT_59 <= inform_L [58][0] ;			OUT_60 <= inform_L [59][0] ;			OUT_61 <= inform_L [60][0] ;			OUT_62 <= inform_L [61][0] ;			OUT_63 <= inform_L [62][0] ;			OUT_64 <= inform_L [63][0] ;			OUT_65 <= inform_L [64][0] ;			OUT_66 <= inform_L [65][0] ;			OUT_67 <= inform_L [66][0] ;			OUT_68 <= inform_L [67][0] ;			OUT_69 <= inform_L [68][0] ;			OUT_70 <= inform_L [69][0] ;			OUT_71 <= inform_L [70][0] ;			OUT_72 <= inform_L [71][0] ;			OUT_73 <= inform_L [72][0] ;			OUT_74 <= inform_L [73][0] ;			OUT_75 <= inform_L [74][0] ;			OUT_76 <= inform_L [75][0] ;			OUT_77 <= inform_L [76][0] ;			OUT_78 <= inform_L [77][0] ;			OUT_79 <= inform_L [78][0] ;			OUT_80 <= inform_L [79][0] ;			OUT_81 <= inform_L [80][0] ;			OUT_82 <= inform_L [81][0] ;			OUT_83 <= inform_L [82][0] ;			OUT_84 <= inform_L [83][0] ;			OUT_85 <= inform_L [84][0] ;			OUT_86 <= inform_L [85][0] ;			OUT_87 <= inform_L [86][0] ;			OUT_88 <= inform_L [87][0] ;			OUT_89 <= inform_L [88][0] ;			OUT_90 <= inform_L [89][0] ;			OUT_91 <= inform_L [90][0] ;			OUT_92 <= inform_L [91][0] ;			OUT_93 <= inform_L [92][0] ;			OUT_94 <= inform_L [93][0] ;			OUT_95 <= inform_L [94][0] ;			OUT_96 <= inform_L [95][0] ;			OUT_97 <= inform_L [96][0] ;			OUT_98 <= inform_L [97][0] ;			OUT_99 <= inform_L [98][0] ;			OUT_100 <= inform_L [99][0] ;			OUT_101 <= inform_L [100][0] ;			OUT_102 <= inform_L [101][0] ;			OUT_103 <= inform_L [102][0] ;			OUT_104 <= inform_L [103][0] ;			OUT_105 <= inform_L [104][0] ;			OUT_106 <= inform_L [105][0] ;			OUT_107 <= inform_L [106][0] ;			OUT_108 <= inform_L [107][0] ;			OUT_109 <= inform_L [108][0] ;			OUT_110 <= inform_L [109][0] ;			OUT_111 <= inform_L [110][0] ;			OUT_112 <= inform_L [111][0] ;			OUT_113 <= inform_L [112][0] ;			OUT_114 <= inform_L [113][0] ;			OUT_115 <= inform_L [114][0] ;			OUT_116 <= inform_L [115][0] ;			OUT_117 <= inform_L [116][0] ;			OUT_118 <= inform_L [117][0] ;			OUT_119 <= inform_L [118][0] ;			OUT_120 <= inform_L [119][0] ;			OUT_121 <= inform_L [120][0] ;			OUT_122 <= inform_L [121][0] ;			OUT_123 <= inform_L [122][0] ;			OUT_124 <= inform_L [123][0] ;			OUT_125 <= inform_L [124][0] ;			OUT_126 <= inform_L [125][0] ;			OUT_127 <= inform_L [126][0] ;			OUT_128 <= inform_L [127][0] ;			OUT_129 <= inform_L [128][0] ;			OUT_130 <= inform_L [129][0] ;			OUT_131 <= inform_L [130][0] ;			OUT_132 <= inform_L [131][0] ;			OUT_133 <= inform_L [132][0] ;			OUT_134 <= inform_L [133][0] ;			OUT_135 <= inform_L [134][0] ;			OUT_136 <= inform_L [135][0] ;			OUT_137 <= inform_L [136][0] ;			OUT_138 <= inform_L [137][0] ;			OUT_139 <= inform_L [138][0] ;			OUT_140 <= inform_L [139][0] ;			OUT_141 <= inform_L [140][0] ;			OUT_142 <= inform_L [141][0] ;			OUT_143 <= inform_L [142][0] ;			OUT_144 <= inform_L [143][0] ;			OUT_145 <= inform_L [144][0] ;			OUT_146 <= inform_L [145][0] ;			OUT_147 <= inform_L [146][0] ;			OUT_148 <= inform_L [147][0] ;			OUT_149 <= inform_L [148][0] ;			OUT_150 <= inform_L [149][0] ;			OUT_151 <= inform_L [150][0] ;			OUT_152 <= inform_L [151][0] ;			OUT_153 <= inform_L [152][0] ;			OUT_154 <= inform_L [153][0] ;			OUT_155 <= inform_L [154][0] ;			OUT_156 <= inform_L [155][0] ;			OUT_157 <= inform_L [156][0] ;			OUT_158 <= inform_L [157][0] ;			OUT_159 <= inform_L [158][0] ;			OUT_160 <= inform_L [159][0] ;			OUT_161 <= inform_L [160][0] ;			OUT_162 <= inform_L [161][0] ;			OUT_163 <= inform_L [162][0] ;			OUT_164 <= inform_L [163][0] ;			OUT_165 <= inform_L [164][0] ;			OUT_166 <= inform_L [165][0] ;			OUT_167 <= inform_L [166][0] ;			OUT_168 <= inform_L [167][0] ;			OUT_169 <= inform_L [168][0] ;			OUT_170 <= inform_L [169][0] ;			OUT_171 <= inform_L [170][0] ;			OUT_172 <= inform_L [171][0] ;			OUT_173 <= inform_L [172][0] ;			OUT_174 <= inform_L [173][0] ;			OUT_175 <= inform_L [174][0] ;			OUT_176 <= inform_L [175][0] ;			OUT_177 <= inform_L [176][0] ;			OUT_178 <= inform_L [177][0] ;			OUT_179 <= inform_L [178][0] ;			OUT_180 <= inform_L [179][0] ;			OUT_181 <= inform_L [180][0] ;			OUT_182 <= inform_L [181][0] ;			OUT_183 <= inform_L [182][0] ;			OUT_184 <= inform_L [183][0] ;			OUT_185 <= inform_L [184][0] ;			OUT_186 <= inform_L [185][0] ;			OUT_187 <= inform_L [186][0] ;			OUT_188 <= inform_L [187][0] ;			OUT_189 <= inform_L [188][0] ;			OUT_190 <= inform_L [189][0] ;			OUT_191 <= inform_L [190][0] ;			OUT_192 <= inform_L [191][0] ;			OUT_193 <= inform_L [192][0] ;			OUT_194 <= inform_L [193][0] ;			OUT_195 <= inform_L [194][0] ;			OUT_196 <= inform_L [195][0] ;			OUT_197 <= inform_L [196][0] ;			OUT_198 <= inform_L [197][0] ;			OUT_199 <= inform_L [198][0] ;			OUT_200 <= inform_L [199][0] ;			OUT_201 <= inform_L [200][0] ;			OUT_202 <= inform_L [201][0] ;			OUT_203 <= inform_L [202][0] ;			OUT_204 <= inform_L [203][0] ;			OUT_205 <= inform_L [204][0] ;			OUT_206 <= inform_L [205][0] ;			OUT_207 <= inform_L [206][0] ;			OUT_208 <= inform_L [207][0] ;			OUT_209 <= inform_L [208][0] ;			OUT_210 <= inform_L [209][0] ;			OUT_211 <= inform_L [210][0] ;			OUT_212 <= inform_L [211][0] ;			OUT_213 <= inform_L [212][0] ;			OUT_214 <= inform_L [213][0] ;			OUT_215 <= inform_L [214][0] ;			OUT_216 <= inform_L [215][0] ;			OUT_217 <= inform_L [216][0] ;			OUT_218 <= inform_L [217][0] ;			OUT_219 <= inform_L [218][0] ;			OUT_220 <= inform_L [219][0] ;			OUT_221 <= inform_L [220][0] ;			OUT_222 <= inform_L [221][0] ;			OUT_223 <= inform_L [222][0] ;			OUT_224 <= inform_L [223][0] ;			OUT_225 <= inform_L [224][0] ;			OUT_226 <= inform_L [225][0] ;			OUT_227 <= inform_L [226][0] ;			OUT_228 <= inform_L [227][0] ;			OUT_229 <= inform_L [228][0] ;			OUT_230 <= inform_L [229][0] ;			OUT_231 <= inform_L [230][0] ;			OUT_232 <= inform_L [231][0] ;			OUT_233 <= inform_L [232][0] ;			OUT_234 <= inform_L [233][0] ;			OUT_235 <= inform_L [234][0] ;			OUT_236 <= inform_L [235][0] ;			OUT_237 <= inform_L [236][0] ;			OUT_238 <= inform_L [237][0] ;			OUT_239 <= inform_L [238][0] ;			OUT_240 <= inform_L [239][0] ;			OUT_241 <= inform_L [240][0] ;			OUT_242 <= inform_L [241][0] ;			OUT_243 <= inform_L [242][0] ;			OUT_244 <= inform_L [243][0] ;			OUT_245 <= inform_L [244][0] ;			OUT_246 <= inform_L [245][0] ;			OUT_247 <= inform_L [246][0] ;			OUT_248 <= inform_L [247][0] ;			OUT_249 <= inform_L [248][0] ;			OUT_250 <= inform_L [249][0] ;			OUT_251 <= inform_L [250][0] ;			OUT_252 <= inform_L [251][0] ;			OUT_253 <= inform_L [252][0] ;			OUT_254 <= inform_L [253][0] ;			OUT_255 <= inform_L [254][0] ;			OUT_256 <= inform_L [255][0] ;		end	end
endmodule