`define iteration_times 40 module bp_1024_720 #(	parameter integer BIT = 8)(	input clk,	input rst_n,	input start,	output reg en_busy,	input [BIT - 1:0] LLR_1,	input [BIT - 1:0] LLR_2,	input [BIT - 1:0] LLR_3,	input [BIT - 1:0] LLR_4,	input [BIT - 1:0] LLR_5,	input [BIT - 1:0] LLR_6,	input [BIT - 1:0] LLR_7,	input [BIT - 1:0] LLR_8,	input [BIT - 1:0] LLR_9,	input [BIT - 1:0] LLR_10,	input [BIT - 1:0] LLR_11,	input [BIT - 1:0] LLR_12,	input [BIT - 1:0] LLR_13,	input [BIT - 1:0] LLR_14,	input [BIT - 1:0] LLR_15,	input [BIT - 1:0] LLR_16,	input [BIT - 1:0] LLR_17,	input [BIT - 1:0] LLR_18,	input [BIT - 1:0] LLR_19,	input [BIT - 1:0] LLR_20,	input [BIT - 1:0] LLR_21,	input [BIT - 1:0] LLR_22,	input [BIT - 1:0] LLR_23,	input [BIT - 1:0] LLR_24,	input [BIT - 1:0] LLR_25,	input [BIT - 1:0] LLR_26,	input [BIT - 1:0] LLR_27,	input [BIT - 1:0] LLR_28,	input [BIT - 1:0] LLR_29,	input [BIT - 1:0] LLR_30,	input [BIT - 1:0] LLR_31,	input [BIT - 1:0] LLR_32,	input [BIT - 1:0] LLR_33,	input [BIT - 1:0] LLR_34,	input [BIT - 1:0] LLR_35,	input [BIT - 1:0] LLR_36,	input [BIT - 1:0] LLR_37,	input [BIT - 1:0] LLR_38,	input [BIT - 1:0] LLR_39,	input [BIT - 1:0] LLR_40,	input [BIT - 1:0] LLR_41,	input [BIT - 1:0] LLR_42,	input [BIT - 1:0] LLR_43,	input [BIT - 1:0] LLR_44,	input [BIT - 1:0] LLR_45,	input [BIT - 1:0] LLR_46,	input [BIT - 1:0] LLR_47,	input [BIT - 1:0] LLR_48,	input [BIT - 1:0] LLR_49,	input [BIT - 1:0] LLR_50,	input [BIT - 1:0] LLR_51,	input [BIT - 1:0] LLR_52,	input [BIT - 1:0] LLR_53,	input [BIT - 1:0] LLR_54,	input [BIT - 1:0] LLR_55,	input [BIT - 1:0] LLR_56,	input [BIT - 1:0] LLR_57,	input [BIT - 1:0] LLR_58,	input [BIT - 1:0] LLR_59,	input [BIT - 1:0] LLR_60,	input [BIT - 1:0] LLR_61,	input [BIT - 1:0] LLR_62,	input [BIT - 1:0] LLR_63,	input [BIT - 1:0] LLR_64,	input [BIT - 1:0] LLR_65,	input [BIT - 1:0] LLR_66,	input [BIT - 1:0] LLR_67,	input [BIT - 1:0] LLR_68,	input [BIT - 1:0] LLR_69,	input [BIT - 1:0] LLR_70,	input [BIT - 1:0] LLR_71,	input [BIT - 1:0] LLR_72,	input [BIT - 1:0] LLR_73,	input [BIT - 1:0] LLR_74,	input [BIT - 1:0] LLR_75,	input [BIT - 1:0] LLR_76,	input [BIT - 1:0] LLR_77,	input [BIT - 1:0] LLR_78,	input [BIT - 1:0] LLR_79,	input [BIT - 1:0] LLR_80,	input [BIT - 1:0] LLR_81,	input [BIT - 1:0] LLR_82,	input [BIT - 1:0] LLR_83,	input [BIT - 1:0] LLR_84,	input [BIT - 1:0] LLR_85,	input [BIT - 1:0] LLR_86,	input [BIT - 1:0] LLR_87,	input [BIT - 1:0] LLR_88,	input [BIT - 1:0] LLR_89,	input [BIT - 1:0] LLR_90,	input [BIT - 1:0] LLR_91,	input [BIT - 1:0] LLR_92,	input [BIT - 1:0] LLR_93,	input [BIT - 1:0] LLR_94,	input [BIT - 1:0] LLR_95,	input [BIT - 1:0] LLR_96,	input [BIT - 1:0] LLR_97,	input [BIT - 1:0] LLR_98,	input [BIT - 1:0] LLR_99,	input [BIT - 1:0] LLR_100,	input [BIT - 1:0] LLR_101,	input [BIT - 1:0] LLR_102,	input [BIT - 1:0] LLR_103,	input [BIT - 1:0] LLR_104,	input [BIT - 1:0] LLR_105,	input [BIT - 1:0] LLR_106,	input [BIT - 1:0] LLR_107,	input [BIT - 1:0] LLR_108,	input [BIT - 1:0] LLR_109,	input [BIT - 1:0] LLR_110,	input [BIT - 1:0] LLR_111,	input [BIT - 1:0] LLR_112,	input [BIT - 1:0] LLR_113,	input [BIT - 1:0] LLR_114,	input [BIT - 1:0] LLR_115,	input [BIT - 1:0] LLR_116,	input [BIT - 1:0] LLR_117,	input [BIT - 1:0] LLR_118,	input [BIT - 1:0] LLR_119,	input [BIT - 1:0] LLR_120,	input [BIT - 1:0] LLR_121,	input [BIT - 1:0] LLR_122,	input [BIT - 1:0] LLR_123,	input [BIT - 1:0] LLR_124,	input [BIT - 1:0] LLR_125,	input [BIT - 1:0] LLR_126,	input [BIT - 1:0] LLR_127,	input [BIT - 1:0] LLR_128,	input [BIT - 1:0] LLR_129,	input [BIT - 1:0] LLR_130,	input [BIT - 1:0] LLR_131,	input [BIT - 1:0] LLR_132,	input [BIT - 1:0] LLR_133,	input [BIT - 1:0] LLR_134,	input [BIT - 1:0] LLR_135,	input [BIT - 1:0] LLR_136,	input [BIT - 1:0] LLR_137,	input [BIT - 1:0] LLR_138,	input [BIT - 1:0] LLR_139,	input [BIT - 1:0] LLR_140,	input [BIT - 1:0] LLR_141,	input [BIT - 1:0] LLR_142,	input [BIT - 1:0] LLR_143,	input [BIT - 1:0] LLR_144,	input [BIT - 1:0] LLR_145,	input [BIT - 1:0] LLR_146,	input [BIT - 1:0] LLR_147,	input [BIT - 1:0] LLR_148,	input [BIT - 1:0] LLR_149,	input [BIT - 1:0] LLR_150,	input [BIT - 1:0] LLR_151,	input [BIT - 1:0] LLR_152,	input [BIT - 1:0] LLR_153,	input [BIT - 1:0] LLR_154,	input [BIT - 1:0] LLR_155,	input [BIT - 1:0] LLR_156,	input [BIT - 1:0] LLR_157,	input [BIT - 1:0] LLR_158,	input [BIT - 1:0] LLR_159,	input [BIT - 1:0] LLR_160,	input [BIT - 1:0] LLR_161,	input [BIT - 1:0] LLR_162,	input [BIT - 1:0] LLR_163,	input [BIT - 1:0] LLR_164,	input [BIT - 1:0] LLR_165,	input [BIT - 1:0] LLR_166,	input [BIT - 1:0] LLR_167,	input [BIT - 1:0] LLR_168,	input [BIT - 1:0] LLR_169,	input [BIT - 1:0] LLR_170,	input [BIT - 1:0] LLR_171,	input [BIT - 1:0] LLR_172,	input [BIT - 1:0] LLR_173,	input [BIT - 1:0] LLR_174,	input [BIT - 1:0] LLR_175,	input [BIT - 1:0] LLR_176,	input [BIT - 1:0] LLR_177,	input [BIT - 1:0] LLR_178,	input [BIT - 1:0] LLR_179,	input [BIT - 1:0] LLR_180,	input [BIT - 1:0] LLR_181,	input [BIT - 1:0] LLR_182,	input [BIT - 1:0] LLR_183,	input [BIT - 1:0] LLR_184,	input [BIT - 1:0] LLR_185,	input [BIT - 1:0] LLR_186,	input [BIT - 1:0] LLR_187,	input [BIT - 1:0] LLR_188,	input [BIT - 1:0] LLR_189,	input [BIT - 1:0] LLR_190,	input [BIT - 1:0] LLR_191,	input [BIT - 1:0] LLR_192,	input [BIT - 1:0] LLR_193,	input [BIT - 1:0] LLR_194,	input [BIT - 1:0] LLR_195,	input [BIT - 1:0] LLR_196,	input [BIT - 1:0] LLR_197,	input [BIT - 1:0] LLR_198,	input [BIT - 1:0] LLR_199,	input [BIT - 1:0] LLR_200,	input [BIT - 1:0] LLR_201,	input [BIT - 1:0] LLR_202,	input [BIT - 1:0] LLR_203,	input [BIT - 1:0] LLR_204,	input [BIT - 1:0] LLR_205,	input [BIT - 1:0] LLR_206,	input [BIT - 1:0] LLR_207,	input [BIT - 1:0] LLR_208,	input [BIT - 1:0] LLR_209,	input [BIT - 1:0] LLR_210,	input [BIT - 1:0] LLR_211,	input [BIT - 1:0] LLR_212,	input [BIT - 1:0] LLR_213,	input [BIT - 1:0] LLR_214,	input [BIT - 1:0] LLR_215,	input [BIT - 1:0] LLR_216,	input [BIT - 1:0] LLR_217,	input [BIT - 1:0] LLR_218,	input [BIT - 1:0] LLR_219,	input [BIT - 1:0] LLR_220,	input [BIT - 1:0] LLR_221,	input [BIT - 1:0] LLR_222,	input [BIT - 1:0] LLR_223,	input [BIT - 1:0] LLR_224,	input [BIT - 1:0] LLR_225,	input [BIT - 1:0] LLR_226,	input [BIT - 1:0] LLR_227,	input [BIT - 1:0] LLR_228,	input [BIT - 1:0] LLR_229,	input [BIT - 1:0] LLR_230,	input [BIT - 1:0] LLR_231,	input [BIT - 1:0] LLR_232,	input [BIT - 1:0] LLR_233,	input [BIT - 1:0] LLR_234,	input [BIT - 1:0] LLR_235,	input [BIT - 1:0] LLR_236,	input [BIT - 1:0] LLR_237,	input [BIT - 1:0] LLR_238,	input [BIT - 1:0] LLR_239,	input [BIT - 1:0] LLR_240,	input [BIT - 1:0] LLR_241,	input [BIT - 1:0] LLR_242,	input [BIT - 1:0] LLR_243,	input [BIT - 1:0] LLR_244,	input [BIT - 1:0] LLR_245,	input [BIT - 1:0] LLR_246,	input [BIT - 1:0] LLR_247,	input [BIT - 1:0] LLR_248,	input [BIT - 1:0] LLR_249,	input [BIT - 1:0] LLR_250,	input [BIT - 1:0] LLR_251,	input [BIT - 1:0] LLR_252,	input [BIT - 1:0] LLR_253,	input [BIT - 1:0] LLR_254,	input [BIT - 1:0] LLR_255,	input [BIT - 1:0] LLR_256,	input [BIT - 1:0] LLR_257,	input [BIT - 1:0] LLR_258,	input [BIT - 1:0] LLR_259,	input [BIT - 1:0] LLR_260,	input [BIT - 1:0] LLR_261,	input [BIT - 1:0] LLR_262,	input [BIT - 1:0] LLR_263,	input [BIT - 1:0] LLR_264,	input [BIT - 1:0] LLR_265,	input [BIT - 1:0] LLR_266,	input [BIT - 1:0] LLR_267,	input [BIT - 1:0] LLR_268,	input [BIT - 1:0] LLR_269,	input [BIT - 1:0] LLR_270,	input [BIT - 1:0] LLR_271,	input [BIT - 1:0] LLR_272,	input [BIT - 1:0] LLR_273,	input [BIT - 1:0] LLR_274,	input [BIT - 1:0] LLR_275,	input [BIT - 1:0] LLR_276,	input [BIT - 1:0] LLR_277,	input [BIT - 1:0] LLR_278,	input [BIT - 1:0] LLR_279,	input [BIT - 1:0] LLR_280,	input [BIT - 1:0] LLR_281,	input [BIT - 1:0] LLR_282,	input [BIT - 1:0] LLR_283,	input [BIT - 1:0] LLR_284,	input [BIT - 1:0] LLR_285,	input [BIT - 1:0] LLR_286,	input [BIT - 1:0] LLR_287,	input [BIT - 1:0] LLR_288,	input [BIT - 1:0] LLR_289,	input [BIT - 1:0] LLR_290,	input [BIT - 1:0] LLR_291,	input [BIT - 1:0] LLR_292,	input [BIT - 1:0] LLR_293,	input [BIT - 1:0] LLR_294,	input [BIT - 1:0] LLR_295,	input [BIT - 1:0] LLR_296,	input [BIT - 1:0] LLR_297,	input [BIT - 1:0] LLR_298,	input [BIT - 1:0] LLR_299,	input [BIT - 1:0] LLR_300,	input [BIT - 1:0] LLR_301,	input [BIT - 1:0] LLR_302,	input [BIT - 1:0] LLR_303,	input [BIT - 1:0] LLR_304,	input [BIT - 1:0] LLR_305,	input [BIT - 1:0] LLR_306,	input [BIT - 1:0] LLR_307,	input [BIT - 1:0] LLR_308,	input [BIT - 1:0] LLR_309,	input [BIT - 1:0] LLR_310,	input [BIT - 1:0] LLR_311,	input [BIT - 1:0] LLR_312,	input [BIT - 1:0] LLR_313,	input [BIT - 1:0] LLR_314,	input [BIT - 1:0] LLR_315,	input [BIT - 1:0] LLR_316,	input [BIT - 1:0] LLR_317,	input [BIT - 1:0] LLR_318,	input [BIT - 1:0] LLR_319,	input [BIT - 1:0] LLR_320,	input [BIT - 1:0] LLR_321,	input [BIT - 1:0] LLR_322,	input [BIT - 1:0] LLR_323,	input [BIT - 1:0] LLR_324,	input [BIT - 1:0] LLR_325,	input [BIT - 1:0] LLR_326,	input [BIT - 1:0] LLR_327,	input [BIT - 1:0] LLR_328,	input [BIT - 1:0] LLR_329,	input [BIT - 1:0] LLR_330,	input [BIT - 1:0] LLR_331,	input [BIT - 1:0] LLR_332,	input [BIT - 1:0] LLR_333,	input [BIT - 1:0] LLR_334,	input [BIT - 1:0] LLR_335,	input [BIT - 1:0] LLR_336,	input [BIT - 1:0] LLR_337,	input [BIT - 1:0] LLR_338,	input [BIT - 1:0] LLR_339,	input [BIT - 1:0] LLR_340,	input [BIT - 1:0] LLR_341,	input [BIT - 1:0] LLR_342,	input [BIT - 1:0] LLR_343,	input [BIT - 1:0] LLR_344,	input [BIT - 1:0] LLR_345,	input [BIT - 1:0] LLR_346,	input [BIT - 1:0] LLR_347,	input [BIT - 1:0] LLR_348,	input [BIT - 1:0] LLR_349,	input [BIT - 1:0] LLR_350,	input [BIT - 1:0] LLR_351,	input [BIT - 1:0] LLR_352,	input [BIT - 1:0] LLR_353,	input [BIT - 1:0] LLR_354,	input [BIT - 1:0] LLR_355,	input [BIT - 1:0] LLR_356,	input [BIT - 1:0] LLR_357,	input [BIT - 1:0] LLR_358,	input [BIT - 1:0] LLR_359,	input [BIT - 1:0] LLR_360,	input [BIT - 1:0] LLR_361,	input [BIT - 1:0] LLR_362,	input [BIT - 1:0] LLR_363,	input [BIT - 1:0] LLR_364,	input [BIT - 1:0] LLR_365,	input [BIT - 1:0] LLR_366,	input [BIT - 1:0] LLR_367,	input [BIT - 1:0] LLR_368,	input [BIT - 1:0] LLR_369,	input [BIT - 1:0] LLR_370,	input [BIT - 1:0] LLR_371,	input [BIT - 1:0] LLR_372,	input [BIT - 1:0] LLR_373,	input [BIT - 1:0] LLR_374,	input [BIT - 1:0] LLR_375,	input [BIT - 1:0] LLR_376,	input [BIT - 1:0] LLR_377,	input [BIT - 1:0] LLR_378,	input [BIT - 1:0] LLR_379,	input [BIT - 1:0] LLR_380,	input [BIT - 1:0] LLR_381,	input [BIT - 1:0] LLR_382,	input [BIT - 1:0] LLR_383,	input [BIT - 1:0] LLR_384,	input [BIT - 1:0] LLR_385,	input [BIT - 1:0] LLR_386,	input [BIT - 1:0] LLR_387,	input [BIT - 1:0] LLR_388,	input [BIT - 1:0] LLR_389,	input [BIT - 1:0] LLR_390,	input [BIT - 1:0] LLR_391,	input [BIT - 1:0] LLR_392,	input [BIT - 1:0] LLR_393,	input [BIT - 1:0] LLR_394,	input [BIT - 1:0] LLR_395,	input [BIT - 1:0] LLR_396,	input [BIT - 1:0] LLR_397,	input [BIT - 1:0] LLR_398,	input [BIT - 1:0] LLR_399,	input [BIT - 1:0] LLR_400,	input [BIT - 1:0] LLR_401,	input [BIT - 1:0] LLR_402,	input [BIT - 1:0] LLR_403,	input [BIT - 1:0] LLR_404,	input [BIT - 1:0] LLR_405,	input [BIT - 1:0] LLR_406,	input [BIT - 1:0] LLR_407,	input [BIT - 1:0] LLR_408,	input [BIT - 1:0] LLR_409,	input [BIT - 1:0] LLR_410,	input [BIT - 1:0] LLR_411,	input [BIT - 1:0] LLR_412,	input [BIT - 1:0] LLR_413,	input [BIT - 1:0] LLR_414,	input [BIT - 1:0] LLR_415,	input [BIT - 1:0] LLR_416,	input [BIT - 1:0] LLR_417,	input [BIT - 1:0] LLR_418,	input [BIT - 1:0] LLR_419,	input [BIT - 1:0] LLR_420,	input [BIT - 1:0] LLR_421,	input [BIT - 1:0] LLR_422,	input [BIT - 1:0] LLR_423,	input [BIT - 1:0] LLR_424,	input [BIT - 1:0] LLR_425,	input [BIT - 1:0] LLR_426,	input [BIT - 1:0] LLR_427,	input [BIT - 1:0] LLR_428,	input [BIT - 1:0] LLR_429,	input [BIT - 1:0] LLR_430,	input [BIT - 1:0] LLR_431,	input [BIT - 1:0] LLR_432,	input [BIT - 1:0] LLR_433,	input [BIT - 1:0] LLR_434,	input [BIT - 1:0] LLR_435,	input [BIT - 1:0] LLR_436,	input [BIT - 1:0] LLR_437,	input [BIT - 1:0] LLR_438,	input [BIT - 1:0] LLR_439,	input [BIT - 1:0] LLR_440,	input [BIT - 1:0] LLR_441,	input [BIT - 1:0] LLR_442,	input [BIT - 1:0] LLR_443,	input [BIT - 1:0] LLR_444,	input [BIT - 1:0] LLR_445,	input [BIT - 1:0] LLR_446,	input [BIT - 1:0] LLR_447,	input [BIT - 1:0] LLR_448,	input [BIT - 1:0] LLR_449,	input [BIT - 1:0] LLR_450,	input [BIT - 1:0] LLR_451,	input [BIT - 1:0] LLR_452,	input [BIT - 1:0] LLR_453,	input [BIT - 1:0] LLR_454,	input [BIT - 1:0] LLR_455,	input [BIT - 1:0] LLR_456,	input [BIT - 1:0] LLR_457,	input [BIT - 1:0] LLR_458,	input [BIT - 1:0] LLR_459,	input [BIT - 1:0] LLR_460,	input [BIT - 1:0] LLR_461,	input [BIT - 1:0] LLR_462,	input [BIT - 1:0] LLR_463,	input [BIT - 1:0] LLR_464,	input [BIT - 1:0] LLR_465,	input [BIT - 1:0] LLR_466,	input [BIT - 1:0] LLR_467,	input [BIT - 1:0] LLR_468,	input [BIT - 1:0] LLR_469,	input [BIT - 1:0] LLR_470,	input [BIT - 1:0] LLR_471,	input [BIT - 1:0] LLR_472,	input [BIT - 1:0] LLR_473,	input [BIT - 1:0] LLR_474,	input [BIT - 1:0] LLR_475,	input [BIT - 1:0] LLR_476,	input [BIT - 1:0] LLR_477,	input [BIT - 1:0] LLR_478,	input [BIT - 1:0] LLR_479,	input [BIT - 1:0] LLR_480,	input [BIT - 1:0] LLR_481,	input [BIT - 1:0] LLR_482,	input [BIT - 1:0] LLR_483,	input [BIT - 1:0] LLR_484,	input [BIT - 1:0] LLR_485,	input [BIT - 1:0] LLR_486,	input [BIT - 1:0] LLR_487,	input [BIT - 1:0] LLR_488,	input [BIT - 1:0] LLR_489,	input [BIT - 1:0] LLR_490,	input [BIT - 1:0] LLR_491,	input [BIT - 1:0] LLR_492,	input [BIT - 1:0] LLR_493,	input [BIT - 1:0] LLR_494,	input [BIT - 1:0] LLR_495,	input [BIT - 1:0] LLR_496,	input [BIT - 1:0] LLR_497,	input [BIT - 1:0] LLR_498,	input [BIT - 1:0] LLR_499,	input [BIT - 1:0] LLR_500,	input [BIT - 1:0] LLR_501,	input [BIT - 1:0] LLR_502,	input [BIT - 1:0] LLR_503,	input [BIT - 1:0] LLR_504,	input [BIT - 1:0] LLR_505,	input [BIT - 1:0] LLR_506,	input [BIT - 1:0] LLR_507,	input [BIT - 1:0] LLR_508,	input [BIT - 1:0] LLR_509,	input [BIT - 1:0] LLR_510,	input [BIT - 1:0] LLR_511,	input [BIT - 1:0] LLR_512,	input [BIT - 1:0] LLR_513,	input [BIT - 1:0] LLR_514,	input [BIT - 1:0] LLR_515,	input [BIT - 1:0] LLR_516,	input [BIT - 1:0] LLR_517,	input [BIT - 1:0] LLR_518,	input [BIT - 1:0] LLR_519,	input [BIT - 1:0] LLR_520,	input [BIT - 1:0] LLR_521,	input [BIT - 1:0] LLR_522,	input [BIT - 1:0] LLR_523,	input [BIT - 1:0] LLR_524,	input [BIT - 1:0] LLR_525,	input [BIT - 1:0] LLR_526,	input [BIT - 1:0] LLR_527,	input [BIT - 1:0] LLR_528,	input [BIT - 1:0] LLR_529,	input [BIT - 1:0] LLR_530,	input [BIT - 1:0] LLR_531,	input [BIT - 1:0] LLR_532,	input [BIT - 1:0] LLR_533,	input [BIT - 1:0] LLR_534,	input [BIT - 1:0] LLR_535,	input [BIT - 1:0] LLR_536,	input [BIT - 1:0] LLR_537,	input [BIT - 1:0] LLR_538,	input [BIT - 1:0] LLR_539,	input [BIT - 1:0] LLR_540,	input [BIT - 1:0] LLR_541,	input [BIT - 1:0] LLR_542,	input [BIT - 1:0] LLR_543,	input [BIT - 1:0] LLR_544,	input [BIT - 1:0] LLR_545,	input [BIT - 1:0] LLR_546,	input [BIT - 1:0] LLR_547,	input [BIT - 1:0] LLR_548,	input [BIT - 1:0] LLR_549,	input [BIT - 1:0] LLR_550,	input [BIT - 1:0] LLR_551,	input [BIT - 1:0] LLR_552,	input [BIT - 1:0] LLR_553,	input [BIT - 1:0] LLR_554,	input [BIT - 1:0] LLR_555,	input [BIT - 1:0] LLR_556,	input [BIT - 1:0] LLR_557,	input [BIT - 1:0] LLR_558,	input [BIT - 1:0] LLR_559,	input [BIT - 1:0] LLR_560,	input [BIT - 1:0] LLR_561,	input [BIT - 1:0] LLR_562,	input [BIT - 1:0] LLR_563,	input [BIT - 1:0] LLR_564,	input [BIT - 1:0] LLR_565,	input [BIT - 1:0] LLR_566,	input [BIT - 1:0] LLR_567,	input [BIT - 1:0] LLR_568,	input [BIT - 1:0] LLR_569,	input [BIT - 1:0] LLR_570,	input [BIT - 1:0] LLR_571,	input [BIT - 1:0] LLR_572,	input [BIT - 1:0] LLR_573,	input [BIT - 1:0] LLR_574,	input [BIT - 1:0] LLR_575,	input [BIT - 1:0] LLR_576,	input [BIT - 1:0] LLR_577,	input [BIT - 1:0] LLR_578,	input [BIT - 1:0] LLR_579,	input [BIT - 1:0] LLR_580,	input [BIT - 1:0] LLR_581,	input [BIT - 1:0] LLR_582,	input [BIT - 1:0] LLR_583,	input [BIT - 1:0] LLR_584,	input [BIT - 1:0] LLR_585,	input [BIT - 1:0] LLR_586,	input [BIT - 1:0] LLR_587,	input [BIT - 1:0] LLR_588,	input [BIT - 1:0] LLR_589,	input [BIT - 1:0] LLR_590,	input [BIT - 1:0] LLR_591,	input [BIT - 1:0] LLR_592,	input [BIT - 1:0] LLR_593,	input [BIT - 1:0] LLR_594,	input [BIT - 1:0] LLR_595,	input [BIT - 1:0] LLR_596,	input [BIT - 1:0] LLR_597,	input [BIT - 1:0] LLR_598,	input [BIT - 1:0] LLR_599,	input [BIT - 1:0] LLR_600,	input [BIT - 1:0] LLR_601,	input [BIT - 1:0] LLR_602,	input [BIT - 1:0] LLR_603,	input [BIT - 1:0] LLR_604,	input [BIT - 1:0] LLR_605,	input [BIT - 1:0] LLR_606,	input [BIT - 1:0] LLR_607,	input [BIT - 1:0] LLR_608,	input [BIT - 1:0] LLR_609,	input [BIT - 1:0] LLR_610,	input [BIT - 1:0] LLR_611,	input [BIT - 1:0] LLR_612,	input [BIT - 1:0] LLR_613,	input [BIT - 1:0] LLR_614,	input [BIT - 1:0] LLR_615,	input [BIT - 1:0] LLR_616,	input [BIT - 1:0] LLR_617,	input [BIT - 1:0] LLR_618,	input [BIT - 1:0] LLR_619,	input [BIT - 1:0] LLR_620,	input [BIT - 1:0] LLR_621,	input [BIT - 1:0] LLR_622,	input [BIT - 1:0] LLR_623,	input [BIT - 1:0] LLR_624,	input [BIT - 1:0] LLR_625,	input [BIT - 1:0] LLR_626,	input [BIT - 1:0] LLR_627,	input [BIT - 1:0] LLR_628,	input [BIT - 1:0] LLR_629,	input [BIT - 1:0] LLR_630,	input [BIT - 1:0] LLR_631,	input [BIT - 1:0] LLR_632,	input [BIT - 1:0] LLR_633,	input [BIT - 1:0] LLR_634,	input [BIT - 1:0] LLR_635,	input [BIT - 1:0] LLR_636,	input [BIT - 1:0] LLR_637,	input [BIT - 1:0] LLR_638,	input [BIT - 1:0] LLR_639,	input [BIT - 1:0] LLR_640,	input [BIT - 1:0] LLR_641,	input [BIT - 1:0] LLR_642,	input [BIT - 1:0] LLR_643,	input [BIT - 1:0] LLR_644,	input [BIT - 1:0] LLR_645,	input [BIT - 1:0] LLR_646,	input [BIT - 1:0] LLR_647,	input [BIT - 1:0] LLR_648,	input [BIT - 1:0] LLR_649,	input [BIT - 1:0] LLR_650,	input [BIT - 1:0] LLR_651,	input [BIT - 1:0] LLR_652,	input [BIT - 1:0] LLR_653,	input [BIT - 1:0] LLR_654,	input [BIT - 1:0] LLR_655,	input [BIT - 1:0] LLR_656,	input [BIT - 1:0] LLR_657,	input [BIT - 1:0] LLR_658,	input [BIT - 1:0] LLR_659,	input [BIT - 1:0] LLR_660,	input [BIT - 1:0] LLR_661,	input [BIT - 1:0] LLR_662,	input [BIT - 1:0] LLR_663,	input [BIT - 1:0] LLR_664,	input [BIT - 1:0] LLR_665,	input [BIT - 1:0] LLR_666,	input [BIT - 1:0] LLR_667,	input [BIT - 1:0] LLR_668,	input [BIT - 1:0] LLR_669,	input [BIT - 1:0] LLR_670,	input [BIT - 1:0] LLR_671,	input [BIT - 1:0] LLR_672,	input [BIT - 1:0] LLR_673,	input [BIT - 1:0] LLR_674,	input [BIT - 1:0] LLR_675,	input [BIT - 1:0] LLR_676,	input [BIT - 1:0] LLR_677,	input [BIT - 1:0] LLR_678,	input [BIT - 1:0] LLR_679,	input [BIT - 1:0] LLR_680,	input [BIT - 1:0] LLR_681,	input [BIT - 1:0] LLR_682,	input [BIT - 1:0] LLR_683,	input [BIT - 1:0] LLR_684,	input [BIT - 1:0] LLR_685,	input [BIT - 1:0] LLR_686,	input [BIT - 1:0] LLR_687,	input [BIT - 1:0] LLR_688,	input [BIT - 1:0] LLR_689,	input [BIT - 1:0] LLR_690,	input [BIT - 1:0] LLR_691,	input [BIT - 1:0] LLR_692,	input [BIT - 1:0] LLR_693,	input [BIT - 1:0] LLR_694,	input [BIT - 1:0] LLR_695,	input [BIT - 1:0] LLR_696,	input [BIT - 1:0] LLR_697,	input [BIT - 1:0] LLR_698,	input [BIT - 1:0] LLR_699,	input [BIT - 1:0] LLR_700,	input [BIT - 1:0] LLR_701,	input [BIT - 1:0] LLR_702,	input [BIT - 1:0] LLR_703,	input [BIT - 1:0] LLR_704,	input [BIT - 1:0] LLR_705,	input [BIT - 1:0] LLR_706,	input [BIT - 1:0] LLR_707,	input [BIT - 1:0] LLR_708,	input [BIT - 1:0] LLR_709,	input [BIT - 1:0] LLR_710,	input [BIT - 1:0] LLR_711,	input [BIT - 1:0] LLR_712,	input [BIT - 1:0] LLR_713,	input [BIT - 1:0] LLR_714,	input [BIT - 1:0] LLR_715,	input [BIT - 1:0] LLR_716,	input [BIT - 1:0] LLR_717,	input [BIT - 1:0] LLR_718,	input [BIT - 1:0] LLR_719,	input [BIT - 1:0] LLR_720,	input [BIT - 1:0] LLR_721,	input [BIT - 1:0] LLR_722,	input [BIT - 1:0] LLR_723,	input [BIT - 1:0] LLR_724,	input [BIT - 1:0] LLR_725,	input [BIT - 1:0] LLR_726,	input [BIT - 1:0] LLR_727,	input [BIT - 1:0] LLR_728,	input [BIT - 1:0] LLR_729,	input [BIT - 1:0] LLR_730,	input [BIT - 1:0] LLR_731,	input [BIT - 1:0] LLR_732,	input [BIT - 1:0] LLR_733,	input [BIT - 1:0] LLR_734,	input [BIT - 1:0] LLR_735,	input [BIT - 1:0] LLR_736,	input [BIT - 1:0] LLR_737,	input [BIT - 1:0] LLR_738,	input [BIT - 1:0] LLR_739,	input [BIT - 1:0] LLR_740,	input [BIT - 1:0] LLR_741,	input [BIT - 1:0] LLR_742,	input [BIT - 1:0] LLR_743,	input [BIT - 1:0] LLR_744,	input [BIT - 1:0] LLR_745,	input [BIT - 1:0] LLR_746,	input [BIT - 1:0] LLR_747,	input [BIT - 1:0] LLR_748,	input [BIT - 1:0] LLR_749,	input [BIT - 1:0] LLR_750,	input [BIT - 1:0] LLR_751,	input [BIT - 1:0] LLR_752,	input [BIT - 1:0] LLR_753,	input [BIT - 1:0] LLR_754,	input [BIT - 1:0] LLR_755,	input [BIT - 1:0] LLR_756,	input [BIT - 1:0] LLR_757,	input [BIT - 1:0] LLR_758,	input [BIT - 1:0] LLR_759,	input [BIT - 1:0] LLR_760,	input [BIT - 1:0] LLR_761,	input [BIT - 1:0] LLR_762,	input [BIT - 1:0] LLR_763,	input [BIT - 1:0] LLR_764,	input [BIT - 1:0] LLR_765,	input [BIT - 1:0] LLR_766,	input [BIT - 1:0] LLR_767,	input [BIT - 1:0] LLR_768,	input [BIT - 1:0] LLR_769,	input [BIT - 1:0] LLR_770,	input [BIT - 1:0] LLR_771,	input [BIT - 1:0] LLR_772,	input [BIT - 1:0] LLR_773,	input [BIT - 1:0] LLR_774,	input [BIT - 1:0] LLR_775,	input [BIT - 1:0] LLR_776,	input [BIT - 1:0] LLR_777,	input [BIT - 1:0] LLR_778,	input [BIT - 1:0] LLR_779,	input [BIT - 1:0] LLR_780,	input [BIT - 1:0] LLR_781,	input [BIT - 1:0] LLR_782,	input [BIT - 1:0] LLR_783,	input [BIT - 1:0] LLR_784,	input [BIT - 1:0] LLR_785,	input [BIT - 1:0] LLR_786,	input [BIT - 1:0] LLR_787,	input [BIT - 1:0] LLR_788,	input [BIT - 1:0] LLR_789,	input [BIT - 1:0] LLR_790,	input [BIT - 1:0] LLR_791,	input [BIT - 1:0] LLR_792,	input [BIT - 1:0] LLR_793,	input [BIT - 1:0] LLR_794,	input [BIT - 1:0] LLR_795,	input [BIT - 1:0] LLR_796,	input [BIT - 1:0] LLR_797,	input [BIT - 1:0] LLR_798,	input [BIT - 1:0] LLR_799,	input [BIT - 1:0] LLR_800,	input [BIT - 1:0] LLR_801,	input [BIT - 1:0] LLR_802,	input [BIT - 1:0] LLR_803,	input [BIT - 1:0] LLR_804,	input [BIT - 1:0] LLR_805,	input [BIT - 1:0] LLR_806,	input [BIT - 1:0] LLR_807,	input [BIT - 1:0] LLR_808,	input [BIT - 1:0] LLR_809,	input [BIT - 1:0] LLR_810,	input [BIT - 1:0] LLR_811,	input [BIT - 1:0] LLR_812,	input [BIT - 1:0] LLR_813,	input [BIT - 1:0] LLR_814,	input [BIT - 1:0] LLR_815,	input [BIT - 1:0] LLR_816,	input [BIT - 1:0] LLR_817,	input [BIT - 1:0] LLR_818,	input [BIT - 1:0] LLR_819,	input [BIT - 1:0] LLR_820,	input [BIT - 1:0] LLR_821,	input [BIT - 1:0] LLR_822,	input [BIT - 1:0] LLR_823,	input [BIT - 1:0] LLR_824,	input [BIT - 1:0] LLR_825,	input [BIT - 1:0] LLR_826,	input [BIT - 1:0] LLR_827,	input [BIT - 1:0] LLR_828,	input [BIT - 1:0] LLR_829,	input [BIT - 1:0] LLR_830,	input [BIT - 1:0] LLR_831,	input [BIT - 1:0] LLR_832,	input [BIT - 1:0] LLR_833,	input [BIT - 1:0] LLR_834,	input [BIT - 1:0] LLR_835,	input [BIT - 1:0] LLR_836,	input [BIT - 1:0] LLR_837,	input [BIT - 1:0] LLR_838,	input [BIT - 1:0] LLR_839,	input [BIT - 1:0] LLR_840,	input [BIT - 1:0] LLR_841,	input [BIT - 1:0] LLR_842,	input [BIT - 1:0] LLR_843,	input [BIT - 1:0] LLR_844,	input [BIT - 1:0] LLR_845,	input [BIT - 1:0] LLR_846,	input [BIT - 1:0] LLR_847,	input [BIT - 1:0] LLR_848,	input [BIT - 1:0] LLR_849,	input [BIT - 1:0] LLR_850,	input [BIT - 1:0] LLR_851,	input [BIT - 1:0] LLR_852,	input [BIT - 1:0] LLR_853,	input [BIT - 1:0] LLR_854,	input [BIT - 1:0] LLR_855,	input [BIT - 1:0] LLR_856,	input [BIT - 1:0] LLR_857,	input [BIT - 1:0] LLR_858,	input [BIT - 1:0] LLR_859,	input [BIT - 1:0] LLR_860,	input [BIT - 1:0] LLR_861,	input [BIT - 1:0] LLR_862,	input [BIT - 1:0] LLR_863,	input [BIT - 1:0] LLR_864,	input [BIT - 1:0] LLR_865,	input [BIT - 1:0] LLR_866,	input [BIT - 1:0] LLR_867,	input [BIT - 1:0] LLR_868,	input [BIT - 1:0] LLR_869,	input [BIT - 1:0] LLR_870,	input [BIT - 1:0] LLR_871,	input [BIT - 1:0] LLR_872,	input [BIT - 1:0] LLR_873,	input [BIT - 1:0] LLR_874,	input [BIT - 1:0] LLR_875,	input [BIT - 1:0] LLR_876,	input [BIT - 1:0] LLR_877,	input [BIT - 1:0] LLR_878,	input [BIT - 1:0] LLR_879,	input [BIT - 1:0] LLR_880,	input [BIT - 1:0] LLR_881,	input [BIT - 1:0] LLR_882,	input [BIT - 1:0] LLR_883,	input [BIT - 1:0] LLR_884,	input [BIT - 1:0] LLR_885,	input [BIT - 1:0] LLR_886,	input [BIT - 1:0] LLR_887,	input [BIT - 1:0] LLR_888,	input [BIT - 1:0] LLR_889,	input [BIT - 1:0] LLR_890,	input [BIT - 1:0] LLR_891,	input [BIT - 1:0] LLR_892,	input [BIT - 1:0] LLR_893,	input [BIT - 1:0] LLR_894,	input [BIT - 1:0] LLR_895,	input [BIT - 1:0] LLR_896,	input [BIT - 1:0] LLR_897,	input [BIT - 1:0] LLR_898,	input [BIT - 1:0] LLR_899,	input [BIT - 1:0] LLR_900,	input [BIT - 1:0] LLR_901,	input [BIT - 1:0] LLR_902,	input [BIT - 1:0] LLR_903,	input [BIT - 1:0] LLR_904,	input [BIT - 1:0] LLR_905,	input [BIT - 1:0] LLR_906,	input [BIT - 1:0] LLR_907,	input [BIT - 1:0] LLR_908,	input [BIT - 1:0] LLR_909,	input [BIT - 1:0] LLR_910,	input [BIT - 1:0] LLR_911,	input [BIT - 1:0] LLR_912,	input [BIT - 1:0] LLR_913,	input [BIT - 1:0] LLR_914,	input [BIT - 1:0] LLR_915,	input [BIT - 1:0] LLR_916,	input [BIT - 1:0] LLR_917,	input [BIT - 1:0] LLR_918,	input [BIT - 1:0] LLR_919,	input [BIT - 1:0] LLR_920,	input [BIT - 1:0] LLR_921,	input [BIT - 1:0] LLR_922,	input [BIT - 1:0] LLR_923,	input [BIT - 1:0] LLR_924,	input [BIT - 1:0] LLR_925,	input [BIT - 1:0] LLR_926,	input [BIT - 1:0] LLR_927,	input [BIT - 1:0] LLR_928,	input [BIT - 1:0] LLR_929,	input [BIT - 1:0] LLR_930,	input [BIT - 1:0] LLR_931,	input [BIT - 1:0] LLR_932,	input [BIT - 1:0] LLR_933,	input [BIT - 1:0] LLR_934,	input [BIT - 1:0] LLR_935,	input [BIT - 1:0] LLR_936,	input [BIT - 1:0] LLR_937,	input [BIT - 1:0] LLR_938,	input [BIT - 1:0] LLR_939,	input [BIT - 1:0] LLR_940,	input [BIT - 1:0] LLR_941,	input [BIT - 1:0] LLR_942,	input [BIT - 1:0] LLR_943,	input [BIT - 1:0] LLR_944,	input [BIT - 1:0] LLR_945,	input [BIT - 1:0] LLR_946,	input [BIT - 1:0] LLR_947,	input [BIT - 1:0] LLR_948,	input [BIT - 1:0] LLR_949,	input [BIT - 1:0] LLR_950,	input [BIT - 1:0] LLR_951,	input [BIT - 1:0] LLR_952,	input [BIT - 1:0] LLR_953,	input [BIT - 1:0] LLR_954,	input [BIT - 1:0] LLR_955,	input [BIT - 1:0] LLR_956,	input [BIT - 1:0] LLR_957,	input [BIT - 1:0] LLR_958,	input [BIT - 1:0] LLR_959,	input [BIT - 1:0] LLR_960,	input [BIT - 1:0] LLR_961,	input [BIT - 1:0] LLR_962,	input [BIT - 1:0] LLR_963,	input [BIT - 1:0] LLR_964,	input [BIT - 1:0] LLR_965,	input [BIT - 1:0] LLR_966,	input [BIT - 1:0] LLR_967,	input [BIT - 1:0] LLR_968,	input [BIT - 1:0] LLR_969,	input [BIT - 1:0] LLR_970,	input [BIT - 1:0] LLR_971,	input [BIT - 1:0] LLR_972,	input [BIT - 1:0] LLR_973,	input [BIT - 1:0] LLR_974,	input [BIT - 1:0] LLR_975,	input [BIT - 1:0] LLR_976,	input [BIT - 1:0] LLR_977,	input [BIT - 1:0] LLR_978,	input [BIT - 1:0] LLR_979,	input [BIT - 1:0] LLR_980,	input [BIT - 1:0] LLR_981,	input [BIT - 1:0] LLR_982,	input [BIT - 1:0] LLR_983,	input [BIT - 1:0] LLR_984,	input [BIT - 1:0] LLR_985,	input [BIT - 1:0] LLR_986,	input [BIT - 1:0] LLR_987,	input [BIT - 1:0] LLR_988,	input [BIT - 1:0] LLR_989,	input [BIT - 1:0] LLR_990,	input [BIT - 1:0] LLR_991,	input [BIT - 1:0] LLR_992,	input [BIT - 1:0] LLR_993,	input [BIT - 1:0] LLR_994,	input [BIT - 1:0] LLR_995,	input [BIT - 1:0] LLR_996,	input [BIT - 1:0] LLR_997,	input [BIT - 1:0] LLR_998,	input [BIT - 1:0] LLR_999,	input [BIT - 1:0] LLR_1000,	input [BIT - 1:0] LLR_1001,	input [BIT - 1:0] LLR_1002,	input [BIT - 1:0] LLR_1003,	input [BIT - 1:0] LLR_1004,	input [BIT - 1:0] LLR_1005,	input [BIT - 1:0] LLR_1006,	input [BIT - 1:0] LLR_1007,	input [BIT - 1:0] LLR_1008,	input [BIT - 1:0] LLR_1009,	input [BIT - 1:0] LLR_1010,	input [BIT - 1:0] LLR_1011,	input [BIT - 1:0] LLR_1012,	input [BIT - 1:0] LLR_1013,	input [BIT - 1:0] LLR_1014,	input [BIT - 1:0] LLR_1015,	input [BIT - 1:0] LLR_1016,	input [BIT - 1:0] LLR_1017,	input [BIT - 1:0] LLR_1018,	input [BIT - 1:0] LLR_1019,	input [BIT - 1:0] LLR_1020,	input [BIT - 1:0] LLR_1021,	input [BIT - 1:0] LLR_1022,	input [BIT - 1:0] LLR_1023,	input [BIT - 1:0] LLR_1024,	output reg [BIT - 1:0] OUT_1,	output reg [BIT - 1:0] OUT_2,	output reg [BIT - 1:0] OUT_3,	output reg [BIT - 1:0] OUT_4,	output reg [BIT - 1:0] OUT_5,	output reg [BIT - 1:0] OUT_6,	output reg [BIT - 1:0] OUT_7,	output reg [BIT - 1:0] OUT_8,	output reg [BIT - 1:0] OUT_9,	output reg [BIT - 1:0] OUT_10,	output reg [BIT - 1:0] OUT_11,	output reg [BIT - 1:0] OUT_12,	output reg [BIT - 1:0] OUT_13,	output reg [BIT - 1:0] OUT_14,	output reg [BIT - 1:0] OUT_15,	output reg [BIT - 1:0] OUT_16,	output reg [BIT - 1:0] OUT_17,	output reg [BIT - 1:0] OUT_18,	output reg [BIT - 1:0] OUT_19,	output reg [BIT - 1:0] OUT_20,	output reg [BIT - 1:0] OUT_21,	output reg [BIT - 1:0] OUT_22,	output reg [BIT - 1:0] OUT_23,	output reg [BIT - 1:0] OUT_24,	output reg [BIT - 1:0] OUT_25,	output reg [BIT - 1:0] OUT_26,	output reg [BIT - 1:0] OUT_27,	output reg [BIT - 1:0] OUT_28,	output reg [BIT - 1:0] OUT_29,	output reg [BIT - 1:0] OUT_30,	output reg [BIT - 1:0] OUT_31,	output reg [BIT - 1:0] OUT_32,	output reg [BIT - 1:0] OUT_33,	output reg [BIT - 1:0] OUT_34,	output reg [BIT - 1:0] OUT_35,	output reg [BIT - 1:0] OUT_36,	output reg [BIT - 1:0] OUT_37,	output reg [BIT - 1:0] OUT_38,	output reg [BIT - 1:0] OUT_39,	output reg [BIT - 1:0] OUT_40,	output reg [BIT - 1:0] OUT_41,	output reg [BIT - 1:0] OUT_42,	output reg [BIT - 1:0] OUT_43,	output reg [BIT - 1:0] OUT_44,	output reg [BIT - 1:0] OUT_45,	output reg [BIT - 1:0] OUT_46,	output reg [BIT - 1:0] OUT_47,	output reg [BIT - 1:0] OUT_48,	output reg [BIT - 1:0] OUT_49,	output reg [BIT - 1:0] OUT_50,	output reg [BIT - 1:0] OUT_51,	output reg [BIT - 1:0] OUT_52,	output reg [BIT - 1:0] OUT_53,	output reg [BIT - 1:0] OUT_54,	output reg [BIT - 1:0] OUT_55,	output reg [BIT - 1:0] OUT_56,	output reg [BIT - 1:0] OUT_57,	output reg [BIT - 1:0] OUT_58,	output reg [BIT - 1:0] OUT_59,	output reg [BIT - 1:0] OUT_60,	output reg [BIT - 1:0] OUT_61,	output reg [BIT - 1:0] OUT_62,	output reg [BIT - 1:0] OUT_63,	output reg [BIT - 1:0] OUT_64,	output reg [BIT - 1:0] OUT_65,	output reg [BIT - 1:0] OUT_66,	output reg [BIT - 1:0] OUT_67,	output reg [BIT - 1:0] OUT_68,	output reg [BIT - 1:0] OUT_69,	output reg [BIT - 1:0] OUT_70,	output reg [BIT - 1:0] OUT_71,	output reg [BIT - 1:0] OUT_72,	output reg [BIT - 1:0] OUT_73,	output reg [BIT - 1:0] OUT_74,	output reg [BIT - 1:0] OUT_75,	output reg [BIT - 1:0] OUT_76,	output reg [BIT - 1:0] OUT_77,	output reg [BIT - 1:0] OUT_78,	output reg [BIT - 1:0] OUT_79,	output reg [BIT - 1:0] OUT_80,	output reg [BIT - 1:0] OUT_81,	output reg [BIT - 1:0] OUT_82,	output reg [BIT - 1:0] OUT_83,	output reg [BIT - 1:0] OUT_84,	output reg [BIT - 1:0] OUT_85,	output reg [BIT - 1:0] OUT_86,	output reg [BIT - 1:0] OUT_87,	output reg [BIT - 1:0] OUT_88,	output reg [BIT - 1:0] OUT_89,	output reg [BIT - 1:0] OUT_90,	output reg [BIT - 1:0] OUT_91,	output reg [BIT - 1:0] OUT_92,	output reg [BIT - 1:0] OUT_93,	output reg [BIT - 1:0] OUT_94,	output reg [BIT - 1:0] OUT_95,	output reg [BIT - 1:0] OUT_96,	output reg [BIT - 1:0] OUT_97,	output reg [BIT - 1:0] OUT_98,	output reg [BIT - 1:0] OUT_99,	output reg [BIT - 1:0] OUT_100,	output reg [BIT - 1:0] OUT_101,	output reg [BIT - 1:0] OUT_102,	output reg [BIT - 1:0] OUT_103,	output reg [BIT - 1:0] OUT_104,	output reg [BIT - 1:0] OUT_105,	output reg [BIT - 1:0] OUT_106,	output reg [BIT - 1:0] OUT_107,	output reg [BIT - 1:0] OUT_108,	output reg [BIT - 1:0] OUT_109,	output reg [BIT - 1:0] OUT_110,	output reg [BIT - 1:0] OUT_111,	output reg [BIT - 1:0] OUT_112,	output reg [BIT - 1:0] OUT_113,	output reg [BIT - 1:0] OUT_114,	output reg [BIT - 1:0] OUT_115,	output reg [BIT - 1:0] OUT_116,	output reg [BIT - 1:0] OUT_117,	output reg [BIT - 1:0] OUT_118,	output reg [BIT - 1:0] OUT_119,	output reg [BIT - 1:0] OUT_120,	output reg [BIT - 1:0] OUT_121,	output reg [BIT - 1:0] OUT_122,	output reg [BIT - 1:0] OUT_123,	output reg [BIT - 1:0] OUT_124,	output reg [BIT - 1:0] OUT_125,	output reg [BIT - 1:0] OUT_126,	output reg [BIT - 1:0] OUT_127,	output reg [BIT - 1:0] OUT_128,	output reg [BIT - 1:0] OUT_129,	output reg [BIT - 1:0] OUT_130,	output reg [BIT - 1:0] OUT_131,	output reg [BIT - 1:0] OUT_132,	output reg [BIT - 1:0] OUT_133,	output reg [BIT - 1:0] OUT_134,	output reg [BIT - 1:0] OUT_135,	output reg [BIT - 1:0] OUT_136,	output reg [BIT - 1:0] OUT_137,	output reg [BIT - 1:0] OUT_138,	output reg [BIT - 1:0] OUT_139,	output reg [BIT - 1:0] OUT_140,	output reg [BIT - 1:0] OUT_141,	output reg [BIT - 1:0] OUT_142,	output reg [BIT - 1:0] OUT_143,	output reg [BIT - 1:0] OUT_144,	output reg [BIT - 1:0] OUT_145,	output reg [BIT - 1:0] OUT_146,	output reg [BIT - 1:0] OUT_147,	output reg [BIT - 1:0] OUT_148,	output reg [BIT - 1:0] OUT_149,	output reg [BIT - 1:0] OUT_150,	output reg [BIT - 1:0] OUT_151,	output reg [BIT - 1:0] OUT_152,	output reg [BIT - 1:0] OUT_153,	output reg [BIT - 1:0] OUT_154,	output reg [BIT - 1:0] OUT_155,	output reg [BIT - 1:0] OUT_156,	output reg [BIT - 1:0] OUT_157,	output reg [BIT - 1:0] OUT_158,	output reg [BIT - 1:0] OUT_159,	output reg [BIT - 1:0] OUT_160,	output reg [BIT - 1:0] OUT_161,	output reg [BIT - 1:0] OUT_162,	output reg [BIT - 1:0] OUT_163,	output reg [BIT - 1:0] OUT_164,	output reg [BIT - 1:0] OUT_165,	output reg [BIT - 1:0] OUT_166,	output reg [BIT - 1:0] OUT_167,	output reg [BIT - 1:0] OUT_168,	output reg [BIT - 1:0] OUT_169,	output reg [BIT - 1:0] OUT_170,	output reg [BIT - 1:0] OUT_171,	output reg [BIT - 1:0] OUT_172,	output reg [BIT - 1:0] OUT_173,	output reg [BIT - 1:0] OUT_174,	output reg [BIT - 1:0] OUT_175,	output reg [BIT - 1:0] OUT_176,	output reg [BIT - 1:0] OUT_177,	output reg [BIT - 1:0] OUT_178,	output reg [BIT - 1:0] OUT_179,	output reg [BIT - 1:0] OUT_180,	output reg [BIT - 1:0] OUT_181,	output reg [BIT - 1:0] OUT_182,	output reg [BIT - 1:0] OUT_183,	output reg [BIT - 1:0] OUT_184,	output reg [BIT - 1:0] OUT_185,	output reg [BIT - 1:0] OUT_186,	output reg [BIT - 1:0] OUT_187,	output reg [BIT - 1:0] OUT_188,	output reg [BIT - 1:0] OUT_189,	output reg [BIT - 1:0] OUT_190,	output reg [BIT - 1:0] OUT_191,	output reg [BIT - 1:0] OUT_192,	output reg [BIT - 1:0] OUT_193,	output reg [BIT - 1:0] OUT_194,	output reg [BIT - 1:0] OUT_195,	output reg [BIT - 1:0] OUT_196,	output reg [BIT - 1:0] OUT_197,	output reg [BIT - 1:0] OUT_198,	output reg [BIT - 1:0] OUT_199,	output reg [BIT - 1:0] OUT_200,	output reg [BIT - 1:0] OUT_201,	output reg [BIT - 1:0] OUT_202,	output reg [BIT - 1:0] OUT_203,	output reg [BIT - 1:0] OUT_204,	output reg [BIT - 1:0] OUT_205,	output reg [BIT - 1:0] OUT_206,	output reg [BIT - 1:0] OUT_207,	output reg [BIT - 1:0] OUT_208,	output reg [BIT - 1:0] OUT_209,	output reg [BIT - 1:0] OUT_210,	output reg [BIT - 1:0] OUT_211,	output reg [BIT - 1:0] OUT_212,	output reg [BIT - 1:0] OUT_213,	output reg [BIT - 1:0] OUT_214,	output reg [BIT - 1:0] OUT_215,	output reg [BIT - 1:0] OUT_216,	output reg [BIT - 1:0] OUT_217,	output reg [BIT - 1:0] OUT_218,	output reg [BIT - 1:0] OUT_219,	output reg [BIT - 1:0] OUT_220,	output reg [BIT - 1:0] OUT_221,	output reg [BIT - 1:0] OUT_222,	output reg [BIT - 1:0] OUT_223,	output reg [BIT - 1:0] OUT_224,	output reg [BIT - 1:0] OUT_225,	output reg [BIT - 1:0] OUT_226,	output reg [BIT - 1:0] OUT_227,	output reg [BIT - 1:0] OUT_228,	output reg [BIT - 1:0] OUT_229,	output reg [BIT - 1:0] OUT_230,	output reg [BIT - 1:0] OUT_231,	output reg [BIT - 1:0] OUT_232,	output reg [BIT - 1:0] OUT_233,	output reg [BIT - 1:0] OUT_234,	output reg [BIT - 1:0] OUT_235,	output reg [BIT - 1:0] OUT_236,	output reg [BIT - 1:0] OUT_237,	output reg [BIT - 1:0] OUT_238,	output reg [BIT - 1:0] OUT_239,	output reg [BIT - 1:0] OUT_240,	output reg [BIT - 1:0] OUT_241,	output reg [BIT - 1:0] OUT_242,	output reg [BIT - 1:0] OUT_243,	output reg [BIT - 1:0] OUT_244,	output reg [BIT - 1:0] OUT_245,	output reg [BIT - 1:0] OUT_246,	output reg [BIT - 1:0] OUT_247,	output reg [BIT - 1:0] OUT_248,	output reg [BIT - 1:0] OUT_249,	output reg [BIT - 1:0] OUT_250,	output reg [BIT - 1:0] OUT_251,	output reg [BIT - 1:0] OUT_252,	output reg [BIT - 1:0] OUT_253,	output reg [BIT - 1:0] OUT_254,	output reg [BIT - 1:0] OUT_255,	output reg [BIT - 1:0] OUT_256,	output reg [BIT - 1:0] OUT_257,	output reg [BIT - 1:0] OUT_258,	output reg [BIT - 1:0] OUT_259,	output reg [BIT - 1:0] OUT_260,	output reg [BIT - 1:0] OUT_261,	output reg [BIT - 1:0] OUT_262,	output reg [BIT - 1:0] OUT_263,	output reg [BIT - 1:0] OUT_264,	output reg [BIT - 1:0] OUT_265,	output reg [BIT - 1:0] OUT_266,	output reg [BIT - 1:0] OUT_267,	output reg [BIT - 1:0] OUT_268,	output reg [BIT - 1:0] OUT_269,	output reg [BIT - 1:0] OUT_270,	output reg [BIT - 1:0] OUT_271,	output reg [BIT - 1:0] OUT_272,	output reg [BIT - 1:0] OUT_273,	output reg [BIT - 1:0] OUT_274,	output reg [BIT - 1:0] OUT_275,	output reg [BIT - 1:0] OUT_276,	output reg [BIT - 1:0] OUT_277,	output reg [BIT - 1:0] OUT_278,	output reg [BIT - 1:0] OUT_279,	output reg [BIT - 1:0] OUT_280,	output reg [BIT - 1:0] OUT_281,	output reg [BIT - 1:0] OUT_282,	output reg [BIT - 1:0] OUT_283,	output reg [BIT - 1:0] OUT_284,	output reg [BIT - 1:0] OUT_285,	output reg [BIT - 1:0] OUT_286,	output reg [BIT - 1:0] OUT_287,	output reg [BIT - 1:0] OUT_288,	output reg [BIT - 1:0] OUT_289,	output reg [BIT - 1:0] OUT_290,	output reg [BIT - 1:0] OUT_291,	output reg [BIT - 1:0] OUT_292,	output reg [BIT - 1:0] OUT_293,	output reg [BIT - 1:0] OUT_294,	output reg [BIT - 1:0] OUT_295,	output reg [BIT - 1:0] OUT_296,	output reg [BIT - 1:0] OUT_297,	output reg [BIT - 1:0] OUT_298,	output reg [BIT - 1:0] OUT_299,	output reg [BIT - 1:0] OUT_300,	output reg [BIT - 1:0] OUT_301,	output reg [BIT - 1:0] OUT_302,	output reg [BIT - 1:0] OUT_303,	output reg [BIT - 1:0] OUT_304,	output reg [BIT - 1:0] OUT_305,	output reg [BIT - 1:0] OUT_306,	output reg [BIT - 1:0] OUT_307,	output reg [BIT - 1:0] OUT_308,	output reg [BIT - 1:0] OUT_309,	output reg [BIT - 1:0] OUT_310,	output reg [BIT - 1:0] OUT_311,	output reg [BIT - 1:0] OUT_312,	output reg [BIT - 1:0] OUT_313,	output reg [BIT - 1:0] OUT_314,	output reg [BIT - 1:0] OUT_315,	output reg [BIT - 1:0] OUT_316,	output reg [BIT - 1:0] OUT_317,	output reg [BIT - 1:0] OUT_318,	output reg [BIT - 1:0] OUT_319,	output reg [BIT - 1:0] OUT_320,	output reg [BIT - 1:0] OUT_321,	output reg [BIT - 1:0] OUT_322,	output reg [BIT - 1:0] OUT_323,	output reg [BIT - 1:0] OUT_324,	output reg [BIT - 1:0] OUT_325,	output reg [BIT - 1:0] OUT_326,	output reg [BIT - 1:0] OUT_327,	output reg [BIT - 1:0] OUT_328,	output reg [BIT - 1:0] OUT_329,	output reg [BIT - 1:0] OUT_330,	output reg [BIT - 1:0] OUT_331,	output reg [BIT - 1:0] OUT_332,	output reg [BIT - 1:0] OUT_333,	output reg [BIT - 1:0] OUT_334,	output reg [BIT - 1:0] OUT_335,	output reg [BIT - 1:0] OUT_336,	output reg [BIT - 1:0] OUT_337,	output reg [BIT - 1:0] OUT_338,	output reg [BIT - 1:0] OUT_339,	output reg [BIT - 1:0] OUT_340,	output reg [BIT - 1:0] OUT_341,	output reg [BIT - 1:0] OUT_342,	output reg [BIT - 1:0] OUT_343,	output reg [BIT - 1:0] OUT_344,	output reg [BIT - 1:0] OUT_345,	output reg [BIT - 1:0] OUT_346,	output reg [BIT - 1:0] OUT_347,	output reg [BIT - 1:0] OUT_348,	output reg [BIT - 1:0] OUT_349,	output reg [BIT - 1:0] OUT_350,	output reg [BIT - 1:0] OUT_351,	output reg [BIT - 1:0] OUT_352,	output reg [BIT - 1:0] OUT_353,	output reg [BIT - 1:0] OUT_354,	output reg [BIT - 1:0] OUT_355,	output reg [BIT - 1:0] OUT_356,	output reg [BIT - 1:0] OUT_357,	output reg [BIT - 1:0] OUT_358,	output reg [BIT - 1:0] OUT_359,	output reg [BIT - 1:0] OUT_360,	output reg [BIT - 1:0] OUT_361,	output reg [BIT - 1:0] OUT_362,	output reg [BIT - 1:0] OUT_363,	output reg [BIT - 1:0] OUT_364,	output reg [BIT - 1:0] OUT_365,	output reg [BIT - 1:0] OUT_366,	output reg [BIT - 1:0] OUT_367,	output reg [BIT - 1:0] OUT_368,	output reg [BIT - 1:0] OUT_369,	output reg [BIT - 1:0] OUT_370,	output reg [BIT - 1:0] OUT_371,	output reg [BIT - 1:0] OUT_372,	output reg [BIT - 1:0] OUT_373,	output reg [BIT - 1:0] OUT_374,	output reg [BIT - 1:0] OUT_375,	output reg [BIT - 1:0] OUT_376,	output reg [BIT - 1:0] OUT_377,	output reg [BIT - 1:0] OUT_378,	output reg [BIT - 1:0] OUT_379,	output reg [BIT - 1:0] OUT_380,	output reg [BIT - 1:0] OUT_381,	output reg [BIT - 1:0] OUT_382,	output reg [BIT - 1:0] OUT_383,	output reg [BIT - 1:0] OUT_384,	output reg [BIT - 1:0] OUT_385,	output reg [BIT - 1:0] OUT_386,	output reg [BIT - 1:0] OUT_387,	output reg [BIT - 1:0] OUT_388,	output reg [BIT - 1:0] OUT_389,	output reg [BIT - 1:0] OUT_390,	output reg [BIT - 1:0] OUT_391,	output reg [BIT - 1:0] OUT_392,	output reg [BIT - 1:0] OUT_393,	output reg [BIT - 1:0] OUT_394,	output reg [BIT - 1:0] OUT_395,	output reg [BIT - 1:0] OUT_396,	output reg [BIT - 1:0] OUT_397,	output reg [BIT - 1:0] OUT_398,	output reg [BIT - 1:0] OUT_399,	output reg [BIT - 1:0] OUT_400,	output reg [BIT - 1:0] OUT_401,	output reg [BIT - 1:0] OUT_402,	output reg [BIT - 1:0] OUT_403,	output reg [BIT - 1:0] OUT_404,	output reg [BIT - 1:0] OUT_405,	output reg [BIT - 1:0] OUT_406,	output reg [BIT - 1:0] OUT_407,	output reg [BIT - 1:0] OUT_408,	output reg [BIT - 1:0] OUT_409,	output reg [BIT - 1:0] OUT_410,	output reg [BIT - 1:0] OUT_411,	output reg [BIT - 1:0] OUT_412,	output reg [BIT - 1:0] OUT_413,	output reg [BIT - 1:0] OUT_414,	output reg [BIT - 1:0] OUT_415,	output reg [BIT - 1:0] OUT_416,	output reg [BIT - 1:0] OUT_417,	output reg [BIT - 1:0] OUT_418,	output reg [BIT - 1:0] OUT_419,	output reg [BIT - 1:0] OUT_420,	output reg [BIT - 1:0] OUT_421,	output reg [BIT - 1:0] OUT_422,	output reg [BIT - 1:0] OUT_423,	output reg [BIT - 1:0] OUT_424,	output reg [BIT - 1:0] OUT_425,	output reg [BIT - 1:0] OUT_426,	output reg [BIT - 1:0] OUT_427,	output reg [BIT - 1:0] OUT_428,	output reg [BIT - 1:0] OUT_429,	output reg [BIT - 1:0] OUT_430,	output reg [BIT - 1:0] OUT_431,	output reg [BIT - 1:0] OUT_432,	output reg [BIT - 1:0] OUT_433,	output reg [BIT - 1:0] OUT_434,	output reg [BIT - 1:0] OUT_435,	output reg [BIT - 1:0] OUT_436,	output reg [BIT - 1:0] OUT_437,	output reg [BIT - 1:0] OUT_438,	output reg [BIT - 1:0] OUT_439,	output reg [BIT - 1:0] OUT_440,	output reg [BIT - 1:0] OUT_441,	output reg [BIT - 1:0] OUT_442,	output reg [BIT - 1:0] OUT_443,	output reg [BIT - 1:0] OUT_444,	output reg [BIT - 1:0] OUT_445,	output reg [BIT - 1:0] OUT_446,	output reg [BIT - 1:0] OUT_447,	output reg [BIT - 1:0] OUT_448,	output reg [BIT - 1:0] OUT_449,	output reg [BIT - 1:0] OUT_450,	output reg [BIT - 1:0] OUT_451,	output reg [BIT - 1:0] OUT_452,	output reg [BIT - 1:0] OUT_453,	output reg [BIT - 1:0] OUT_454,	output reg [BIT - 1:0] OUT_455,	output reg [BIT - 1:0] OUT_456,	output reg [BIT - 1:0] OUT_457,	output reg [BIT - 1:0] OUT_458,	output reg [BIT - 1:0] OUT_459,	output reg [BIT - 1:0] OUT_460,	output reg [BIT - 1:0] OUT_461,	output reg [BIT - 1:0] OUT_462,	output reg [BIT - 1:0] OUT_463,	output reg [BIT - 1:0] OUT_464,	output reg [BIT - 1:0] OUT_465,	output reg [BIT - 1:0] OUT_466,	output reg [BIT - 1:0] OUT_467,	output reg [BIT - 1:0] OUT_468,	output reg [BIT - 1:0] OUT_469,	output reg [BIT - 1:0] OUT_470,	output reg [BIT - 1:0] OUT_471,	output reg [BIT - 1:0] OUT_472,	output reg [BIT - 1:0] OUT_473,	output reg [BIT - 1:0] OUT_474,	output reg [BIT - 1:0] OUT_475,	output reg [BIT - 1:0] OUT_476,	output reg [BIT - 1:0] OUT_477,	output reg [BIT - 1:0] OUT_478,	output reg [BIT - 1:0] OUT_479,	output reg [BIT - 1:0] OUT_480,	output reg [BIT - 1:0] OUT_481,	output reg [BIT - 1:0] OUT_482,	output reg [BIT - 1:0] OUT_483,	output reg [BIT - 1:0] OUT_484,	output reg [BIT - 1:0] OUT_485,	output reg [BIT - 1:0] OUT_486,	output reg [BIT - 1:0] OUT_487,	output reg [BIT - 1:0] OUT_488,	output reg [BIT - 1:0] OUT_489,	output reg [BIT - 1:0] OUT_490,	output reg [BIT - 1:0] OUT_491,	output reg [BIT - 1:0] OUT_492,	output reg [BIT - 1:0] OUT_493,	output reg [BIT - 1:0] OUT_494,	output reg [BIT - 1:0] OUT_495,	output reg [BIT - 1:0] OUT_496,	output reg [BIT - 1:0] OUT_497,	output reg [BIT - 1:0] OUT_498,	output reg [BIT - 1:0] OUT_499,	output reg [BIT - 1:0] OUT_500,	output reg [BIT - 1:0] OUT_501,	output reg [BIT - 1:0] OUT_502,	output reg [BIT - 1:0] OUT_503,	output reg [BIT - 1:0] OUT_504,	output reg [BIT - 1:0] OUT_505,	output reg [BIT - 1:0] OUT_506,	output reg [BIT - 1:0] OUT_507,	output reg [BIT - 1:0] OUT_508,	output reg [BIT - 1:0] OUT_509,	output reg [BIT - 1:0] OUT_510,	output reg [BIT - 1:0] OUT_511,	output reg [BIT - 1:0] OUT_512,	output reg [BIT - 1:0] OUT_513,	output reg [BIT - 1:0] OUT_514,	output reg [BIT - 1:0] OUT_515,	output reg [BIT - 1:0] OUT_516,	output reg [BIT - 1:0] OUT_517,	output reg [BIT - 1:0] OUT_518,	output reg [BIT - 1:0] OUT_519,	output reg [BIT - 1:0] OUT_520,	output reg [BIT - 1:0] OUT_521,	output reg [BIT - 1:0] OUT_522,	output reg [BIT - 1:0] OUT_523,	output reg [BIT - 1:0] OUT_524,	output reg [BIT - 1:0] OUT_525,	output reg [BIT - 1:0] OUT_526,	output reg [BIT - 1:0] OUT_527,	output reg [BIT - 1:0] OUT_528,	output reg [BIT - 1:0] OUT_529,	output reg [BIT - 1:0] OUT_530,	output reg [BIT - 1:0] OUT_531,	output reg [BIT - 1:0] OUT_532,	output reg [BIT - 1:0] OUT_533,	output reg [BIT - 1:0] OUT_534,	output reg [BIT - 1:0] OUT_535,	output reg [BIT - 1:0] OUT_536,	output reg [BIT - 1:0] OUT_537,	output reg [BIT - 1:0] OUT_538,	output reg [BIT - 1:0] OUT_539,	output reg [BIT - 1:0] OUT_540,	output reg [BIT - 1:0] OUT_541,	output reg [BIT - 1:0] OUT_542,	output reg [BIT - 1:0] OUT_543,	output reg [BIT - 1:0] OUT_544,	output reg [BIT - 1:0] OUT_545,	output reg [BIT - 1:0] OUT_546,	output reg [BIT - 1:0] OUT_547,	output reg [BIT - 1:0] OUT_548,	output reg [BIT - 1:0] OUT_549,	output reg [BIT - 1:0] OUT_550,	output reg [BIT - 1:0] OUT_551,	output reg [BIT - 1:0] OUT_552,	output reg [BIT - 1:0] OUT_553,	output reg [BIT - 1:0] OUT_554,	output reg [BIT - 1:0] OUT_555,	output reg [BIT - 1:0] OUT_556,	output reg [BIT - 1:0] OUT_557,	output reg [BIT - 1:0] OUT_558,	output reg [BIT - 1:0] OUT_559,	output reg [BIT - 1:0] OUT_560,	output reg [BIT - 1:0] OUT_561,	output reg [BIT - 1:0] OUT_562,	output reg [BIT - 1:0] OUT_563,	output reg [BIT - 1:0] OUT_564,	output reg [BIT - 1:0] OUT_565,	output reg [BIT - 1:0] OUT_566,	output reg [BIT - 1:0] OUT_567,	output reg [BIT - 1:0] OUT_568,	output reg [BIT - 1:0] OUT_569,	output reg [BIT - 1:0] OUT_570,	output reg [BIT - 1:0] OUT_571,	output reg [BIT - 1:0] OUT_572,	output reg [BIT - 1:0] OUT_573,	output reg [BIT - 1:0] OUT_574,	output reg [BIT - 1:0] OUT_575,	output reg [BIT - 1:0] OUT_576,	output reg [BIT - 1:0] OUT_577,	output reg [BIT - 1:0] OUT_578,	output reg [BIT - 1:0] OUT_579,	output reg [BIT - 1:0] OUT_580,	output reg [BIT - 1:0] OUT_581,	output reg [BIT - 1:0] OUT_582,	output reg [BIT - 1:0] OUT_583,	output reg [BIT - 1:0] OUT_584,	output reg [BIT - 1:0] OUT_585,	output reg [BIT - 1:0] OUT_586,	output reg [BIT - 1:0] OUT_587,	output reg [BIT - 1:0] OUT_588,	output reg [BIT - 1:0] OUT_589,	output reg [BIT - 1:0] OUT_590,	output reg [BIT - 1:0] OUT_591,	output reg [BIT - 1:0] OUT_592,	output reg [BIT - 1:0] OUT_593,	output reg [BIT - 1:0] OUT_594,	output reg [BIT - 1:0] OUT_595,	output reg [BIT - 1:0] OUT_596,	output reg [BIT - 1:0] OUT_597,	output reg [BIT - 1:0] OUT_598,	output reg [BIT - 1:0] OUT_599,	output reg [BIT - 1:0] OUT_600,	output reg [BIT - 1:0] OUT_601,	output reg [BIT - 1:0] OUT_602,	output reg [BIT - 1:0] OUT_603,	output reg [BIT - 1:0] OUT_604,	output reg [BIT - 1:0] OUT_605,	output reg [BIT - 1:0] OUT_606,	output reg [BIT - 1:0] OUT_607,	output reg [BIT - 1:0] OUT_608,	output reg [BIT - 1:0] OUT_609,	output reg [BIT - 1:0] OUT_610,	output reg [BIT - 1:0] OUT_611,	output reg [BIT - 1:0] OUT_612,	output reg [BIT - 1:0] OUT_613,	output reg [BIT - 1:0] OUT_614,	output reg [BIT - 1:0] OUT_615,	output reg [BIT - 1:0] OUT_616,	output reg [BIT - 1:0] OUT_617,	output reg [BIT - 1:0] OUT_618,	output reg [BIT - 1:0] OUT_619,	output reg [BIT - 1:0] OUT_620,	output reg [BIT - 1:0] OUT_621,	output reg [BIT - 1:0] OUT_622,	output reg [BIT - 1:0] OUT_623,	output reg [BIT - 1:0] OUT_624,	output reg [BIT - 1:0] OUT_625,	output reg [BIT - 1:0] OUT_626,	output reg [BIT - 1:0] OUT_627,	output reg [BIT - 1:0] OUT_628,	output reg [BIT - 1:0] OUT_629,	output reg [BIT - 1:0] OUT_630,	output reg [BIT - 1:0] OUT_631,	output reg [BIT - 1:0] OUT_632,	output reg [BIT - 1:0] OUT_633,	output reg [BIT - 1:0] OUT_634,	output reg [BIT - 1:0] OUT_635,	output reg [BIT - 1:0] OUT_636,	output reg [BIT - 1:0] OUT_637,	output reg [BIT - 1:0] OUT_638,	output reg [BIT - 1:0] OUT_639,	output reg [BIT - 1:0] OUT_640,	output reg [BIT - 1:0] OUT_641,	output reg [BIT - 1:0] OUT_642,	output reg [BIT - 1:0] OUT_643,	output reg [BIT - 1:0] OUT_644,	output reg [BIT - 1:0] OUT_645,	output reg [BIT - 1:0] OUT_646,	output reg [BIT - 1:0] OUT_647,	output reg [BIT - 1:0] OUT_648,	output reg [BIT - 1:0] OUT_649,	output reg [BIT - 1:0] OUT_650,	output reg [BIT - 1:0] OUT_651,	output reg [BIT - 1:0] OUT_652,	output reg [BIT - 1:0] OUT_653,	output reg [BIT - 1:0] OUT_654,	output reg [BIT - 1:0] OUT_655,	output reg [BIT - 1:0] OUT_656,	output reg [BIT - 1:0] OUT_657,	output reg [BIT - 1:0] OUT_658,	output reg [BIT - 1:0] OUT_659,	output reg [BIT - 1:0] OUT_660,	output reg [BIT - 1:0] OUT_661,	output reg [BIT - 1:0] OUT_662,	output reg [BIT - 1:0] OUT_663,	output reg [BIT - 1:0] OUT_664,	output reg [BIT - 1:0] OUT_665,	output reg [BIT - 1:0] OUT_666,	output reg [BIT - 1:0] OUT_667,	output reg [BIT - 1:0] OUT_668,	output reg [BIT - 1:0] OUT_669,	output reg [BIT - 1:0] OUT_670,	output reg [BIT - 1:0] OUT_671,	output reg [BIT - 1:0] OUT_672,	output reg [BIT - 1:0] OUT_673,	output reg [BIT - 1:0] OUT_674,	output reg [BIT - 1:0] OUT_675,	output reg [BIT - 1:0] OUT_676,	output reg [BIT - 1:0] OUT_677,	output reg [BIT - 1:0] OUT_678,	output reg [BIT - 1:0] OUT_679,	output reg [BIT - 1:0] OUT_680,	output reg [BIT - 1:0] OUT_681,	output reg [BIT - 1:0] OUT_682,	output reg [BIT - 1:0] OUT_683,	output reg [BIT - 1:0] OUT_684,	output reg [BIT - 1:0] OUT_685,	output reg [BIT - 1:0] OUT_686,	output reg [BIT - 1:0] OUT_687,	output reg [BIT - 1:0] OUT_688,	output reg [BIT - 1:0] OUT_689,	output reg [BIT - 1:0] OUT_690,	output reg [BIT - 1:0] OUT_691,	output reg [BIT - 1:0] OUT_692,	output reg [BIT - 1:0] OUT_693,	output reg [BIT - 1:0] OUT_694,	output reg [BIT - 1:0] OUT_695,	output reg [BIT - 1:0] OUT_696,	output reg [BIT - 1:0] OUT_697,	output reg [BIT - 1:0] OUT_698,	output reg [BIT - 1:0] OUT_699,	output reg [BIT - 1:0] OUT_700,	output reg [BIT - 1:0] OUT_701,	output reg [BIT - 1:0] OUT_702,	output reg [BIT - 1:0] OUT_703,	output reg [BIT - 1:0] OUT_704,	output reg [BIT - 1:0] OUT_705,	output reg [BIT - 1:0] OUT_706,	output reg [BIT - 1:0] OUT_707,	output reg [BIT - 1:0] OUT_708,	output reg [BIT - 1:0] OUT_709,	output reg [BIT - 1:0] OUT_710,	output reg [BIT - 1:0] OUT_711,	output reg [BIT - 1:0] OUT_712,	output reg [BIT - 1:0] OUT_713,	output reg [BIT - 1:0] OUT_714,	output reg [BIT - 1:0] OUT_715,	output reg [BIT - 1:0] OUT_716,	output reg [BIT - 1:0] OUT_717,	output reg [BIT - 1:0] OUT_718,	output reg [BIT - 1:0] OUT_719,	output reg [BIT - 1:0] OUT_720,	output reg [BIT - 1:0] OUT_721,	output reg [BIT - 1:0] OUT_722,	output reg [BIT - 1:0] OUT_723,	output reg [BIT - 1:0] OUT_724,	output reg [BIT - 1:0] OUT_725,	output reg [BIT - 1:0] OUT_726,	output reg [BIT - 1:0] OUT_727,	output reg [BIT - 1:0] OUT_728,	output reg [BIT - 1:0] OUT_729,	output reg [BIT - 1:0] OUT_730,	output reg [BIT - 1:0] OUT_731,	output reg [BIT - 1:0] OUT_732,	output reg [BIT - 1:0] OUT_733,	output reg [BIT - 1:0] OUT_734,	output reg [BIT - 1:0] OUT_735,	output reg [BIT - 1:0] OUT_736,	output reg [BIT - 1:0] OUT_737,	output reg [BIT - 1:0] OUT_738,	output reg [BIT - 1:0] OUT_739,	output reg [BIT - 1:0] OUT_740,	output reg [BIT - 1:0] OUT_741,	output reg [BIT - 1:0] OUT_742,	output reg [BIT - 1:0] OUT_743,	output reg [BIT - 1:0] OUT_744,	output reg [BIT - 1:0] OUT_745,	output reg [BIT - 1:0] OUT_746,	output reg [BIT - 1:0] OUT_747,	output reg [BIT - 1:0] OUT_748,	output reg [BIT - 1:0] OUT_749,	output reg [BIT - 1:0] OUT_750,	output reg [BIT - 1:0] OUT_751,	output reg [BIT - 1:0] OUT_752,	output reg [BIT - 1:0] OUT_753,	output reg [BIT - 1:0] OUT_754,	output reg [BIT - 1:0] OUT_755,	output reg [BIT - 1:0] OUT_756,	output reg [BIT - 1:0] OUT_757,	output reg [BIT - 1:0] OUT_758,	output reg [BIT - 1:0] OUT_759,	output reg [BIT - 1:0] OUT_760,	output reg [BIT - 1:0] OUT_761,	output reg [BIT - 1:0] OUT_762,	output reg [BIT - 1:0] OUT_763,	output reg [BIT - 1:0] OUT_764,	output reg [BIT - 1:0] OUT_765,	output reg [BIT - 1:0] OUT_766,	output reg [BIT - 1:0] OUT_767,	output reg [BIT - 1:0] OUT_768,	output reg [BIT - 1:0] OUT_769,	output reg [BIT - 1:0] OUT_770,	output reg [BIT - 1:0] OUT_771,	output reg [BIT - 1:0] OUT_772,	output reg [BIT - 1:0] OUT_773,	output reg [BIT - 1:0] OUT_774,	output reg [BIT - 1:0] OUT_775,	output reg [BIT - 1:0] OUT_776,	output reg [BIT - 1:0] OUT_777,	output reg [BIT - 1:0] OUT_778,	output reg [BIT - 1:0] OUT_779,	output reg [BIT - 1:0] OUT_780,	output reg [BIT - 1:0] OUT_781,	output reg [BIT - 1:0] OUT_782,	output reg [BIT - 1:0] OUT_783,	output reg [BIT - 1:0] OUT_784,	output reg [BIT - 1:0] OUT_785,	output reg [BIT - 1:0] OUT_786,	output reg [BIT - 1:0] OUT_787,	output reg [BIT - 1:0] OUT_788,	output reg [BIT - 1:0] OUT_789,	output reg [BIT - 1:0] OUT_790,	output reg [BIT - 1:0] OUT_791,	output reg [BIT - 1:0] OUT_792,	output reg [BIT - 1:0] OUT_793,	output reg [BIT - 1:0] OUT_794,	output reg [BIT - 1:0] OUT_795,	output reg [BIT - 1:0] OUT_796,	output reg [BIT - 1:0] OUT_797,	output reg [BIT - 1:0] OUT_798,	output reg [BIT - 1:0] OUT_799,	output reg [BIT - 1:0] OUT_800,	output reg [BIT - 1:0] OUT_801,	output reg [BIT - 1:0] OUT_802,	output reg [BIT - 1:0] OUT_803,	output reg [BIT - 1:0] OUT_804,	output reg [BIT - 1:0] OUT_805,	output reg [BIT - 1:0] OUT_806,	output reg [BIT - 1:0] OUT_807,	output reg [BIT - 1:0] OUT_808,	output reg [BIT - 1:0] OUT_809,	output reg [BIT - 1:0] OUT_810,	output reg [BIT - 1:0] OUT_811,	output reg [BIT - 1:0] OUT_812,	output reg [BIT - 1:0] OUT_813,	output reg [BIT - 1:0] OUT_814,	output reg [BIT - 1:0] OUT_815,	output reg [BIT - 1:0] OUT_816,	output reg [BIT - 1:0] OUT_817,	output reg [BIT - 1:0] OUT_818,	output reg [BIT - 1:0] OUT_819,	output reg [BIT - 1:0] OUT_820,	output reg [BIT - 1:0] OUT_821,	output reg [BIT - 1:0] OUT_822,	output reg [BIT - 1:0] OUT_823,	output reg [BIT - 1:0] OUT_824,	output reg [BIT - 1:0] OUT_825,	output reg [BIT - 1:0] OUT_826,	output reg [BIT - 1:0] OUT_827,	output reg [BIT - 1:0] OUT_828,	output reg [BIT - 1:0] OUT_829,	output reg [BIT - 1:0] OUT_830,	output reg [BIT - 1:0] OUT_831,	output reg [BIT - 1:0] OUT_832,	output reg [BIT - 1:0] OUT_833,	output reg [BIT - 1:0] OUT_834,	output reg [BIT - 1:0] OUT_835,	output reg [BIT - 1:0] OUT_836,	output reg [BIT - 1:0] OUT_837,	output reg [BIT - 1:0] OUT_838,	output reg [BIT - 1:0] OUT_839,	output reg [BIT - 1:0] OUT_840,	output reg [BIT - 1:0] OUT_841,	output reg [BIT - 1:0] OUT_842,	output reg [BIT - 1:0] OUT_843,	output reg [BIT - 1:0] OUT_844,	output reg [BIT - 1:0] OUT_845,	output reg [BIT - 1:0] OUT_846,	output reg [BIT - 1:0] OUT_847,	output reg [BIT - 1:0] OUT_848,	output reg [BIT - 1:0] OUT_849,	output reg [BIT - 1:0] OUT_850,	output reg [BIT - 1:0] OUT_851,	output reg [BIT - 1:0] OUT_852,	output reg [BIT - 1:0] OUT_853,	output reg [BIT - 1:0] OUT_854,	output reg [BIT - 1:0] OUT_855,	output reg [BIT - 1:0] OUT_856,	output reg [BIT - 1:0] OUT_857,	output reg [BIT - 1:0] OUT_858,	output reg [BIT - 1:0] OUT_859,	output reg [BIT - 1:0] OUT_860,	output reg [BIT - 1:0] OUT_861,	output reg [BIT - 1:0] OUT_862,	output reg [BIT - 1:0] OUT_863,	output reg [BIT - 1:0] OUT_864,	output reg [BIT - 1:0] OUT_865,	output reg [BIT - 1:0] OUT_866,	output reg [BIT - 1:0] OUT_867,	output reg [BIT - 1:0] OUT_868,	output reg [BIT - 1:0] OUT_869,	output reg [BIT - 1:0] OUT_870,	output reg [BIT - 1:0] OUT_871,	output reg [BIT - 1:0] OUT_872,	output reg [BIT - 1:0] OUT_873,	output reg [BIT - 1:0] OUT_874,	output reg [BIT - 1:0] OUT_875,	output reg [BIT - 1:0] OUT_876,	output reg [BIT - 1:0] OUT_877,	output reg [BIT - 1:0] OUT_878,	output reg [BIT - 1:0] OUT_879,	output reg [BIT - 1:0] OUT_880,	output reg [BIT - 1:0] OUT_881,	output reg [BIT - 1:0] OUT_882,	output reg [BIT - 1:0] OUT_883,	output reg [BIT - 1:0] OUT_884,	output reg [BIT - 1:0] OUT_885,	output reg [BIT - 1:0] OUT_886,	output reg [BIT - 1:0] OUT_887,	output reg [BIT - 1:0] OUT_888,	output reg [BIT - 1:0] OUT_889,	output reg [BIT - 1:0] OUT_890,	output reg [BIT - 1:0] OUT_891,	output reg [BIT - 1:0] OUT_892,	output reg [BIT - 1:0] OUT_893,	output reg [BIT - 1:0] OUT_894,	output reg [BIT - 1:0] OUT_895,	output reg [BIT - 1:0] OUT_896,	output reg [BIT - 1:0] OUT_897,	output reg [BIT - 1:0] OUT_898,	output reg [BIT - 1:0] OUT_899,	output reg [BIT - 1:0] OUT_900,	output reg [BIT - 1:0] OUT_901,	output reg [BIT - 1:0] OUT_902,	output reg [BIT - 1:0] OUT_903,	output reg [BIT - 1:0] OUT_904,	output reg [BIT - 1:0] OUT_905,	output reg [BIT - 1:0] OUT_906,	output reg [BIT - 1:0] OUT_907,	output reg [BIT - 1:0] OUT_908,	output reg [BIT - 1:0] OUT_909,	output reg [BIT - 1:0] OUT_910,	output reg [BIT - 1:0] OUT_911,	output reg [BIT - 1:0] OUT_912,	output reg [BIT - 1:0] OUT_913,	output reg [BIT - 1:0] OUT_914,	output reg [BIT - 1:0] OUT_915,	output reg [BIT - 1:0] OUT_916,	output reg [BIT - 1:0] OUT_917,	output reg [BIT - 1:0] OUT_918,	output reg [BIT - 1:0] OUT_919,	output reg [BIT - 1:0] OUT_920,	output reg [BIT - 1:0] OUT_921,	output reg [BIT - 1:0] OUT_922,	output reg [BIT - 1:0] OUT_923,	output reg [BIT - 1:0] OUT_924,	output reg [BIT - 1:0] OUT_925,	output reg [BIT - 1:0] OUT_926,	output reg [BIT - 1:0] OUT_927,	output reg [BIT - 1:0] OUT_928,	output reg [BIT - 1:0] OUT_929,	output reg [BIT - 1:0] OUT_930,	output reg [BIT - 1:0] OUT_931,	output reg [BIT - 1:0] OUT_932,	output reg [BIT - 1:0] OUT_933,	output reg [BIT - 1:0] OUT_934,	output reg [BIT - 1:0] OUT_935,	output reg [BIT - 1:0] OUT_936,	output reg [BIT - 1:0] OUT_937,	output reg [BIT - 1:0] OUT_938,	output reg [BIT - 1:0] OUT_939,	output reg [BIT - 1:0] OUT_940,	output reg [BIT - 1:0] OUT_941,	output reg [BIT - 1:0] OUT_942,	output reg [BIT - 1:0] OUT_943,	output reg [BIT - 1:0] OUT_944,	output reg [BIT - 1:0] OUT_945,	output reg [BIT - 1:0] OUT_946,	output reg [BIT - 1:0] OUT_947,	output reg [BIT - 1:0] OUT_948,	output reg [BIT - 1:0] OUT_949,	output reg [BIT - 1:0] OUT_950,	output reg [BIT - 1:0] OUT_951,	output reg [BIT - 1:0] OUT_952,	output reg [BIT - 1:0] OUT_953,	output reg [BIT - 1:0] OUT_954,	output reg [BIT - 1:0] OUT_955,	output reg [BIT - 1:0] OUT_956,	output reg [BIT - 1:0] OUT_957,	output reg [BIT - 1:0] OUT_958,	output reg [BIT - 1:0] OUT_959,	output reg [BIT - 1:0] OUT_960,	output reg [BIT - 1:0] OUT_961,	output reg [BIT - 1:0] OUT_962,	output reg [BIT - 1:0] OUT_963,	output reg [BIT - 1:0] OUT_964,	output reg [BIT - 1:0] OUT_965,	output reg [BIT - 1:0] OUT_966,	output reg [BIT - 1:0] OUT_967,	output reg [BIT - 1:0] OUT_968,	output reg [BIT - 1:0] OUT_969,	output reg [BIT - 1:0] OUT_970,	output reg [BIT - 1:0] OUT_971,	output reg [BIT - 1:0] OUT_972,	output reg [BIT - 1:0] OUT_973,	output reg [BIT - 1:0] OUT_974,	output reg [BIT - 1:0] OUT_975,	output reg [BIT - 1:0] OUT_976,	output reg [BIT - 1:0] OUT_977,	output reg [BIT - 1:0] OUT_978,	output reg [BIT - 1:0] OUT_979,	output reg [BIT - 1:0] OUT_980,	output reg [BIT - 1:0] OUT_981,	output reg [BIT - 1:0] OUT_982,	output reg [BIT - 1:0] OUT_983,	output reg [BIT - 1:0] OUT_984,	output reg [BIT - 1:0] OUT_985,	output reg [BIT - 1:0] OUT_986,	output reg [BIT - 1:0] OUT_987,	output reg [BIT - 1:0] OUT_988,	output reg [BIT - 1:0] OUT_989,	output reg [BIT - 1:0] OUT_990,	output reg [BIT - 1:0] OUT_991,	output reg [BIT - 1:0] OUT_992,	output reg [BIT - 1:0] OUT_993,	output reg [BIT - 1:0] OUT_994,	output reg [BIT - 1:0] OUT_995,	output reg [BIT - 1:0] OUT_996,	output reg [BIT - 1:0] OUT_997,	output reg [BIT - 1:0] OUT_998,	output reg [BIT - 1:0] OUT_999,	output reg [BIT - 1:0] OUT_1000,	output reg [BIT - 1:0] OUT_1001,	output reg [BIT - 1:0] OUT_1002,	output reg [BIT - 1:0] OUT_1003,	output reg [BIT - 1:0] OUT_1004,	output reg [BIT - 1:0] OUT_1005,	output reg [BIT - 1:0] OUT_1006,	output reg [BIT - 1:0] OUT_1007,	output reg [BIT - 1:0] OUT_1008,	output reg [BIT - 1:0] OUT_1009,	output reg [BIT - 1:0] OUT_1010,	output reg [BIT - 1:0] OUT_1011,	output reg [BIT - 1:0] OUT_1012,	output reg [BIT - 1:0] OUT_1013,	output reg [BIT - 1:0] OUT_1014,	output reg [BIT - 1:0] OUT_1015,	output reg [BIT - 1:0] OUT_1016,	output reg [BIT - 1:0] OUT_1017,	output reg [BIT - 1:0] OUT_1018,	output reg [BIT - 1:0] OUT_1019,	output reg [BIT - 1:0] OUT_1020,	output reg [BIT - 1:0] OUT_1021,	output reg [BIT - 1:0] OUT_1022,	output reg [BIT - 1:0] OUT_1023,	output reg [BIT - 1:0] OUT_1024);	integer x, y;
	reg [BIT - 1:0] inform_R [1024-1:0][11-1:0];	reg [BIT - 1:0] inform_L [1024-1:0][11-1:0];	localparam IDLE = 2'b00;	localparam BUSY_LEFT = 2'b01;	localparam BUSY_RIGHT = 2'b10;	reg [1:0] bp_state,bp_next_state;	reg [10-1:0] cell_enable,w2r,w2r_delay;	reg left_over_flag,right_over_flag,init_over_flag;	wire bp_over_flag;	reg [6:0]itera_time;
	always @(posedge clk or negedge rst_n) begin		if (!rst_n) begin			bp_state <= IDLE;		end		else begin			bp_state <= bp_next_state;		end	end
	always @(*) begin		case (bp_state)			IDLE:			if (init_over_flag) begin				bp_next_state <= BUSY_LEFT;			end			else begin				bp_next_state <= IDLE;			end
			BUSY_LEFT:			if (left_over_flag) begin				bp_next_state <= BUSY_RIGHT;			end			else begin				 bp_next_state <= BUSY_LEFT;			end
			BUSY_RIGHT:			if (bp_over_flag) begin				bp_next_state <= IDLE;			end			else if (right_over_flag) begin				bp_next_state <= BUSY_LEFT;			end			else begin				 bp_next_state <= BUSY_RIGHT;			end
			default: bp_next_state <= IDLE;		endcase	end
	reg [1:0] clk_counter;
	always @(posedge clk) begin		case (bp_next_state)			IDLE:			begin				left_over_flag <= 0;				right_over_flag <= 0;				itera_time <= 7'b0;				clk_counter <= 2'b0;				if (start) begin					cell_enable <=10'b1;					w2r <= 10;					init_over_flag <= 1;					en_busy <= 1;				end				else begin					cell_enable <=10'b0;					w2r <= 0;					init_over_flag <= 0;					en_busy <= 0;				end			end
			BUSY_LEFT:			begin				init_over_flag <= 0;				en_busy <= 1;				right_over_flag <= 0;				if (clk_counter == 2'b11) begin					clk_counter <= 2'b00;					if (cell_enable == 512) begin						left_over_flag <= 1;						cell_enable <= cell_enable >> 1;						w2r <= w2r + 1;					end					else begin						left_over_flag <= 0;						cell_enable <= cell_enable << 1;						w2r <= w2r - 1;					end				end				else begin					clk_counter <= clk_counter + 1;				end			end
			BUSY_RIGHT:			begin				en_busy <= 1;				left_over_flag <= 0;				if (clk_counter == 2'b11) begin					clk_counter <= 2'b00;					if (cell_enable == 1) begin						right_over_flag <= 1;						itera_time <= itera_time + 1;						cell_enable <= cell_enable << 1;						w2r <= w2r - 1;					end					else begin						right_over_flag <= 0;						cell_enable <= cell_enable >> 1;						w2r <= w2r + 1;					end				end				else begin					clk_counter <= clk_counter + 1;				end			end
			default:			begin				left_over_flag <= 0;				right_over_flag <= 0;				itera_time <= 7'b0;				clk_counter <= 2'b0;				if (start) begin					cell_enable <=10'b1;					w2r <= 10;					init_over_flag <= 1;					en_busy <= 1;				end				else begin					cell_enable <=10'b0;					w2r <= 0;					init_over_flag <= 0;					en_busy <= 0;				end			end
		endcase	end
	reg[BIT - 1:0] r_cell_reg[1024-1:0];	reg[BIT - 1:0] l_cell_reg[1024-1:0];	wire[BIT - 1:0] r_cell_wire[1024-1:0];	wire[BIT - 1:0] l_cell_wire[1024-1:0];
	always @(posedge clk) begin		case (bp_next_state)			IDLE:			begin				if (start) begin					inform_R [0][0] <= 8'b0111_1111;					inform_R [1][0] <= 8'b0111_1111;					inform_R [2][0] <= 8'b0111_1111;					inform_R [3][0] <= 8'b0111_1111;					inform_R [4][0] <= 8'b0111_1111;					inform_R [5][0] <= 8'b0111_1111;					inform_R [6][0] <= 8'b0111_1111;					inform_R [7][0] <= 8'b0111_1111;					inform_R [8][0] <= 8'b0111_1111;					inform_R [9][0] <= 8'b0111_1111;					inform_R [10][0] <= 8'b0111_1111;					inform_R [11][0] <= 8'b0111_1111;					inform_R [12][0] <= 8'b0111_1111;					inform_R [13][0] <= 8'b0111_1111;					inform_R [14][0] <= 8'b0111_1111;					inform_R [15][0] <= 8'b0111_1111;					inform_R [16][0] <= 8'b0111_1111;					inform_R [17][0] <= 8'b0111_1111;					inform_R [18][0] <= 8'b0111_1111;					inform_R [19][0] <= 8'b0111_1111;					inform_R [20][0] <= 8'b0111_1111;					inform_R [21][0] <= 8'b0111_1111;					inform_R [22][0] <= 8'b0111_1111;					inform_R [23][0] <= 8'b0111_1111;					inform_R [24][0] <= 8'b0111_1111;					inform_R [25][0] <= 8'b0111_1111;					inform_R [26][0] <= 8'b0111_1111;					inform_R [27][0] <= 8'b0111_1111;					inform_R [28][0] <= 8'b0111_1111;					inform_R [29][0] <= 8'b0111_1111;					inform_R [30][0] <= 8'b0111_1111;					inform_R [31][0] <= 8'b0111_1111;					inform_R [32][0] <= 8'b0111_1111;					inform_R [33][0] <= 8'b0111_1111;					inform_R [34][0] <= 8'b0111_1111;					inform_R [35][0] <= 8'b0111_1111;					inform_R [36][0] <= 8'b0111_1111;					inform_R [37][0] <= 8'b0111_1111;					inform_R [38][0] <= 8'b0111_1111;					inform_R [39][0] <= 8'b0111_1111;					inform_R [40][0] <= 8'b0111_1111;					inform_R [41][0] <= 8'b0111_1111;					inform_R [42][0] <= 8'b0111_1111;					inform_R [43][0] <= 8'b0111_1111;					inform_R [44][0] <= 8'b0111_1111;					inform_R [45][0] <= 8'b0111_1111;					inform_R [46][0] <= 8'b0111_1111;					inform_R [47][0] <= 8'b0111_1111;					inform_R [48][0] <= 8'b0111_1111;					inform_R [49][0] <= 8'b0111_1111;					inform_R [50][0] <= 8'b0111_1111;					inform_R [51][0] <= 8'b0111_1111;					inform_R [52][0] <= 8'b0111_1111;					inform_R [53][0] <= 8'b0111_1111;					inform_R [54][0] <= 8'b0111_1111;					inform_R [55][0] <= 8'b0111_1111;					inform_R [56][0] <= 8'b0111_1111;					inform_R [57][0] <= 8'b0111_1111;					inform_R [58][0] <= 8'b0111_1111;					inform_R [59][0] <= 8'b0111_1111;					inform_R [60][0] <= 8'b0111_1111;					inform_R [61][0] <= 8'b0111_1111;					inform_R [62][0] <= 8'b0111_1111;					inform_R [63][0] <= 8'b0000_0000;					inform_R [64][0] <= 8'b0111_1111;					inform_R [65][0] <= 8'b0111_1111;					inform_R [66][0] <= 8'b0111_1111;					inform_R [67][0] <= 8'b0111_1111;					inform_R [68][0] <= 8'b0111_1111;					inform_R [69][0] <= 8'b0111_1111;					inform_R [70][0] <= 8'b0111_1111;					inform_R [71][0] <= 8'b0111_1111;					inform_R [72][0] <= 8'b0111_1111;					inform_R [73][0] <= 8'b0111_1111;					inform_R [74][0] <= 8'b0111_1111;					inform_R [75][0] <= 8'b0111_1111;					inform_R [76][0] <= 8'b0111_1111;					inform_R [77][0] <= 8'b0111_1111;					inform_R [78][0] <= 8'b0111_1111;					inform_R [79][0] <= 8'b0111_1111;					inform_R [80][0] <= 8'b0111_1111;					inform_R [81][0] <= 8'b0111_1111;					inform_R [82][0] <= 8'b0111_1111;					inform_R [83][0] <= 8'b0111_1111;					inform_R [84][0] <= 8'b0111_1111;					inform_R [85][0] <= 8'b0111_1111;					inform_R [86][0] <= 8'b0111_1111;					inform_R [87][0] <= 8'b0111_1111;					inform_R [88][0] <= 8'b0111_1111;					inform_R [89][0] <= 8'b0111_1111;					inform_R [90][0] <= 8'b0111_1111;					inform_R [91][0] <= 8'b0111_1111;					inform_R [92][0] <= 8'b0111_1111;					inform_R [93][0] <= 8'b0111_1111;					inform_R [94][0] <= 8'b0111_1111;					inform_R [95][0] <= 8'b0000_0000;					inform_R [96][0] <= 8'b0111_1111;					inform_R [97][0] <= 8'b0111_1111;					inform_R [98][0] <= 8'b0111_1111;					inform_R [99][0] <= 8'b0111_1111;					inform_R [100][0] <= 8'b0111_1111;					inform_R [101][0] <= 8'b0111_1111;					inform_R [102][0] <= 8'b0111_1111;					inform_R [103][0] <= 8'b0111_1111;					inform_R [104][0] <= 8'b0111_1111;					inform_R [105][0] <= 8'b0111_1111;					inform_R [106][0] <= 8'b0111_1111;					inform_R [107][0] <= 8'b0111_1111;					inform_R [108][0] <= 8'b0111_1111;					inform_R [109][0] <= 8'b0111_1111;					inform_R [110][0] <= 8'b0111_1111;					inform_R [111][0] <= 8'b0000_0000;					inform_R [112][0] <= 8'b0111_1111;					inform_R [113][0] <= 8'b0111_1111;					inform_R [114][0] <= 8'b0111_1111;					inform_R [115][0] <= 8'b0111_1111;					inform_R [116][0] <= 8'b0111_1111;					inform_R [117][0] <= 8'b0111_1111;					inform_R [118][0] <= 8'b0111_1111;					inform_R [119][0] <= 8'b0000_0000;					inform_R [120][0] <= 8'b0111_1111;					inform_R [121][0] <= 8'b0111_1111;					inform_R [122][0] <= 8'b0000_0000;					inform_R [123][0] <= 8'b0000_0000;					inform_R [124][0] <= 8'b0000_0000;					inform_R [125][0] <= 8'b0000_0000;					inform_R [126][0] <= 8'b0000_0000;					inform_R [127][0] <= 8'b0000_0000;					inform_R [128][0] <= 8'b0111_1111;					inform_R [129][0] <= 8'b0111_1111;					inform_R [130][0] <= 8'b0111_1111;					inform_R [131][0] <= 8'b0111_1111;					inform_R [132][0] <= 8'b0111_1111;					inform_R [133][0] <= 8'b0111_1111;					inform_R [134][0] <= 8'b0111_1111;					inform_R [135][0] <= 8'b0111_1111;					inform_R [136][0] <= 8'b0111_1111;					inform_R [137][0] <= 8'b0111_1111;					inform_R [138][0] <= 8'b0111_1111;					inform_R [139][0] <= 8'b0111_1111;					inform_R [140][0] <= 8'b0111_1111;					inform_R [141][0] <= 8'b0111_1111;					inform_R [142][0] <= 8'b0111_1111;					inform_R [143][0] <= 8'b0111_1111;					inform_R [144][0] <= 8'b0111_1111;					inform_R [145][0] <= 8'b0111_1111;					inform_R [146][0] <= 8'b0111_1111;					inform_R [147][0] <= 8'b0111_1111;					inform_R [148][0] <= 8'b0111_1111;					inform_R [149][0] <= 8'b0111_1111;					inform_R [150][0] <= 8'b0111_1111;					inform_R [151][0] <= 8'b0111_1111;					inform_R [152][0] <= 8'b0111_1111;					inform_R [153][0] <= 8'b0111_1111;					inform_R [154][0] <= 8'b0111_1111;					inform_R [155][0] <= 8'b0111_1111;					inform_R [156][0] <= 8'b0111_1111;					inform_R [157][0] <= 8'b0111_1111;					inform_R [158][0] <= 8'b0111_1111;					inform_R [159][0] <= 8'b0000_0000;					inform_R [160][0] <= 8'b0111_1111;					inform_R [161][0] <= 8'b0111_1111;					inform_R [162][0] <= 8'b0111_1111;					inform_R [163][0] <= 8'b0111_1111;					inform_R [164][0] <= 8'b0111_1111;					inform_R [165][0] <= 8'b0111_1111;					inform_R [166][0] <= 8'b0111_1111;					inform_R [167][0] <= 8'b0111_1111;					inform_R [168][0] <= 8'b0111_1111;					inform_R [169][0] <= 8'b0111_1111;					inform_R [170][0] <= 8'b0111_1111;					inform_R [171][0] <= 8'b0111_1111;					inform_R [172][0] <= 8'b0111_1111;					inform_R [173][0] <= 8'b0111_1111;					inform_R [174][0] <= 8'b0111_1111;					inform_R [175][0] <= 8'b0000_0000;					inform_R [176][0] <= 8'b0111_1111;					inform_R [177][0] <= 8'b0111_1111;					inform_R [178][0] <= 8'b0111_1111;					inform_R [179][0] <= 8'b0111_1111;					inform_R [180][0] <= 8'b0111_1111;					inform_R [181][0] <= 8'b0000_0000;					inform_R [182][0] <= 8'b0000_0000;					inform_R [183][0] <= 8'b0000_0000;					inform_R [184][0] <= 8'b0111_1111;					inform_R [185][0] <= 8'b0000_0000;					inform_R [186][0] <= 8'b0000_0000;					inform_R [187][0] <= 8'b0000_0000;					inform_R [188][0] <= 8'b0000_0000;					inform_R [189][0] <= 8'b0000_0000;					inform_R [190][0] <= 8'b0000_0000;					inform_R [191][0] <= 8'b0000_0000;					inform_R [192][0] <= 8'b0111_1111;					inform_R [193][0] <= 8'b0111_1111;					inform_R [194][0] <= 8'b0111_1111;					inform_R [195][0] <= 8'b0111_1111;					inform_R [196][0] <= 8'b0111_1111;					inform_R [197][0] <= 8'b0111_1111;					inform_R [198][0] <= 8'b0111_1111;					inform_R [199][0] <= 8'b0000_0000;					inform_R [200][0] <= 8'b0111_1111;					inform_R [201][0] <= 8'b0111_1111;					inform_R [202][0] <= 8'b0111_1111;					inform_R [203][0] <= 8'b0000_0000;					inform_R [204][0] <= 8'b0111_1111;					inform_R [205][0] <= 8'b0000_0000;					inform_R [206][0] <= 8'b0000_0000;					inform_R [207][0] <= 8'b0000_0000;					inform_R [208][0] <= 8'b0111_1111;					inform_R [209][0] <= 8'b0111_1111;					inform_R [210][0] <= 8'b0111_1111;					inform_R [211][0] <= 8'b0000_0000;					inform_R [212][0] <= 8'b0111_1111;					inform_R [213][0] <= 8'b0000_0000;					inform_R [214][0] <= 8'b0000_0000;					inform_R [215][0] <= 8'b0000_0000;					inform_R [216][0] <= 8'b0111_1111;					inform_R [217][0] <= 8'b0000_0000;					inform_R [218][0] <= 8'b0000_0000;					inform_R [219][0] <= 8'b0000_0000;					inform_R [220][0] <= 8'b0000_0000;					inform_R [221][0] <= 8'b0000_0000;					inform_R [222][0] <= 8'b0000_0000;					inform_R [223][0] <= 8'b0000_0000;					inform_R [224][0] <= 8'b0111_1111;					inform_R [225][0] <= 8'b0111_1111;					inform_R [226][0] <= 8'b0111_1111;					inform_R [227][0] <= 8'b0000_0000;					inform_R [228][0] <= 8'b0111_1111;					inform_R [229][0] <= 8'b0000_0000;					inform_R [230][0] <= 8'b0000_0000;					inform_R [231][0] <= 8'b0000_0000;					inform_R [232][0] <= 8'b0000_0000;					inform_R [233][0] <= 8'b0000_0000;					inform_R [234][0] <= 8'b0000_0000;					inform_R [235][0] <= 8'b0000_0000;					inform_R [236][0] <= 8'b0000_0000;					inform_R [237][0] <= 8'b0000_0000;					inform_R [238][0] <= 8'b0000_0000;					inform_R [239][0] <= 8'b0000_0000;					inform_R [240][0] <= 8'b0000_0000;					inform_R [241][0] <= 8'b0000_0000;					inform_R [242][0] <= 8'b0000_0000;					inform_R [243][0] <= 8'b0000_0000;					inform_R [244][0] <= 8'b0000_0000;					inform_R [245][0] <= 8'b0000_0000;					inform_R [246][0] <= 8'b0000_0000;					inform_R [247][0] <= 8'b0000_0000;					inform_R [248][0] <= 8'b0000_0000;					inform_R [249][0] <= 8'b0000_0000;					inform_R [250][0] <= 8'b0000_0000;					inform_R [251][0] <= 8'b0000_0000;					inform_R [252][0] <= 8'b0000_0000;					inform_R [253][0] <= 8'b0000_0000;					inform_R [254][0] <= 8'b0000_0000;					inform_R [255][0] <= 8'b0000_0000;					inform_R [256][0] <= 8'b0111_1111;					inform_R [257][0] <= 8'b0111_1111;					inform_R [258][0] <= 8'b0111_1111;					inform_R [259][0] <= 8'b0111_1111;					inform_R [260][0] <= 8'b0111_1111;					inform_R [261][0] <= 8'b0111_1111;					inform_R [262][0] <= 8'b0111_1111;					inform_R [263][0] <= 8'b0111_1111;					inform_R [264][0] <= 8'b0111_1111;					inform_R [265][0] <= 8'b0111_1111;					inform_R [266][0] <= 8'b0111_1111;					inform_R [267][0] <= 8'b0111_1111;					inform_R [268][0] <= 8'b0111_1111;					inform_R [269][0] <= 8'b0111_1111;					inform_R [270][0] <= 8'b0111_1111;					inform_R [271][0] <= 8'b0111_1111;					inform_R [272][0] <= 8'b0111_1111;					inform_R [273][0] <= 8'b0111_1111;					inform_R [274][0] <= 8'b0111_1111;					inform_R [275][0] <= 8'b0111_1111;					inform_R [276][0] <= 8'b0111_1111;					inform_R [277][0] <= 8'b0111_1111;					inform_R [278][0] <= 8'b0111_1111;					inform_R [279][0] <= 8'b0000_0000;					inform_R [280][0] <= 8'b0111_1111;					inform_R [281][0] <= 8'b0111_1111;					inform_R [282][0] <= 8'b0111_1111;					inform_R [283][0] <= 8'b0000_0000;					inform_R [284][0] <= 8'b0111_1111;					inform_R [285][0] <= 8'b0000_0000;					inform_R [286][0] <= 8'b0000_0000;					inform_R [287][0] <= 8'b0000_0000;					inform_R [288][0] <= 8'b0111_1111;					inform_R [289][0] <= 8'b0111_1111;					inform_R [290][0] <= 8'b0111_1111;					inform_R [291][0] <= 8'b0111_1111;					inform_R [292][0] <= 8'b0111_1111;					inform_R [293][0] <= 8'b0111_1111;					inform_R [294][0] <= 8'b0111_1111;					inform_R [295][0] <= 8'b0000_0000;					inform_R [296][0] <= 8'b0111_1111;					inform_R [297][0] <= 8'b0111_1111;					inform_R [298][0] <= 8'b0111_1111;					inform_R [299][0] <= 8'b0000_0000;					inform_R [300][0] <= 8'b0111_1111;					inform_R [301][0] <= 8'b0000_0000;					inform_R [302][0] <= 8'b0000_0000;					inform_R [303][0] <= 8'b0000_0000;					inform_R [304][0] <= 8'b0111_1111;					inform_R [305][0] <= 8'b0111_1111;					inform_R [306][0] <= 8'b0111_1111;					inform_R [307][0] <= 8'b0000_0000;					inform_R [308][0] <= 8'b0111_1111;					inform_R [309][0] <= 8'b0000_0000;					inform_R [310][0] <= 8'b0000_0000;					inform_R [311][0] <= 8'b0000_0000;					inform_R [312][0] <= 8'b0111_1111;					inform_R [313][0] <= 8'b0000_0000;					inform_R [314][0] <= 8'b0000_0000;					inform_R [315][0] <= 8'b0000_0000;					inform_R [316][0] <= 8'b0000_0000;					inform_R [317][0] <= 8'b0000_0000;					inform_R [318][0] <= 8'b0000_0000;					inform_R [319][0] <= 8'b0000_0000;					inform_R [320][0] <= 8'b0111_1111;					inform_R [321][0] <= 8'b0111_1111;					inform_R [322][0] <= 8'b0111_1111;					inform_R [323][0] <= 8'b0111_1111;					inform_R [324][0] <= 8'b0111_1111;					inform_R [325][0] <= 8'b0111_1111;					inform_R [326][0] <= 8'b0111_1111;					inform_R [327][0] <= 8'b0000_0000;					inform_R [328][0] <= 8'b0111_1111;					inform_R [329][0] <= 8'b0111_1111;					inform_R [330][0] <= 8'b0111_1111;					inform_R [331][0] <= 8'b0000_0000;					inform_R [332][0] <= 8'b0111_1111;					inform_R [333][0] <= 8'b0000_0000;					inform_R [334][0] <= 8'b0000_0000;					inform_R [335][0] <= 8'b0000_0000;					inform_R [336][0] <= 8'b0111_1111;					inform_R [337][0] <= 8'b0111_1111;					inform_R [338][0] <= 8'b0111_1111;					inform_R [339][0] <= 8'b0000_0000;					inform_R [340][0] <= 8'b0000_0000;					inform_R [341][0] <= 8'b0000_0000;					inform_R [342][0] <= 8'b0000_0000;					inform_R [343][0] <= 8'b0000_0000;					inform_R [344][0] <= 8'b0000_0000;					inform_R [345][0] <= 8'b0000_0000;					inform_R [346][0] <= 8'b0000_0000;					inform_R [347][0] <= 8'b0000_0000;					inform_R [348][0] <= 8'b0000_0000;					inform_R [349][0] <= 8'b0000_0000;					inform_R [350][0] <= 8'b0000_0000;					inform_R [351][0] <= 8'b0000_0000;					inform_R [352][0] <= 8'b0111_1111;					inform_R [353][0] <= 8'b0000_0000;					inform_R [354][0] <= 8'b0000_0000;					inform_R [355][0] <= 8'b0000_0000;					inform_R [356][0] <= 8'b0000_0000;					inform_R [357][0] <= 8'b0000_0000;					inform_R [358][0] <= 8'b0000_0000;					inform_R [359][0] <= 8'b0000_0000;					inform_R [360][0] <= 8'b0000_0000;					inform_R [361][0] <= 8'b0000_0000;					inform_R [362][0] <= 8'b0000_0000;					inform_R [363][0] <= 8'b0000_0000;					inform_R [364][0] <= 8'b0000_0000;					inform_R [365][0] <= 8'b0000_0000;					inform_R [366][0] <= 8'b0000_0000;					inform_R [367][0] <= 8'b0000_0000;					inform_R [368][0] <= 8'b0000_0000;					inform_R [369][0] <= 8'b0000_0000;					inform_R [370][0] <= 8'b0000_0000;					inform_R [371][0] <= 8'b0000_0000;					inform_R [372][0] <= 8'b0000_0000;					inform_R [373][0] <= 8'b0000_0000;					inform_R [374][0] <= 8'b0000_0000;					inform_R [375][0] <= 8'b0000_0000;					inform_R [376][0] <= 8'b0000_0000;					inform_R [377][0] <= 8'b0000_0000;					inform_R [378][0] <= 8'b0000_0000;					inform_R [379][0] <= 8'b0000_0000;					inform_R [380][0] <= 8'b0000_0000;					inform_R [381][0] <= 8'b0000_0000;					inform_R [382][0] <= 8'b0000_0000;					inform_R [383][0] <= 8'b0000_0000;					inform_R [384][0] <= 8'b0111_1111;					inform_R [385][0] <= 8'b0111_1111;					inform_R [386][0] <= 8'b0111_1111;					inform_R [387][0] <= 8'b0111_1111;					inform_R [388][0] <= 8'b0111_1111;					inform_R [389][0] <= 8'b0111_1111;					inform_R [390][0] <= 8'b0000_0000;					inform_R [391][0] <= 8'b0000_0000;					inform_R [392][0] <= 8'b0111_1111;					inform_R [393][0] <= 8'b0000_0000;					inform_R [394][0] <= 8'b0000_0000;					inform_R [395][0] <= 8'b0000_0000;					inform_R [396][0] <= 8'b0000_0000;					inform_R [397][0] <= 8'b0000_0000;					inform_R [398][0] <= 8'b0000_0000;					inform_R [399][0] <= 8'b0000_0000;					inform_R [400][0] <= 8'b0111_1111;					inform_R [401][0] <= 8'b0000_0000;					inform_R [402][0] <= 8'b0000_0000;					inform_R [403][0] <= 8'b0000_0000;					inform_R [404][0] <= 8'b0000_0000;					inform_R [405][0] <= 8'b0000_0000;					inform_R [406][0] <= 8'b0000_0000;					inform_R [407][0] <= 8'b0000_0000;					inform_R [408][0] <= 8'b0000_0000;					inform_R [409][0] <= 8'b0000_0000;					inform_R [410][0] <= 8'b0000_0000;					inform_R [411][0] <= 8'b0000_0000;					inform_R [412][0] <= 8'b0000_0000;					inform_R [413][0] <= 8'b0000_0000;					inform_R [414][0] <= 8'b0000_0000;					inform_R [415][0] <= 8'b0000_0000;					inform_R [416][0] <= 8'b0111_1111;					inform_R [417][0] <= 8'b0000_0000;					inform_R [418][0] <= 8'b0000_0000;					inform_R [419][0] <= 8'b0000_0000;					inform_R [420][0] <= 8'b0000_0000;					inform_R [421][0] <= 8'b0000_0000;					inform_R [422][0] <= 8'b0000_0000;					inform_R [423][0] <= 8'b0000_0000;					inform_R [424][0] <= 8'b0000_0000;					inform_R [425][0] <= 8'b0000_0000;					inform_R [426][0] <= 8'b0000_0000;					inform_R [427][0] <= 8'b0000_0000;					inform_R [428][0] <= 8'b0000_0000;					inform_R [429][0] <= 8'b0000_0000;					inform_R [430][0] <= 8'b0000_0000;					inform_R [431][0] <= 8'b0000_0000;					inform_R [432][0] <= 8'b0000_0000;					inform_R [433][0] <= 8'b0000_0000;					inform_R [434][0] <= 8'b0000_0000;					inform_R [435][0] <= 8'b0000_0000;					inform_R [436][0] <= 8'b0000_0000;					inform_R [437][0] <= 8'b0000_0000;					inform_R [438][0] <= 8'b0000_0000;					inform_R [439][0] <= 8'b0000_0000;					inform_R [440][0] <= 8'b0000_0000;					inform_R [441][0] <= 8'b0000_0000;					inform_R [442][0] <= 8'b0000_0000;					inform_R [443][0] <= 8'b0000_0000;					inform_R [444][0] <= 8'b0000_0000;					inform_R [445][0] <= 8'b0000_0000;					inform_R [446][0] <= 8'b0000_0000;					inform_R [447][0] <= 8'b0000_0000;					inform_R [448][0] <= 8'b0000_0000;					inform_R [449][0] <= 8'b0000_0000;					inform_R [450][0] <= 8'b0000_0000;					inform_R [451][0] <= 8'b0000_0000;					inform_R [452][0] <= 8'b0000_0000;					inform_R [453][0] <= 8'b0000_0000;					inform_R [454][0] <= 8'b0000_0000;					inform_R [455][0] <= 8'b0000_0000;					inform_R [456][0] <= 8'b0000_0000;					inform_R [457][0] <= 8'b0000_0000;					inform_R [458][0] <= 8'b0000_0000;					inform_R [459][0] <= 8'b0000_0000;					inform_R [460][0] <= 8'b0000_0000;					inform_R [461][0] <= 8'b0000_0000;					inform_R [462][0] <= 8'b0000_0000;					inform_R [463][0] <= 8'b0000_0000;					inform_R [464][0] <= 8'b0000_0000;					inform_R [465][0] <= 8'b0000_0000;					inform_R [466][0] <= 8'b0000_0000;					inform_R [467][0] <= 8'b0000_0000;					inform_R [468][0] <= 8'b0000_0000;					inform_R [469][0] <= 8'b0000_0000;					inform_R [470][0] <= 8'b0000_0000;					inform_R [471][0] <= 8'b0000_0000;					inform_R [472][0] <= 8'b0000_0000;					inform_R [473][0] <= 8'b0000_0000;					inform_R [474][0] <= 8'b0000_0000;					inform_R [475][0] <= 8'b0000_0000;					inform_R [476][0] <= 8'b0000_0000;					inform_R [477][0] <= 8'b0000_0000;					inform_R [478][0] <= 8'b0000_0000;					inform_R [479][0] <= 8'b0000_0000;					inform_R [480][0] <= 8'b0000_0000;					inform_R [481][0] <= 8'b0000_0000;					inform_R [482][0] <= 8'b0000_0000;					inform_R [483][0] <= 8'b0000_0000;					inform_R [484][0] <= 8'b0000_0000;					inform_R [485][0] <= 8'b0000_0000;					inform_R [486][0] <= 8'b0000_0000;					inform_R [487][0] <= 8'b0000_0000;					inform_R [488][0] <= 8'b0000_0000;					inform_R [489][0] <= 8'b0000_0000;					inform_R [490][0] <= 8'b0000_0000;					inform_R [491][0] <= 8'b0000_0000;					inform_R [492][0] <= 8'b0000_0000;					inform_R [493][0] <= 8'b0000_0000;					inform_R [494][0] <= 8'b0000_0000;					inform_R [495][0] <= 8'b0000_0000;					inform_R [496][0] <= 8'b0000_0000;					inform_R [497][0] <= 8'b0000_0000;					inform_R [498][0] <= 8'b0000_0000;					inform_R [499][0] <= 8'b0000_0000;					inform_R [500][0] <= 8'b0000_0000;					inform_R [501][0] <= 8'b0000_0000;					inform_R [502][0] <= 8'b0000_0000;					inform_R [503][0] <= 8'b0000_0000;					inform_R [504][0] <= 8'b0000_0000;					inform_R [505][0] <= 8'b0000_0000;					inform_R [506][0] <= 8'b0000_0000;					inform_R [507][0] <= 8'b0000_0000;					inform_R [508][0] <= 8'b0000_0000;					inform_R [509][0] <= 8'b0000_0000;					inform_R [510][0] <= 8'b0000_0000;					inform_R [511][0] <= 8'b0000_0000;					inform_R [512][0] <= 8'b0111_1111;					inform_R [513][0] <= 8'b0111_1111;					inform_R [514][0] <= 8'b0111_1111;					inform_R [515][0] <= 8'b0111_1111;					inform_R [516][0] <= 8'b0111_1111;					inform_R [517][0] <= 8'b0111_1111;					inform_R [518][0] <= 8'b0111_1111;					inform_R [519][0] <= 8'b0111_1111;					inform_R [520][0] <= 8'b0111_1111;					inform_R [521][0] <= 8'b0111_1111;					inform_R [522][0] <= 8'b0111_1111;					inform_R [523][0] <= 8'b0111_1111;					inform_R [524][0] <= 8'b0111_1111;					inform_R [525][0] <= 8'b0111_1111;					inform_R [526][0] <= 8'b0111_1111;					inform_R [527][0] <= 8'b0000_0000;					inform_R [528][0] <= 8'b0111_1111;					inform_R [529][0] <= 8'b0111_1111;					inform_R [530][0] <= 8'b0111_1111;					inform_R [531][0] <= 8'b0111_1111;					inform_R [532][0] <= 8'b0111_1111;					inform_R [533][0] <= 8'b0111_1111;					inform_R [534][0] <= 8'b0111_1111;					inform_R [535][0] <= 8'b0000_0000;					inform_R [536][0] <= 8'b0111_1111;					inform_R [537][0] <= 8'b0111_1111;					inform_R [538][0] <= 8'b0111_1111;					inform_R [539][0] <= 8'b0000_0000;					inform_R [540][0] <= 8'b0111_1111;					inform_R [541][0] <= 8'b0000_0000;					inform_R [542][0] <= 8'b0000_0000;					inform_R [543][0] <= 8'b0000_0000;					inform_R [544][0] <= 8'b0111_1111;					inform_R [545][0] <= 8'b0111_1111;					inform_R [546][0] <= 8'b0111_1111;					inform_R [547][0] <= 8'b0111_1111;					inform_R [548][0] <= 8'b0111_1111;					inform_R [549][0] <= 8'b0111_1111;					inform_R [550][0] <= 8'b0111_1111;					inform_R [551][0] <= 8'b0000_0000;					inform_R [552][0] <= 8'b0111_1111;					inform_R [553][0] <= 8'b0111_1111;					inform_R [554][0] <= 8'b0000_0000;					inform_R [555][0] <= 8'b0000_0000;					inform_R [556][0] <= 8'b0000_0000;					inform_R [557][0] <= 8'b0000_0000;					inform_R [558][0] <= 8'b0000_0000;					inform_R [559][0] <= 8'b0000_0000;					inform_R [560][0] <= 8'b0111_1111;					inform_R [561][0] <= 8'b0000_0000;					inform_R [562][0] <= 8'b0000_0000;					inform_R [563][0] <= 8'b0000_0000;					inform_R [564][0] <= 8'b0000_0000;					inform_R [565][0] <= 8'b0000_0000;					inform_R [566][0] <= 8'b0000_0000;					inform_R [567][0] <= 8'b0000_0000;					inform_R [568][0] <= 8'b0000_0000;					inform_R [569][0] <= 8'b0000_0000;					inform_R [570][0] <= 8'b0000_0000;					inform_R [571][0] <= 8'b0000_0000;					inform_R [572][0] <= 8'b0000_0000;					inform_R [573][0] <= 8'b0000_0000;					inform_R [574][0] <= 8'b0000_0000;					inform_R [575][0] <= 8'b0000_0000;					inform_R [576][0] <= 8'b0111_1111;					inform_R [577][0] <= 8'b0111_1111;					inform_R [578][0] <= 8'b0111_1111;					inform_R [579][0] <= 8'b0000_0000;					inform_R [580][0] <= 8'b0111_1111;					inform_R [581][0] <= 8'b0000_0000;					inform_R [582][0] <= 8'b0000_0000;					inform_R [583][0] <= 8'b0000_0000;					inform_R [584][0] <= 8'b0111_1111;					inform_R [585][0] <= 8'b0000_0000;					inform_R [586][0] <= 8'b0000_0000;					inform_R [587][0] <= 8'b0000_0000;					inform_R [588][0] <= 8'b0000_0000;					inform_R [589][0] <= 8'b0000_0000;					inform_R [590][0] <= 8'b0000_0000;					inform_R [591][0] <= 8'b0000_0000;					inform_R [592][0] <= 8'b0111_1111;					inform_R [593][0] <= 8'b0000_0000;					inform_R [594][0] <= 8'b0000_0000;					inform_R [595][0] <= 8'b0000_0000;					inform_R [596][0] <= 8'b0000_0000;					inform_R [597][0] <= 8'b0000_0000;					inform_R [598][0] <= 8'b0000_0000;					inform_R [599][0] <= 8'b0000_0000;					inform_R [600][0] <= 8'b0000_0000;					inform_R [601][0] <= 8'b0000_0000;					inform_R [602][0] <= 8'b0000_0000;					inform_R [603][0] <= 8'b0000_0000;					inform_R [604][0] <= 8'b0000_0000;					inform_R [605][0] <= 8'b0000_0000;					inform_R [606][0] <= 8'b0000_0000;					inform_R [607][0] <= 8'b0000_0000;					inform_R [608][0] <= 8'b0000_0000;					inform_R [609][0] <= 8'b0000_0000;					inform_R [610][0] <= 8'b0000_0000;					inform_R [611][0] <= 8'b0000_0000;					inform_R [612][0] <= 8'b0000_0000;					inform_R [613][0] <= 8'b0000_0000;					inform_R [614][0] <= 8'b0000_0000;					inform_R [615][0] <= 8'b0000_0000;					inform_R [616][0] <= 8'b0000_0000;					inform_R [617][0] <= 8'b0000_0000;					inform_R [618][0] <= 8'b0000_0000;					inform_R [619][0] <= 8'b0000_0000;					inform_R [620][0] <= 8'b0000_0000;					inform_R [621][0] <= 8'b0000_0000;					inform_R [622][0] <= 8'b0000_0000;					inform_R [623][0] <= 8'b0000_0000;					inform_R [624][0] <= 8'b0000_0000;					inform_R [625][0] <= 8'b0000_0000;					inform_R [626][0] <= 8'b0000_0000;					inform_R [627][0] <= 8'b0000_0000;					inform_R [628][0] <= 8'b0000_0000;					inform_R [629][0] <= 8'b0000_0000;					inform_R [630][0] <= 8'b0000_0000;					inform_R [631][0] <= 8'b0000_0000;					inform_R [632][0] <= 8'b0000_0000;					inform_R [633][0] <= 8'b0000_0000;					inform_R [634][0] <= 8'b0000_0000;					inform_R [635][0] <= 8'b0000_0000;					inform_R [636][0] <= 8'b0000_0000;					inform_R [637][0] <= 8'b0000_0000;					inform_R [638][0] <= 8'b0000_0000;					inform_R [639][0] <= 8'b0000_0000;					inform_R [640][0] <= 8'b0111_1111;					inform_R [641][0] <= 8'b0111_1111;					inform_R [642][0] <= 8'b0111_1111;					inform_R [643][0] <= 8'b0000_0000;					inform_R [644][0] <= 8'b0111_1111;					inform_R [645][0] <= 8'b0000_0000;					inform_R [646][0] <= 8'b0000_0000;					inform_R [647][0] <= 8'b0000_0000;					inform_R [648][0] <= 8'b0000_0000;					inform_R [649][0] <= 8'b0000_0000;					inform_R [650][0] <= 8'b0000_0000;					inform_R [651][0] <= 8'b0000_0000;					inform_R [652][0] <= 8'b0000_0000;					inform_R [653][0] <= 8'b0000_0000;					inform_R [654][0] <= 8'b0000_0000;					inform_R [655][0] <= 8'b0000_0000;					inform_R [656][0] <= 8'b0000_0000;					inform_R [657][0] <= 8'b0000_0000;					inform_R [658][0] <= 8'b0000_0000;					inform_R [659][0] <= 8'b0000_0000;					inform_R [660][0] <= 8'b0000_0000;					inform_R [661][0] <= 8'b0000_0000;					inform_R [662][0] <= 8'b0000_0000;					inform_R [663][0] <= 8'b0000_0000;					inform_R [664][0] <= 8'b0000_0000;					inform_R [665][0] <= 8'b0000_0000;					inform_R [666][0] <= 8'b0000_0000;					inform_R [667][0] <= 8'b0000_0000;					inform_R [668][0] <= 8'b0000_0000;					inform_R [669][0] <= 8'b0000_0000;					inform_R [670][0] <= 8'b0000_0000;					inform_R [671][0] <= 8'b0000_0000;					inform_R [672][0] <= 8'b0000_0000;					inform_R [673][0] <= 8'b0000_0000;					inform_R [674][0] <= 8'b0000_0000;					inform_R [675][0] <= 8'b0000_0000;					inform_R [676][0] <= 8'b0000_0000;					inform_R [677][0] <= 8'b0000_0000;					inform_R [678][0] <= 8'b0000_0000;					inform_R [679][0] <= 8'b0000_0000;					inform_R [680][0] <= 8'b0000_0000;					inform_R [681][0] <= 8'b0000_0000;					inform_R [682][0] <= 8'b0000_0000;					inform_R [683][0] <= 8'b0000_0000;					inform_R [684][0] <= 8'b0000_0000;					inform_R [685][0] <= 8'b0000_0000;					inform_R [686][0] <= 8'b0000_0000;					inform_R [687][0] <= 8'b0000_0000;					inform_R [688][0] <= 8'b0000_0000;					inform_R [689][0] <= 8'b0000_0000;					inform_R [690][0] <= 8'b0000_0000;					inform_R [691][0] <= 8'b0000_0000;					inform_R [692][0] <= 8'b0000_0000;					inform_R [693][0] <= 8'b0000_0000;					inform_R [694][0] <= 8'b0000_0000;					inform_R [695][0] <= 8'b0000_0000;					inform_R [696][0] <= 8'b0000_0000;					inform_R [697][0] <= 8'b0000_0000;					inform_R [698][0] <= 8'b0000_0000;					inform_R [699][0] <= 8'b0000_0000;					inform_R [700][0] <= 8'b0000_0000;					inform_R [701][0] <= 8'b0000_0000;					inform_R [702][0] <= 8'b0000_0000;					inform_R [703][0] <= 8'b0000_0000;					inform_R [704][0] <= 8'b0000_0000;					inform_R [705][0] <= 8'b0000_0000;					inform_R [706][0] <= 8'b0000_0000;					inform_R [707][0] <= 8'b0000_0000;					inform_R [708][0] <= 8'b0000_0000;					inform_R [709][0] <= 8'b0000_0000;					inform_R [710][0] <= 8'b0000_0000;					inform_R [711][0] <= 8'b0000_0000;					inform_R [712][0] <= 8'b0000_0000;					inform_R [713][0] <= 8'b0000_0000;					inform_R [714][0] <= 8'b0000_0000;					inform_R [715][0] <= 8'b0000_0000;					inform_R [716][0] <= 8'b0000_0000;					inform_R [717][0] <= 8'b0000_0000;					inform_R [718][0] <= 8'b0000_0000;					inform_R [719][0] <= 8'b0000_0000;					inform_R [720][0] <= 8'b0000_0000;					inform_R [721][0] <= 8'b0000_0000;					inform_R [722][0] <= 8'b0000_0000;					inform_R [723][0] <= 8'b0000_0000;					inform_R [724][0] <= 8'b0000_0000;					inform_R [725][0] <= 8'b0000_0000;					inform_R [726][0] <= 8'b0000_0000;					inform_R [727][0] <= 8'b0000_0000;					inform_R [728][0] <= 8'b0000_0000;					inform_R [729][0] <= 8'b0000_0000;					inform_R [730][0] <= 8'b0000_0000;					inform_R [731][0] <= 8'b0000_0000;					inform_R [732][0] <= 8'b0000_0000;					inform_R [733][0] <= 8'b0000_0000;					inform_R [734][0] <= 8'b0000_0000;					inform_R [735][0] <= 8'b0000_0000;					inform_R [736][0] <= 8'b0000_0000;					inform_R [737][0] <= 8'b0000_0000;					inform_R [738][0] <= 8'b0000_0000;					inform_R [739][0] <= 8'b0000_0000;					inform_R [740][0] <= 8'b0000_0000;					inform_R [741][0] <= 8'b0000_0000;					inform_R [742][0] <= 8'b0000_0000;					inform_R [743][0] <= 8'b0000_0000;					inform_R [744][0] <= 8'b0000_0000;					inform_R [745][0] <= 8'b0000_0000;					inform_R [746][0] <= 8'b0000_0000;					inform_R [747][0] <= 8'b0000_0000;					inform_R [748][0] <= 8'b0000_0000;					inform_R [749][0] <= 8'b0000_0000;					inform_R [750][0] <= 8'b0000_0000;					inform_R [751][0] <= 8'b0000_0000;					inform_R [752][0] <= 8'b0000_0000;					inform_R [753][0] <= 8'b0000_0000;					inform_R [754][0] <= 8'b0000_0000;					inform_R [755][0] <= 8'b0000_0000;					inform_R [756][0] <= 8'b0000_0000;					inform_R [757][0] <= 8'b0000_0000;					inform_R [758][0] <= 8'b0000_0000;					inform_R [759][0] <= 8'b0000_0000;					inform_R [760][0] <= 8'b0000_0000;					inform_R [761][0] <= 8'b0000_0000;					inform_R [762][0] <= 8'b0000_0000;					inform_R [763][0] <= 8'b0000_0000;					inform_R [764][0] <= 8'b0000_0000;					inform_R [765][0] <= 8'b0000_0000;					inform_R [766][0] <= 8'b0000_0000;					inform_R [767][0] <= 8'b0000_0000;					inform_R [768][0] <= 8'b0111_1111;					inform_R [769][0] <= 8'b0000_0000;					inform_R [770][0] <= 8'b0000_0000;					inform_R [771][0] <= 8'b0000_0000;					inform_R [772][0] <= 8'b0000_0000;					inform_R [773][0] <= 8'b0000_0000;					inform_R [774][0] <= 8'b0000_0000;					inform_R [775][0] <= 8'b0000_0000;					inform_R [776][0] <= 8'b0000_0000;					inform_R [777][0] <= 8'b0000_0000;					inform_R [778][0] <= 8'b0000_0000;					inform_R [779][0] <= 8'b0000_0000;					inform_R [780][0] <= 8'b0000_0000;					inform_R [781][0] <= 8'b0000_0000;					inform_R [782][0] <= 8'b0000_0000;					inform_R [783][0] <= 8'b0000_0000;					inform_R [784][0] <= 8'b0000_0000;					inform_R [785][0] <= 8'b0000_0000;					inform_R [786][0] <= 8'b0000_0000;					inform_R [787][0] <= 8'b0000_0000;					inform_R [788][0] <= 8'b0000_0000;					inform_R [789][0] <= 8'b0000_0000;					inform_R [790][0] <= 8'b0000_0000;					inform_R [791][0] <= 8'b0000_0000;					inform_R [792][0] <= 8'b0000_0000;					inform_R [793][0] <= 8'b0000_0000;					inform_R [794][0] <= 8'b0000_0000;					inform_R [795][0] <= 8'b0000_0000;					inform_R [796][0] <= 8'b0000_0000;					inform_R [797][0] <= 8'b0000_0000;					inform_R [798][0] <= 8'b0000_0000;					inform_R [799][0] <= 8'b0000_0000;					inform_R [800][0] <= 8'b0000_0000;					inform_R [801][0] <= 8'b0000_0000;					inform_R [802][0] <= 8'b0000_0000;					inform_R [803][0] <= 8'b0000_0000;					inform_R [804][0] <= 8'b0000_0000;					inform_R [805][0] <= 8'b0000_0000;					inform_R [806][0] <= 8'b0000_0000;					inform_R [807][0] <= 8'b0000_0000;					inform_R [808][0] <= 8'b0000_0000;					inform_R [809][0] <= 8'b0000_0000;					inform_R [810][0] <= 8'b0000_0000;					inform_R [811][0] <= 8'b0000_0000;					inform_R [812][0] <= 8'b0000_0000;					inform_R [813][0] <= 8'b0000_0000;					inform_R [814][0] <= 8'b0000_0000;					inform_R [815][0] <= 8'b0000_0000;					inform_R [816][0] <= 8'b0000_0000;					inform_R [817][0] <= 8'b0000_0000;					inform_R [818][0] <= 8'b0000_0000;					inform_R [819][0] <= 8'b0000_0000;					inform_R [820][0] <= 8'b0000_0000;					inform_R [821][0] <= 8'b0000_0000;					inform_R [822][0] <= 8'b0000_0000;					inform_R [823][0] <= 8'b0000_0000;					inform_R [824][0] <= 8'b0000_0000;					inform_R [825][0] <= 8'b0000_0000;					inform_R [826][0] <= 8'b0000_0000;					inform_R [827][0] <= 8'b0000_0000;					inform_R [828][0] <= 8'b0000_0000;					inform_R [829][0] <= 8'b0000_0000;					inform_R [830][0] <= 8'b0000_0000;					inform_R [831][0] <= 8'b0000_0000;					inform_R [832][0] <= 8'b0000_0000;					inform_R [833][0] <= 8'b0000_0000;					inform_R [834][0] <= 8'b0000_0000;					inform_R [835][0] <= 8'b0000_0000;					inform_R [836][0] <= 8'b0000_0000;					inform_R [837][0] <= 8'b0000_0000;					inform_R [838][0] <= 8'b0000_0000;					inform_R [839][0] <= 8'b0000_0000;					inform_R [840][0] <= 8'b0000_0000;					inform_R [841][0] <= 8'b0000_0000;					inform_R [842][0] <= 8'b0000_0000;					inform_R [843][0] <= 8'b0000_0000;					inform_R [844][0] <= 8'b0000_0000;					inform_R [845][0] <= 8'b0000_0000;					inform_R [846][0] <= 8'b0000_0000;					inform_R [847][0] <= 8'b0000_0000;					inform_R [848][0] <= 8'b0000_0000;					inform_R [849][0] <= 8'b0000_0000;					inform_R [850][0] <= 8'b0000_0000;					inform_R [851][0] <= 8'b0000_0000;					inform_R [852][0] <= 8'b0000_0000;					inform_R [853][0] <= 8'b0000_0000;					inform_R [854][0] <= 8'b0000_0000;					inform_R [855][0] <= 8'b0000_0000;					inform_R [856][0] <= 8'b0000_0000;					inform_R [857][0] <= 8'b0000_0000;					inform_R [858][0] <= 8'b0000_0000;					inform_R [859][0] <= 8'b0000_0000;					inform_R [860][0] <= 8'b0000_0000;					inform_R [861][0] <= 8'b0000_0000;					inform_R [862][0] <= 8'b0000_0000;					inform_R [863][0] <= 8'b0000_0000;					inform_R [864][0] <= 8'b0000_0000;					inform_R [865][0] <= 8'b0000_0000;					inform_R [866][0] <= 8'b0000_0000;					inform_R [867][0] <= 8'b0000_0000;					inform_R [868][0] <= 8'b0000_0000;					inform_R [869][0] <= 8'b0000_0000;					inform_R [870][0] <= 8'b0000_0000;					inform_R [871][0] <= 8'b0000_0000;					inform_R [872][0] <= 8'b0000_0000;					inform_R [873][0] <= 8'b0000_0000;					inform_R [874][0] <= 8'b0000_0000;					inform_R [875][0] <= 8'b0000_0000;					inform_R [876][0] <= 8'b0000_0000;					inform_R [877][0] <= 8'b0000_0000;					inform_R [878][0] <= 8'b0000_0000;					inform_R [879][0] <= 8'b0000_0000;					inform_R [880][0] <= 8'b0000_0000;					inform_R [881][0] <= 8'b0000_0000;					inform_R [882][0] <= 8'b0000_0000;					inform_R [883][0] <= 8'b0000_0000;					inform_R [884][0] <= 8'b0000_0000;					inform_R [885][0] <= 8'b0000_0000;					inform_R [886][0] <= 8'b0000_0000;					inform_R [887][0] <= 8'b0000_0000;					inform_R [888][0] <= 8'b0000_0000;					inform_R [889][0] <= 8'b0000_0000;					inform_R [890][0] <= 8'b0000_0000;					inform_R [891][0] <= 8'b0000_0000;					inform_R [892][0] <= 8'b0000_0000;					inform_R [893][0] <= 8'b0000_0000;					inform_R [894][0] <= 8'b0000_0000;					inform_R [895][0] <= 8'b0000_0000;					inform_R [896][0] <= 8'b0000_0000;					inform_R [897][0] <= 8'b0000_0000;					inform_R [898][0] <= 8'b0000_0000;					inform_R [899][0] <= 8'b0000_0000;					inform_R [900][0] <= 8'b0000_0000;					inform_R [901][0] <= 8'b0000_0000;					inform_R [902][0] <= 8'b0000_0000;					inform_R [903][0] <= 8'b0000_0000;					inform_R [904][0] <= 8'b0000_0000;					inform_R [905][0] <= 8'b0000_0000;					inform_R [906][0] <= 8'b0000_0000;					inform_R [907][0] <= 8'b0000_0000;					inform_R [908][0] <= 8'b0000_0000;					inform_R [909][0] <= 8'b0000_0000;					inform_R [910][0] <= 8'b0000_0000;					inform_R [911][0] <= 8'b0000_0000;					inform_R [912][0] <= 8'b0000_0000;					inform_R [913][0] <= 8'b0000_0000;					inform_R [914][0] <= 8'b0000_0000;					inform_R [915][0] <= 8'b0000_0000;					inform_R [916][0] <= 8'b0000_0000;					inform_R [917][0] <= 8'b0000_0000;					inform_R [918][0] <= 8'b0000_0000;					inform_R [919][0] <= 8'b0000_0000;					inform_R [920][0] <= 8'b0000_0000;					inform_R [921][0] <= 8'b0000_0000;					inform_R [922][0] <= 8'b0000_0000;					inform_R [923][0] <= 8'b0000_0000;					inform_R [924][0] <= 8'b0000_0000;					inform_R [925][0] <= 8'b0000_0000;					inform_R [926][0] <= 8'b0000_0000;					inform_R [927][0] <= 8'b0000_0000;					inform_R [928][0] <= 8'b0000_0000;					inform_R [929][0] <= 8'b0000_0000;					inform_R [930][0] <= 8'b0000_0000;					inform_R [931][0] <= 8'b0000_0000;					inform_R [932][0] <= 8'b0000_0000;					inform_R [933][0] <= 8'b0000_0000;					inform_R [934][0] <= 8'b0000_0000;					inform_R [935][0] <= 8'b0000_0000;					inform_R [936][0] <= 8'b0000_0000;					inform_R [937][0] <= 8'b0000_0000;					inform_R [938][0] <= 8'b0000_0000;					inform_R [939][0] <= 8'b0000_0000;					inform_R [940][0] <= 8'b0000_0000;					inform_R [941][0] <= 8'b0000_0000;					inform_R [942][0] <= 8'b0000_0000;					inform_R [943][0] <= 8'b0000_0000;					inform_R [944][0] <= 8'b0000_0000;					inform_R [945][0] <= 8'b0000_0000;					inform_R [946][0] <= 8'b0000_0000;					inform_R [947][0] <= 8'b0000_0000;					inform_R [948][0] <= 8'b0000_0000;					inform_R [949][0] <= 8'b0000_0000;					inform_R [950][0] <= 8'b0000_0000;					inform_R [951][0] <= 8'b0000_0000;					inform_R [952][0] <= 8'b0000_0000;					inform_R [953][0] <= 8'b0000_0000;					inform_R [954][0] <= 8'b0000_0000;					inform_R [955][0] <= 8'b0000_0000;					inform_R [956][0] <= 8'b0000_0000;					inform_R [957][0] <= 8'b0000_0000;					inform_R [958][0] <= 8'b0000_0000;					inform_R [959][0] <= 8'b0000_0000;					inform_R [960][0] <= 8'b0000_0000;					inform_R [961][0] <= 8'b0000_0000;					inform_R [962][0] <= 8'b0000_0000;					inform_R [963][0] <= 8'b0000_0000;					inform_R [964][0] <= 8'b0000_0000;					inform_R [965][0] <= 8'b0000_0000;					inform_R [966][0] <= 8'b0000_0000;					inform_R [967][0] <= 8'b0000_0000;					inform_R [968][0] <= 8'b0000_0000;					inform_R [969][0] <= 8'b0000_0000;					inform_R [970][0] <= 8'b0000_0000;					inform_R [971][0] <= 8'b0000_0000;					inform_R [972][0] <= 8'b0000_0000;					inform_R [973][0] <= 8'b0000_0000;					inform_R [974][0] <= 8'b0000_0000;					inform_R [975][0] <= 8'b0000_0000;					inform_R [976][0] <= 8'b0000_0000;					inform_R [977][0] <= 8'b0000_0000;					inform_R [978][0] <= 8'b0000_0000;					inform_R [979][0] <= 8'b0000_0000;					inform_R [980][0] <= 8'b0000_0000;					inform_R [981][0] <= 8'b0000_0000;					inform_R [982][0] <= 8'b0000_0000;					inform_R [983][0] <= 8'b0000_0000;					inform_R [984][0] <= 8'b0000_0000;					inform_R [985][0] <= 8'b0000_0000;					inform_R [986][0] <= 8'b0000_0000;					inform_R [987][0] <= 8'b0000_0000;					inform_R [988][0] <= 8'b0000_0000;					inform_R [989][0] <= 8'b0000_0000;					inform_R [990][0] <= 8'b0000_0000;					inform_R [991][0] <= 8'b0000_0000;					inform_R [992][0] <= 8'b0000_0000;					inform_R [993][0] <= 8'b0000_0000;					inform_R [994][0] <= 8'b0000_0000;					inform_R [995][0] <= 8'b0000_0000;					inform_R [996][0] <= 8'b0000_0000;					inform_R [997][0] <= 8'b0000_0000;					inform_R [998][0] <= 8'b0000_0000;					inform_R [999][0] <= 8'b0000_0000;					inform_R [1000][0] <= 8'b0000_0000;					inform_R [1001][0] <= 8'b0000_0000;					inform_R [1002][0] <= 8'b0000_0000;					inform_R [1003][0] <= 8'b0000_0000;					inform_R [1004][0] <= 8'b0000_0000;					inform_R [1005][0] <= 8'b0000_0000;					inform_R [1006][0] <= 8'b0000_0000;					inform_R [1007][0] <= 8'b0000_0000;					inform_R [1008][0] <= 8'b0000_0000;					inform_R [1009][0] <= 8'b0000_0000;					inform_R [1010][0] <= 8'b0000_0000;					inform_R [1011][0] <= 8'b0000_0000;					inform_R [1012][0] <= 8'b0000_0000;					inform_R [1013][0] <= 8'b0000_0000;					inform_R [1014][0] <= 8'b0000_0000;					inform_R [1015][0] <= 8'b0000_0000;					inform_R [1016][0] <= 8'b0000_0000;					inform_R [1017][0] <= 8'b0000_0000;					inform_R [1018][0] <= 8'b0000_0000;					inform_R [1019][0] <= 8'b0000_0000;					inform_R [1020][0] <= 8'b0000_0000;					inform_R [1021][0] <= 8'b0000_0000;					inform_R [1022][0] <= 8'b0000_0000;					inform_R [1023][0] <= 8'b0000_0000;					inform_L [0][10] <= LLR_1;					inform_L [1][10] <= LLR_2;					inform_L [2][10] <= LLR_3;					inform_L [3][10] <= LLR_4;					inform_L [4][10] <= LLR_5;					inform_L [5][10] <= LLR_6;					inform_L [6][10] <= LLR_7;					inform_L [7][10] <= LLR_8;					inform_L [8][10] <= LLR_9;					inform_L [9][10] <= LLR_10;					inform_L [10][10] <= LLR_11;					inform_L [11][10] <= LLR_12;					inform_L [12][10] <= LLR_13;					inform_L [13][10] <= LLR_14;					inform_L [14][10] <= LLR_15;					inform_L [15][10] <= LLR_16;					inform_L [16][10] <= LLR_17;					inform_L [17][10] <= LLR_18;					inform_L [18][10] <= LLR_19;					inform_L [19][10] <= LLR_20;					inform_L [20][10] <= LLR_21;					inform_L [21][10] <= LLR_22;					inform_L [22][10] <= LLR_23;					inform_L [23][10] <= LLR_24;					inform_L [24][10] <= LLR_25;					inform_L [25][10] <= LLR_26;					inform_L [26][10] <= LLR_27;					inform_L [27][10] <= LLR_28;					inform_L [28][10] <= LLR_29;					inform_L [29][10] <= LLR_30;					inform_L [30][10] <= LLR_31;					inform_L [31][10] <= LLR_32;					inform_L [32][10] <= LLR_33;					inform_L [33][10] <= LLR_34;					inform_L [34][10] <= LLR_35;					inform_L [35][10] <= LLR_36;					inform_L [36][10] <= LLR_37;					inform_L [37][10] <= LLR_38;					inform_L [38][10] <= LLR_39;					inform_L [39][10] <= LLR_40;					inform_L [40][10] <= LLR_41;					inform_L [41][10] <= LLR_42;					inform_L [42][10] <= LLR_43;					inform_L [43][10] <= LLR_44;					inform_L [44][10] <= LLR_45;					inform_L [45][10] <= LLR_46;					inform_L [46][10] <= LLR_47;					inform_L [47][10] <= LLR_48;					inform_L [48][10] <= LLR_49;					inform_L [49][10] <= LLR_50;					inform_L [50][10] <= LLR_51;					inform_L [51][10] <= LLR_52;					inform_L [52][10] <= LLR_53;					inform_L [53][10] <= LLR_54;					inform_L [54][10] <= LLR_55;					inform_L [55][10] <= LLR_56;					inform_L [56][10] <= LLR_57;					inform_L [57][10] <= LLR_58;					inform_L [58][10] <= LLR_59;					inform_L [59][10] <= LLR_60;					inform_L [60][10] <= LLR_61;					inform_L [61][10] <= LLR_62;					inform_L [62][10] <= LLR_63;					inform_L [63][10] <= LLR_64;					inform_L [64][10] <= LLR_65;					inform_L [65][10] <= LLR_66;					inform_L [66][10] <= LLR_67;					inform_L [67][10] <= LLR_68;					inform_L [68][10] <= LLR_69;					inform_L [69][10] <= LLR_70;					inform_L [70][10] <= LLR_71;					inform_L [71][10] <= LLR_72;					inform_L [72][10] <= LLR_73;					inform_L [73][10] <= LLR_74;					inform_L [74][10] <= LLR_75;					inform_L [75][10] <= LLR_76;					inform_L [76][10] <= LLR_77;					inform_L [77][10] <= LLR_78;					inform_L [78][10] <= LLR_79;					inform_L [79][10] <= LLR_80;					inform_L [80][10] <= LLR_81;					inform_L [81][10] <= LLR_82;					inform_L [82][10] <= LLR_83;					inform_L [83][10] <= LLR_84;					inform_L [84][10] <= LLR_85;					inform_L [85][10] <= LLR_86;					inform_L [86][10] <= LLR_87;					inform_L [87][10] <= LLR_88;					inform_L [88][10] <= LLR_89;					inform_L [89][10] <= LLR_90;					inform_L [90][10] <= LLR_91;					inform_L [91][10] <= LLR_92;					inform_L [92][10] <= LLR_93;					inform_L [93][10] <= LLR_94;					inform_L [94][10] <= LLR_95;					inform_L [95][10] <= LLR_96;					inform_L [96][10] <= LLR_97;					inform_L [97][10] <= LLR_98;					inform_L [98][10] <= LLR_99;					inform_L [99][10] <= LLR_100;					inform_L [100][10] <= LLR_101;					inform_L [101][10] <= LLR_102;					inform_L [102][10] <= LLR_103;					inform_L [103][10] <= LLR_104;					inform_L [104][10] <= LLR_105;					inform_L [105][10] <= LLR_106;					inform_L [106][10] <= LLR_107;					inform_L [107][10] <= LLR_108;					inform_L [108][10] <= LLR_109;					inform_L [109][10] <= LLR_110;					inform_L [110][10] <= LLR_111;					inform_L [111][10] <= LLR_112;					inform_L [112][10] <= LLR_113;					inform_L [113][10] <= LLR_114;					inform_L [114][10] <= LLR_115;					inform_L [115][10] <= LLR_116;					inform_L [116][10] <= LLR_117;					inform_L [117][10] <= LLR_118;					inform_L [118][10] <= LLR_119;					inform_L [119][10] <= LLR_120;					inform_L [120][10] <= LLR_121;					inform_L [121][10] <= LLR_122;					inform_L [122][10] <= LLR_123;					inform_L [123][10] <= LLR_124;					inform_L [124][10] <= LLR_125;					inform_L [125][10] <= LLR_126;					inform_L [126][10] <= LLR_127;					inform_L [127][10] <= LLR_128;					inform_L [128][10] <= LLR_129;					inform_L [129][10] <= LLR_130;					inform_L [130][10] <= LLR_131;					inform_L [131][10] <= LLR_132;					inform_L [132][10] <= LLR_133;					inform_L [133][10] <= LLR_134;					inform_L [134][10] <= LLR_135;					inform_L [135][10] <= LLR_136;					inform_L [136][10] <= LLR_137;					inform_L [137][10] <= LLR_138;					inform_L [138][10] <= LLR_139;					inform_L [139][10] <= LLR_140;					inform_L [140][10] <= LLR_141;					inform_L [141][10] <= LLR_142;					inform_L [142][10] <= LLR_143;					inform_L [143][10] <= LLR_144;					inform_L [144][10] <= LLR_145;					inform_L [145][10] <= LLR_146;					inform_L [146][10] <= LLR_147;					inform_L [147][10] <= LLR_148;					inform_L [148][10] <= LLR_149;					inform_L [149][10] <= LLR_150;					inform_L [150][10] <= LLR_151;					inform_L [151][10] <= LLR_152;					inform_L [152][10] <= LLR_153;					inform_L [153][10] <= LLR_154;					inform_L [154][10] <= LLR_155;					inform_L [155][10] <= LLR_156;					inform_L [156][10] <= LLR_157;					inform_L [157][10] <= LLR_158;					inform_L [158][10] <= LLR_159;					inform_L [159][10] <= LLR_160;					inform_L [160][10] <= LLR_161;					inform_L [161][10] <= LLR_162;					inform_L [162][10] <= LLR_163;					inform_L [163][10] <= LLR_164;					inform_L [164][10] <= LLR_165;					inform_L [165][10] <= LLR_166;					inform_L [166][10] <= LLR_167;					inform_L [167][10] <= LLR_168;					inform_L [168][10] <= LLR_169;					inform_L [169][10] <= LLR_170;					inform_L [170][10] <= LLR_171;					inform_L [171][10] <= LLR_172;					inform_L [172][10] <= LLR_173;					inform_L [173][10] <= LLR_174;					inform_L [174][10] <= LLR_175;					inform_L [175][10] <= LLR_176;					inform_L [176][10] <= LLR_177;					inform_L [177][10] <= LLR_178;					inform_L [178][10] <= LLR_179;					inform_L [179][10] <= LLR_180;					inform_L [180][10] <= LLR_181;					inform_L [181][10] <= LLR_182;					inform_L [182][10] <= LLR_183;					inform_L [183][10] <= LLR_184;					inform_L [184][10] <= LLR_185;					inform_L [185][10] <= LLR_186;					inform_L [186][10] <= LLR_187;					inform_L [187][10] <= LLR_188;					inform_L [188][10] <= LLR_189;					inform_L [189][10] <= LLR_190;					inform_L [190][10] <= LLR_191;					inform_L [191][10] <= LLR_192;					inform_L [192][10] <= LLR_193;					inform_L [193][10] <= LLR_194;					inform_L [194][10] <= LLR_195;					inform_L [195][10] <= LLR_196;					inform_L [196][10] <= LLR_197;					inform_L [197][10] <= LLR_198;					inform_L [198][10] <= LLR_199;					inform_L [199][10] <= LLR_200;					inform_L [200][10] <= LLR_201;					inform_L [201][10] <= LLR_202;					inform_L [202][10] <= LLR_203;					inform_L [203][10] <= LLR_204;					inform_L [204][10] <= LLR_205;					inform_L [205][10] <= LLR_206;					inform_L [206][10] <= LLR_207;					inform_L [207][10] <= LLR_208;					inform_L [208][10] <= LLR_209;					inform_L [209][10] <= LLR_210;					inform_L [210][10] <= LLR_211;					inform_L [211][10] <= LLR_212;					inform_L [212][10] <= LLR_213;					inform_L [213][10] <= LLR_214;					inform_L [214][10] <= LLR_215;					inform_L [215][10] <= LLR_216;					inform_L [216][10] <= LLR_217;					inform_L [217][10] <= LLR_218;					inform_L [218][10] <= LLR_219;					inform_L [219][10] <= LLR_220;					inform_L [220][10] <= LLR_221;					inform_L [221][10] <= LLR_222;					inform_L [222][10] <= LLR_223;					inform_L [223][10] <= LLR_224;					inform_L [224][10] <= LLR_225;					inform_L [225][10] <= LLR_226;					inform_L [226][10] <= LLR_227;					inform_L [227][10] <= LLR_228;					inform_L [228][10] <= LLR_229;					inform_L [229][10] <= LLR_230;					inform_L [230][10] <= LLR_231;					inform_L [231][10] <= LLR_232;					inform_L [232][10] <= LLR_233;					inform_L [233][10] <= LLR_234;					inform_L [234][10] <= LLR_235;					inform_L [235][10] <= LLR_236;					inform_L [236][10] <= LLR_237;					inform_L [237][10] <= LLR_238;					inform_L [238][10] <= LLR_239;					inform_L [239][10] <= LLR_240;					inform_L [240][10] <= LLR_241;					inform_L [241][10] <= LLR_242;					inform_L [242][10] <= LLR_243;					inform_L [243][10] <= LLR_244;					inform_L [244][10] <= LLR_245;					inform_L [245][10] <= LLR_246;					inform_L [246][10] <= LLR_247;					inform_L [247][10] <= LLR_248;					inform_L [248][10] <= LLR_249;					inform_L [249][10] <= LLR_250;					inform_L [250][10] <= LLR_251;					inform_L [251][10] <= LLR_252;					inform_L [252][10] <= LLR_253;					inform_L [253][10] <= LLR_254;					inform_L [254][10] <= LLR_255;					inform_L [255][10] <= LLR_256;					inform_L [256][10] <= LLR_257;					inform_L [257][10] <= LLR_258;					inform_L [258][10] <= LLR_259;					inform_L [259][10] <= LLR_260;					inform_L [260][10] <= LLR_261;					inform_L [261][10] <= LLR_262;					inform_L [262][10] <= LLR_263;					inform_L [263][10] <= LLR_264;					inform_L [264][10] <= LLR_265;					inform_L [265][10] <= LLR_266;					inform_L [266][10] <= LLR_267;					inform_L [267][10] <= LLR_268;					inform_L [268][10] <= LLR_269;					inform_L [269][10] <= LLR_270;					inform_L [270][10] <= LLR_271;					inform_L [271][10] <= LLR_272;					inform_L [272][10] <= LLR_273;					inform_L [273][10] <= LLR_274;					inform_L [274][10] <= LLR_275;					inform_L [275][10] <= LLR_276;					inform_L [276][10] <= LLR_277;					inform_L [277][10] <= LLR_278;					inform_L [278][10] <= LLR_279;					inform_L [279][10] <= LLR_280;					inform_L [280][10] <= LLR_281;					inform_L [281][10] <= LLR_282;					inform_L [282][10] <= LLR_283;					inform_L [283][10] <= LLR_284;					inform_L [284][10] <= LLR_285;					inform_L [285][10] <= LLR_286;					inform_L [286][10] <= LLR_287;					inform_L [287][10] <= LLR_288;					inform_L [288][10] <= LLR_289;					inform_L [289][10] <= LLR_290;					inform_L [290][10] <= LLR_291;					inform_L [291][10] <= LLR_292;					inform_L [292][10] <= LLR_293;					inform_L [293][10] <= LLR_294;					inform_L [294][10] <= LLR_295;					inform_L [295][10] <= LLR_296;					inform_L [296][10] <= LLR_297;					inform_L [297][10] <= LLR_298;					inform_L [298][10] <= LLR_299;					inform_L [299][10] <= LLR_300;					inform_L [300][10] <= LLR_301;					inform_L [301][10] <= LLR_302;					inform_L [302][10] <= LLR_303;					inform_L [303][10] <= LLR_304;					inform_L [304][10] <= LLR_305;					inform_L [305][10] <= LLR_306;					inform_L [306][10] <= LLR_307;					inform_L [307][10] <= LLR_308;					inform_L [308][10] <= LLR_309;					inform_L [309][10] <= LLR_310;					inform_L [310][10] <= LLR_311;					inform_L [311][10] <= LLR_312;					inform_L [312][10] <= LLR_313;					inform_L [313][10] <= LLR_314;					inform_L [314][10] <= LLR_315;					inform_L [315][10] <= LLR_316;					inform_L [316][10] <= LLR_317;					inform_L [317][10] <= LLR_318;					inform_L [318][10] <= LLR_319;					inform_L [319][10] <= LLR_320;					inform_L [320][10] <= LLR_321;					inform_L [321][10] <= LLR_322;					inform_L [322][10] <= LLR_323;					inform_L [323][10] <= LLR_324;					inform_L [324][10] <= LLR_325;					inform_L [325][10] <= LLR_326;					inform_L [326][10] <= LLR_327;					inform_L [327][10] <= LLR_328;					inform_L [328][10] <= LLR_329;					inform_L [329][10] <= LLR_330;					inform_L [330][10] <= LLR_331;					inform_L [331][10] <= LLR_332;					inform_L [332][10] <= LLR_333;					inform_L [333][10] <= LLR_334;					inform_L [334][10] <= LLR_335;					inform_L [335][10] <= LLR_336;					inform_L [336][10] <= LLR_337;					inform_L [337][10] <= LLR_338;					inform_L [338][10] <= LLR_339;					inform_L [339][10] <= LLR_340;					inform_L [340][10] <= LLR_341;					inform_L [341][10] <= LLR_342;					inform_L [342][10] <= LLR_343;					inform_L [343][10] <= LLR_344;					inform_L [344][10] <= LLR_345;					inform_L [345][10] <= LLR_346;					inform_L [346][10] <= LLR_347;					inform_L [347][10] <= LLR_348;					inform_L [348][10] <= LLR_349;					inform_L [349][10] <= LLR_350;					inform_L [350][10] <= LLR_351;					inform_L [351][10] <= LLR_352;					inform_L [352][10] <= LLR_353;					inform_L [353][10] <= LLR_354;					inform_L [354][10] <= LLR_355;					inform_L [355][10] <= LLR_356;					inform_L [356][10] <= LLR_357;					inform_L [357][10] <= LLR_358;					inform_L [358][10] <= LLR_359;					inform_L [359][10] <= LLR_360;					inform_L [360][10] <= LLR_361;					inform_L [361][10] <= LLR_362;					inform_L [362][10] <= LLR_363;					inform_L [363][10] <= LLR_364;					inform_L [364][10] <= LLR_365;					inform_L [365][10] <= LLR_366;					inform_L [366][10] <= LLR_367;					inform_L [367][10] <= LLR_368;					inform_L [368][10] <= LLR_369;					inform_L [369][10] <= LLR_370;					inform_L [370][10] <= LLR_371;					inform_L [371][10] <= LLR_372;					inform_L [372][10] <= LLR_373;					inform_L [373][10] <= LLR_374;					inform_L [374][10] <= LLR_375;					inform_L [375][10] <= LLR_376;					inform_L [376][10] <= LLR_377;					inform_L [377][10] <= LLR_378;					inform_L [378][10] <= LLR_379;					inform_L [379][10] <= LLR_380;					inform_L [380][10] <= LLR_381;					inform_L [381][10] <= LLR_382;					inform_L [382][10] <= LLR_383;					inform_L [383][10] <= LLR_384;					inform_L [384][10] <= LLR_385;					inform_L [385][10] <= LLR_386;					inform_L [386][10] <= LLR_387;					inform_L [387][10] <= LLR_388;					inform_L [388][10] <= LLR_389;					inform_L [389][10] <= LLR_390;					inform_L [390][10] <= LLR_391;					inform_L [391][10] <= LLR_392;					inform_L [392][10] <= LLR_393;					inform_L [393][10] <= LLR_394;					inform_L [394][10] <= LLR_395;					inform_L [395][10] <= LLR_396;					inform_L [396][10] <= LLR_397;					inform_L [397][10] <= LLR_398;					inform_L [398][10] <= LLR_399;					inform_L [399][10] <= LLR_400;					inform_L [400][10] <= LLR_401;					inform_L [401][10] <= LLR_402;					inform_L [402][10] <= LLR_403;					inform_L [403][10] <= LLR_404;					inform_L [404][10] <= LLR_405;					inform_L [405][10] <= LLR_406;					inform_L [406][10] <= LLR_407;					inform_L [407][10] <= LLR_408;					inform_L [408][10] <= LLR_409;					inform_L [409][10] <= LLR_410;					inform_L [410][10] <= LLR_411;					inform_L [411][10] <= LLR_412;					inform_L [412][10] <= LLR_413;					inform_L [413][10] <= LLR_414;					inform_L [414][10] <= LLR_415;					inform_L [415][10] <= LLR_416;					inform_L [416][10] <= LLR_417;					inform_L [417][10] <= LLR_418;					inform_L [418][10] <= LLR_419;					inform_L [419][10] <= LLR_420;					inform_L [420][10] <= LLR_421;					inform_L [421][10] <= LLR_422;					inform_L [422][10] <= LLR_423;					inform_L [423][10] <= LLR_424;					inform_L [424][10] <= LLR_425;					inform_L [425][10] <= LLR_426;					inform_L [426][10] <= LLR_427;					inform_L [427][10] <= LLR_428;					inform_L [428][10] <= LLR_429;					inform_L [429][10] <= LLR_430;					inform_L [430][10] <= LLR_431;					inform_L [431][10] <= LLR_432;					inform_L [432][10] <= LLR_433;					inform_L [433][10] <= LLR_434;					inform_L [434][10] <= LLR_435;					inform_L [435][10] <= LLR_436;					inform_L [436][10] <= LLR_437;					inform_L [437][10] <= LLR_438;					inform_L [438][10] <= LLR_439;					inform_L [439][10] <= LLR_440;					inform_L [440][10] <= LLR_441;					inform_L [441][10] <= LLR_442;					inform_L [442][10] <= LLR_443;					inform_L [443][10] <= LLR_444;					inform_L [444][10] <= LLR_445;					inform_L [445][10] <= LLR_446;					inform_L [446][10] <= LLR_447;					inform_L [447][10] <= LLR_448;					inform_L [448][10] <= LLR_449;					inform_L [449][10] <= LLR_450;					inform_L [450][10] <= LLR_451;					inform_L [451][10] <= LLR_452;					inform_L [452][10] <= LLR_453;					inform_L [453][10] <= LLR_454;					inform_L [454][10] <= LLR_455;					inform_L [455][10] <= LLR_456;					inform_L [456][10] <= LLR_457;					inform_L [457][10] <= LLR_458;					inform_L [458][10] <= LLR_459;					inform_L [459][10] <= LLR_460;					inform_L [460][10] <= LLR_461;					inform_L [461][10] <= LLR_462;					inform_L [462][10] <= LLR_463;					inform_L [463][10] <= LLR_464;					inform_L [464][10] <= LLR_465;					inform_L [465][10] <= LLR_466;					inform_L [466][10] <= LLR_467;					inform_L [467][10] <= LLR_468;					inform_L [468][10] <= LLR_469;					inform_L [469][10] <= LLR_470;					inform_L [470][10] <= LLR_471;					inform_L [471][10] <= LLR_472;					inform_L [472][10] <= LLR_473;					inform_L [473][10] <= LLR_474;					inform_L [474][10] <= LLR_475;					inform_L [475][10] <= LLR_476;					inform_L [476][10] <= LLR_477;					inform_L [477][10] <= LLR_478;					inform_L [478][10] <= LLR_479;					inform_L [479][10] <= LLR_480;					inform_L [480][10] <= LLR_481;					inform_L [481][10] <= LLR_482;					inform_L [482][10] <= LLR_483;					inform_L [483][10] <= LLR_484;					inform_L [484][10] <= LLR_485;					inform_L [485][10] <= LLR_486;					inform_L [486][10] <= LLR_487;					inform_L [487][10] <= LLR_488;					inform_L [488][10] <= LLR_489;					inform_L [489][10] <= LLR_490;					inform_L [490][10] <= LLR_491;					inform_L [491][10] <= LLR_492;					inform_L [492][10] <= LLR_493;					inform_L [493][10] <= LLR_494;					inform_L [494][10] <= LLR_495;					inform_L [495][10] <= LLR_496;					inform_L [496][10] <= LLR_497;					inform_L [497][10] <= LLR_498;					inform_L [498][10] <= LLR_499;					inform_L [499][10] <= LLR_500;					inform_L [500][10] <= LLR_501;					inform_L [501][10] <= LLR_502;					inform_L [502][10] <= LLR_503;					inform_L [503][10] <= LLR_504;					inform_L [504][10] <= LLR_505;					inform_L [505][10] <= LLR_506;					inform_L [506][10] <= LLR_507;					inform_L [507][10] <= LLR_508;					inform_L [508][10] <= LLR_509;					inform_L [509][10] <= LLR_510;					inform_L [510][10] <= LLR_511;					inform_L [511][10] <= LLR_512;					inform_L [512][10] <= LLR_513;					inform_L [513][10] <= LLR_514;					inform_L [514][10] <= LLR_515;					inform_L [515][10] <= LLR_516;					inform_L [516][10] <= LLR_517;					inform_L [517][10] <= LLR_518;					inform_L [518][10] <= LLR_519;					inform_L [519][10] <= LLR_520;					inform_L [520][10] <= LLR_521;					inform_L [521][10] <= LLR_522;					inform_L [522][10] <= LLR_523;					inform_L [523][10] <= LLR_524;					inform_L [524][10] <= LLR_525;					inform_L [525][10] <= LLR_526;					inform_L [526][10] <= LLR_527;					inform_L [527][10] <= LLR_528;					inform_L [528][10] <= LLR_529;					inform_L [529][10] <= LLR_530;					inform_L [530][10] <= LLR_531;					inform_L [531][10] <= LLR_532;					inform_L [532][10] <= LLR_533;					inform_L [533][10] <= LLR_534;					inform_L [534][10] <= LLR_535;					inform_L [535][10] <= LLR_536;					inform_L [536][10] <= LLR_537;					inform_L [537][10] <= LLR_538;					inform_L [538][10] <= LLR_539;					inform_L [539][10] <= LLR_540;					inform_L [540][10] <= LLR_541;					inform_L [541][10] <= LLR_542;					inform_L [542][10] <= LLR_543;					inform_L [543][10] <= LLR_544;					inform_L [544][10] <= LLR_545;					inform_L [545][10] <= LLR_546;					inform_L [546][10] <= LLR_547;					inform_L [547][10] <= LLR_548;					inform_L [548][10] <= LLR_549;					inform_L [549][10] <= LLR_550;					inform_L [550][10] <= LLR_551;					inform_L [551][10] <= LLR_552;					inform_L [552][10] <= LLR_553;					inform_L [553][10] <= LLR_554;					inform_L [554][10] <= LLR_555;					inform_L [555][10] <= LLR_556;					inform_L [556][10] <= LLR_557;					inform_L [557][10] <= LLR_558;					inform_L [558][10] <= LLR_559;					inform_L [559][10] <= LLR_560;					inform_L [560][10] <= LLR_561;					inform_L [561][10] <= LLR_562;					inform_L [562][10] <= LLR_563;					inform_L [563][10] <= LLR_564;					inform_L [564][10] <= LLR_565;					inform_L [565][10] <= LLR_566;					inform_L [566][10] <= LLR_567;					inform_L [567][10] <= LLR_568;					inform_L [568][10] <= LLR_569;					inform_L [569][10] <= LLR_570;					inform_L [570][10] <= LLR_571;					inform_L [571][10] <= LLR_572;					inform_L [572][10] <= LLR_573;					inform_L [573][10] <= LLR_574;					inform_L [574][10] <= LLR_575;					inform_L [575][10] <= LLR_576;					inform_L [576][10] <= LLR_577;					inform_L [577][10] <= LLR_578;					inform_L [578][10] <= LLR_579;					inform_L [579][10] <= LLR_580;					inform_L [580][10] <= LLR_581;					inform_L [581][10] <= LLR_582;					inform_L [582][10] <= LLR_583;					inform_L [583][10] <= LLR_584;					inform_L [584][10] <= LLR_585;					inform_L [585][10] <= LLR_586;					inform_L [586][10] <= LLR_587;					inform_L [587][10] <= LLR_588;					inform_L [588][10] <= LLR_589;					inform_L [589][10] <= LLR_590;					inform_L [590][10] <= LLR_591;					inform_L [591][10] <= LLR_592;					inform_L [592][10] <= LLR_593;					inform_L [593][10] <= LLR_594;					inform_L [594][10] <= LLR_595;					inform_L [595][10] <= LLR_596;					inform_L [596][10] <= LLR_597;					inform_L [597][10] <= LLR_598;					inform_L [598][10] <= LLR_599;					inform_L [599][10] <= LLR_600;					inform_L [600][10] <= LLR_601;					inform_L [601][10] <= LLR_602;					inform_L [602][10] <= LLR_603;					inform_L [603][10] <= LLR_604;					inform_L [604][10] <= LLR_605;					inform_L [605][10] <= LLR_606;					inform_L [606][10] <= LLR_607;					inform_L [607][10] <= LLR_608;					inform_L [608][10] <= LLR_609;					inform_L [609][10] <= LLR_610;					inform_L [610][10] <= LLR_611;					inform_L [611][10] <= LLR_612;					inform_L [612][10] <= LLR_613;					inform_L [613][10] <= LLR_614;					inform_L [614][10] <= LLR_615;					inform_L [615][10] <= LLR_616;					inform_L [616][10] <= LLR_617;					inform_L [617][10] <= LLR_618;					inform_L [618][10] <= LLR_619;					inform_L [619][10] <= LLR_620;					inform_L [620][10] <= LLR_621;					inform_L [621][10] <= LLR_622;					inform_L [622][10] <= LLR_623;					inform_L [623][10] <= LLR_624;					inform_L [624][10] <= LLR_625;					inform_L [625][10] <= LLR_626;					inform_L [626][10] <= LLR_627;					inform_L [627][10] <= LLR_628;					inform_L [628][10] <= LLR_629;					inform_L [629][10] <= LLR_630;					inform_L [630][10] <= LLR_631;					inform_L [631][10] <= LLR_632;					inform_L [632][10] <= LLR_633;					inform_L [633][10] <= LLR_634;					inform_L [634][10] <= LLR_635;					inform_L [635][10] <= LLR_636;					inform_L [636][10] <= LLR_637;					inform_L [637][10] <= LLR_638;					inform_L [638][10] <= LLR_639;					inform_L [639][10] <= LLR_640;					inform_L [640][10] <= LLR_641;					inform_L [641][10] <= LLR_642;					inform_L [642][10] <= LLR_643;					inform_L [643][10] <= LLR_644;					inform_L [644][10] <= LLR_645;					inform_L [645][10] <= LLR_646;					inform_L [646][10] <= LLR_647;					inform_L [647][10] <= LLR_648;					inform_L [648][10] <= LLR_649;					inform_L [649][10] <= LLR_650;					inform_L [650][10] <= LLR_651;					inform_L [651][10] <= LLR_652;					inform_L [652][10] <= LLR_653;					inform_L [653][10] <= LLR_654;					inform_L [654][10] <= LLR_655;					inform_L [655][10] <= LLR_656;					inform_L [656][10] <= LLR_657;					inform_L [657][10] <= LLR_658;					inform_L [658][10] <= LLR_659;					inform_L [659][10] <= LLR_660;					inform_L [660][10] <= LLR_661;					inform_L [661][10] <= LLR_662;					inform_L [662][10] <= LLR_663;					inform_L [663][10] <= LLR_664;					inform_L [664][10] <= LLR_665;					inform_L [665][10] <= LLR_666;					inform_L [666][10] <= LLR_667;					inform_L [667][10] <= LLR_668;					inform_L [668][10] <= LLR_669;					inform_L [669][10] <= LLR_670;					inform_L [670][10] <= LLR_671;					inform_L [671][10] <= LLR_672;					inform_L [672][10] <= LLR_673;					inform_L [673][10] <= LLR_674;					inform_L [674][10] <= LLR_675;					inform_L [675][10] <= LLR_676;					inform_L [676][10] <= LLR_677;					inform_L [677][10] <= LLR_678;					inform_L [678][10] <= LLR_679;					inform_L [679][10] <= LLR_680;					inform_L [680][10] <= LLR_681;					inform_L [681][10] <= LLR_682;					inform_L [682][10] <= LLR_683;					inform_L [683][10] <= LLR_684;					inform_L [684][10] <= LLR_685;					inform_L [685][10] <= LLR_686;					inform_L [686][10] <= LLR_687;					inform_L [687][10] <= LLR_688;					inform_L [688][10] <= LLR_689;					inform_L [689][10] <= LLR_690;					inform_L [690][10] <= LLR_691;					inform_L [691][10] <= LLR_692;					inform_L [692][10] <= LLR_693;					inform_L [693][10] <= LLR_694;					inform_L [694][10] <= LLR_695;					inform_L [695][10] <= LLR_696;					inform_L [696][10] <= LLR_697;					inform_L [697][10] <= LLR_698;					inform_L [698][10] <= LLR_699;					inform_L [699][10] <= LLR_700;					inform_L [700][10] <= LLR_701;					inform_L [701][10] <= LLR_702;					inform_L [702][10] <= LLR_703;					inform_L [703][10] <= LLR_704;					inform_L [704][10] <= LLR_705;					inform_L [705][10] <= LLR_706;					inform_L [706][10] <= LLR_707;					inform_L [707][10] <= LLR_708;					inform_L [708][10] <= LLR_709;					inform_L [709][10] <= LLR_710;					inform_L [710][10] <= LLR_711;					inform_L [711][10] <= LLR_712;					inform_L [712][10] <= LLR_713;					inform_L [713][10] <= LLR_714;					inform_L [714][10] <= LLR_715;					inform_L [715][10] <= LLR_716;					inform_L [716][10] <= LLR_717;					inform_L [717][10] <= LLR_718;					inform_L [718][10] <= LLR_719;					inform_L [719][10] <= LLR_720;					inform_L [720][10] <= LLR_721;					inform_L [721][10] <= LLR_722;					inform_L [722][10] <= LLR_723;					inform_L [723][10] <= LLR_724;					inform_L [724][10] <= LLR_725;					inform_L [725][10] <= LLR_726;					inform_L [726][10] <= LLR_727;					inform_L [727][10] <= LLR_728;					inform_L [728][10] <= LLR_729;					inform_L [729][10] <= LLR_730;					inform_L [730][10] <= LLR_731;					inform_L [731][10] <= LLR_732;					inform_L [732][10] <= LLR_733;					inform_L [733][10] <= LLR_734;					inform_L [734][10] <= LLR_735;					inform_L [735][10] <= LLR_736;					inform_L [736][10] <= LLR_737;					inform_L [737][10] <= LLR_738;					inform_L [738][10] <= LLR_739;					inform_L [739][10] <= LLR_740;					inform_L [740][10] <= LLR_741;					inform_L [741][10] <= LLR_742;					inform_L [742][10] <= LLR_743;					inform_L [743][10] <= LLR_744;					inform_L [744][10] <= LLR_745;					inform_L [745][10] <= LLR_746;					inform_L [746][10] <= LLR_747;					inform_L [747][10] <= LLR_748;					inform_L [748][10] <= LLR_749;					inform_L [749][10] <= LLR_750;					inform_L [750][10] <= LLR_751;					inform_L [751][10] <= LLR_752;					inform_L [752][10] <= LLR_753;					inform_L [753][10] <= LLR_754;					inform_L [754][10] <= LLR_755;					inform_L [755][10] <= LLR_756;					inform_L [756][10] <= LLR_757;					inform_L [757][10] <= LLR_758;					inform_L [758][10] <= LLR_759;					inform_L [759][10] <= LLR_760;					inform_L [760][10] <= LLR_761;					inform_L [761][10] <= LLR_762;					inform_L [762][10] <= LLR_763;					inform_L [763][10] <= LLR_764;					inform_L [764][10] <= LLR_765;					inform_L [765][10] <= LLR_766;					inform_L [766][10] <= LLR_767;					inform_L [767][10] <= LLR_768;					inform_L [768][10] <= LLR_769;					inform_L [769][10] <= LLR_770;					inform_L [770][10] <= LLR_771;					inform_L [771][10] <= LLR_772;					inform_L [772][10] <= LLR_773;					inform_L [773][10] <= LLR_774;					inform_L [774][10] <= LLR_775;					inform_L [775][10] <= LLR_776;					inform_L [776][10] <= LLR_777;					inform_L [777][10] <= LLR_778;					inform_L [778][10] <= LLR_779;					inform_L [779][10] <= LLR_780;					inform_L [780][10] <= LLR_781;					inform_L [781][10] <= LLR_782;					inform_L [782][10] <= LLR_783;					inform_L [783][10] <= LLR_784;					inform_L [784][10] <= LLR_785;					inform_L [785][10] <= LLR_786;					inform_L [786][10] <= LLR_787;					inform_L [787][10] <= LLR_788;					inform_L [788][10] <= LLR_789;					inform_L [789][10] <= LLR_790;					inform_L [790][10] <= LLR_791;					inform_L [791][10] <= LLR_792;					inform_L [792][10] <= LLR_793;					inform_L [793][10] <= LLR_794;					inform_L [794][10] <= LLR_795;					inform_L [795][10] <= LLR_796;					inform_L [796][10] <= LLR_797;					inform_L [797][10] <= LLR_798;					inform_L [798][10] <= LLR_799;					inform_L [799][10] <= LLR_800;					inform_L [800][10] <= LLR_801;					inform_L [801][10] <= LLR_802;					inform_L [802][10] <= LLR_803;					inform_L [803][10] <= LLR_804;					inform_L [804][10] <= LLR_805;					inform_L [805][10] <= LLR_806;					inform_L [806][10] <= LLR_807;					inform_L [807][10] <= LLR_808;					inform_L [808][10] <= LLR_809;					inform_L [809][10] <= LLR_810;					inform_L [810][10] <= LLR_811;					inform_L [811][10] <= LLR_812;					inform_L [812][10] <= LLR_813;					inform_L [813][10] <= LLR_814;					inform_L [814][10] <= LLR_815;					inform_L [815][10] <= LLR_816;					inform_L [816][10] <= LLR_817;					inform_L [817][10] <= LLR_818;					inform_L [818][10] <= LLR_819;					inform_L [819][10] <= LLR_820;					inform_L [820][10] <= LLR_821;					inform_L [821][10] <= LLR_822;					inform_L [822][10] <= LLR_823;					inform_L [823][10] <= LLR_824;					inform_L [824][10] <= LLR_825;					inform_L [825][10] <= LLR_826;					inform_L [826][10] <= LLR_827;					inform_L [827][10] <= LLR_828;					inform_L [828][10] <= LLR_829;					inform_L [829][10] <= LLR_830;					inform_L [830][10] <= LLR_831;					inform_L [831][10] <= LLR_832;					inform_L [832][10] <= LLR_833;					inform_L [833][10] <= LLR_834;					inform_L [834][10] <= LLR_835;					inform_L [835][10] <= LLR_836;					inform_L [836][10] <= LLR_837;					inform_L [837][10] <= LLR_838;					inform_L [838][10] <= LLR_839;					inform_L [839][10] <= LLR_840;					inform_L [840][10] <= LLR_841;					inform_L [841][10] <= LLR_842;					inform_L [842][10] <= LLR_843;					inform_L [843][10] <= LLR_844;					inform_L [844][10] <= LLR_845;					inform_L [845][10] <= LLR_846;					inform_L [846][10] <= LLR_847;					inform_L [847][10] <= LLR_848;					inform_L [848][10] <= LLR_849;					inform_L [849][10] <= LLR_850;					inform_L [850][10] <= LLR_851;					inform_L [851][10] <= LLR_852;					inform_L [852][10] <= LLR_853;					inform_L [853][10] <= LLR_854;					inform_L [854][10] <= LLR_855;					inform_L [855][10] <= LLR_856;					inform_L [856][10] <= LLR_857;					inform_L [857][10] <= LLR_858;					inform_L [858][10] <= LLR_859;					inform_L [859][10] <= LLR_860;					inform_L [860][10] <= LLR_861;					inform_L [861][10] <= LLR_862;					inform_L [862][10] <= LLR_863;					inform_L [863][10] <= LLR_864;					inform_L [864][10] <= LLR_865;					inform_L [865][10] <= LLR_866;					inform_L [866][10] <= LLR_867;					inform_L [867][10] <= LLR_868;					inform_L [868][10] <= LLR_869;					inform_L [869][10] <= LLR_870;					inform_L [870][10] <= LLR_871;					inform_L [871][10] <= LLR_872;					inform_L [872][10] <= LLR_873;					inform_L [873][10] <= LLR_874;					inform_L [874][10] <= LLR_875;					inform_L [875][10] <= LLR_876;					inform_L [876][10] <= LLR_877;					inform_L [877][10] <= LLR_878;					inform_L [878][10] <= LLR_879;					inform_L [879][10] <= LLR_880;					inform_L [880][10] <= LLR_881;					inform_L [881][10] <= LLR_882;					inform_L [882][10] <= LLR_883;					inform_L [883][10] <= LLR_884;					inform_L [884][10] <= LLR_885;					inform_L [885][10] <= LLR_886;					inform_L [886][10] <= LLR_887;					inform_L [887][10] <= LLR_888;					inform_L [888][10] <= LLR_889;					inform_L [889][10] <= LLR_890;					inform_L [890][10] <= LLR_891;					inform_L [891][10] <= LLR_892;					inform_L [892][10] <= LLR_893;					inform_L [893][10] <= LLR_894;					inform_L [894][10] <= LLR_895;					inform_L [895][10] <= LLR_896;					inform_L [896][10] <= LLR_897;					inform_L [897][10] <= LLR_898;					inform_L [898][10] <= LLR_899;					inform_L [899][10] <= LLR_900;					inform_L [900][10] <= LLR_901;					inform_L [901][10] <= LLR_902;					inform_L [902][10] <= LLR_903;					inform_L [903][10] <= LLR_904;					inform_L [904][10] <= LLR_905;					inform_L [905][10] <= LLR_906;					inform_L [906][10] <= LLR_907;					inform_L [907][10] <= LLR_908;					inform_L [908][10] <= LLR_909;					inform_L [909][10] <= LLR_910;					inform_L [910][10] <= LLR_911;					inform_L [911][10] <= LLR_912;					inform_L [912][10] <= LLR_913;					inform_L [913][10] <= LLR_914;					inform_L [914][10] <= LLR_915;					inform_L [915][10] <= LLR_916;					inform_L [916][10] <= LLR_917;					inform_L [917][10] <= LLR_918;					inform_L [918][10] <= LLR_919;					inform_L [919][10] <= LLR_920;					inform_L [920][10] <= LLR_921;					inform_L [921][10] <= LLR_922;					inform_L [922][10] <= LLR_923;					inform_L [923][10] <= LLR_924;					inform_L [924][10] <= LLR_925;					inform_L [925][10] <= LLR_926;					inform_L [926][10] <= LLR_927;					inform_L [927][10] <= LLR_928;					inform_L [928][10] <= LLR_929;					inform_L [929][10] <= LLR_930;					inform_L [930][10] <= LLR_931;					inform_L [931][10] <= LLR_932;					inform_L [932][10] <= LLR_933;					inform_L [933][10] <= LLR_934;					inform_L [934][10] <= LLR_935;					inform_L [935][10] <= LLR_936;					inform_L [936][10] <= LLR_937;					inform_L [937][10] <= LLR_938;					inform_L [938][10] <= LLR_939;					inform_L [939][10] <= LLR_940;					inform_L [940][10] <= LLR_941;					inform_L [941][10] <= LLR_942;					inform_L [942][10] <= LLR_943;					inform_L [943][10] <= LLR_944;					inform_L [944][10] <= LLR_945;					inform_L [945][10] <= LLR_946;					inform_L [946][10] <= LLR_947;					inform_L [947][10] <= LLR_948;					inform_L [948][10] <= LLR_949;					inform_L [949][10] <= LLR_950;					inform_L [950][10] <= LLR_951;					inform_L [951][10] <= LLR_952;					inform_L [952][10] <= LLR_953;					inform_L [953][10] <= LLR_954;					inform_L [954][10] <= LLR_955;					inform_L [955][10] <= LLR_956;					inform_L [956][10] <= LLR_957;					inform_L [957][10] <= LLR_958;					inform_L [958][10] <= LLR_959;					inform_L [959][10] <= LLR_960;					inform_L [960][10] <= LLR_961;					inform_L [961][10] <= LLR_962;					inform_L [962][10] <= LLR_963;					inform_L [963][10] <= LLR_964;					inform_L [964][10] <= LLR_965;					inform_L [965][10] <= LLR_966;					inform_L [966][10] <= LLR_967;					inform_L [967][10] <= LLR_968;					inform_L [968][10] <= LLR_969;					inform_L [969][10] <= LLR_970;					inform_L [970][10] <= LLR_971;					inform_L [971][10] <= LLR_972;					inform_L [972][10] <= LLR_973;					inform_L [973][10] <= LLR_974;					inform_L [974][10] <= LLR_975;					inform_L [975][10] <= LLR_976;					inform_L [976][10] <= LLR_977;					inform_L [977][10] <= LLR_978;					inform_L [978][10] <= LLR_979;					inform_L [979][10] <= LLR_980;					inform_L [980][10] <= LLR_981;					inform_L [981][10] <= LLR_982;					inform_L [982][10] <= LLR_983;					inform_L [983][10] <= LLR_984;					inform_L [984][10] <= LLR_985;					inform_L [985][10] <= LLR_986;					inform_L [986][10] <= LLR_987;					inform_L [987][10] <= LLR_988;					inform_L [988][10] <= LLR_989;					inform_L [989][10] <= LLR_990;					inform_L [990][10] <= LLR_991;					inform_L [991][10] <= LLR_992;					inform_L [992][10] <= LLR_993;					inform_L [993][10] <= LLR_994;					inform_L [994][10] <= LLR_995;					inform_L [995][10] <= LLR_996;					inform_L [996][10] <= LLR_997;					inform_L [997][10] <= LLR_998;					inform_L [998][10] <= LLR_999;					inform_L [999][10] <= LLR_1000;					inform_L [1000][10] <= LLR_1001;					inform_L [1001][10] <= LLR_1002;					inform_L [1002][10] <= LLR_1003;					inform_L [1003][10] <= LLR_1004;					inform_L [1004][10] <= LLR_1005;					inform_L [1005][10] <= LLR_1006;					inform_L [1006][10] <= LLR_1007;					inform_L [1007][10] <= LLR_1008;					inform_L [1008][10] <= LLR_1009;					inform_L [1009][10] <= LLR_1010;					inform_L [1010][10] <= LLR_1011;					inform_L [1011][10] <= LLR_1012;					inform_L [1012][10] <= LLR_1013;					inform_L [1013][10] <= LLR_1014;					inform_L [1014][10] <= LLR_1015;					inform_L [1015][10] <= LLR_1016;					inform_L [1016][10] <= LLR_1017;					inform_L [1017][10] <= LLR_1018;					inform_L [1018][10] <= LLR_1019;					inform_L [1019][10] <= LLR_1020;					inform_L [1020][10] <= LLR_1021;					inform_L [1021][10] <= LLR_1022;					inform_L [1022][10] <= LLR_1023;					inform_L [1023][10] <= LLR_1024;				end				for (x = 0; x < 1024; x = x + 1)					for (y = 0; y < 10; y = y + 1)					begin						inform_R[x][y+1] <= 8'd0;						inform_L[x][y] <= 8'd0;					end			end
			BUSY_LEFT:			begin				if(clk_counter == 2'b11)begin					case (w2r)						1:						begin							inform_R[0][1] = r_cell_wire[0];							inform_R[1][1] = r_cell_wire[1];							inform_R[2][1] = r_cell_wire[2];							inform_R[3][1] = r_cell_wire[3];							inform_R[4][1] = r_cell_wire[4];							inform_R[5][1] = r_cell_wire[5];							inform_R[6][1] = r_cell_wire[6];							inform_R[7][1] = r_cell_wire[7];							inform_R[8][1] = r_cell_wire[8];							inform_R[9][1] = r_cell_wire[9];							inform_R[10][1] = r_cell_wire[10];							inform_R[11][1] = r_cell_wire[11];							inform_R[12][1] = r_cell_wire[12];							inform_R[13][1] = r_cell_wire[13];							inform_R[14][1] = r_cell_wire[14];							inform_R[15][1] = r_cell_wire[15];							inform_R[16][1] = r_cell_wire[16];							inform_R[17][1] = r_cell_wire[17];							inform_R[18][1] = r_cell_wire[18];							inform_R[19][1] = r_cell_wire[19];							inform_R[20][1] = r_cell_wire[20];							inform_R[21][1] = r_cell_wire[21];							inform_R[22][1] = r_cell_wire[22];							inform_R[23][1] = r_cell_wire[23];							inform_R[24][1] = r_cell_wire[24];							inform_R[25][1] = r_cell_wire[25];							inform_R[26][1] = r_cell_wire[26];							inform_R[27][1] = r_cell_wire[27];							inform_R[28][1] = r_cell_wire[28];							inform_R[29][1] = r_cell_wire[29];							inform_R[30][1] = r_cell_wire[30];							inform_R[31][1] = r_cell_wire[31];							inform_R[32][1] = r_cell_wire[32];							inform_R[33][1] = r_cell_wire[33];							inform_R[34][1] = r_cell_wire[34];							inform_R[35][1] = r_cell_wire[35];							inform_R[36][1] = r_cell_wire[36];							inform_R[37][1] = r_cell_wire[37];							inform_R[38][1] = r_cell_wire[38];							inform_R[39][1] = r_cell_wire[39];							inform_R[40][1] = r_cell_wire[40];							inform_R[41][1] = r_cell_wire[41];							inform_R[42][1] = r_cell_wire[42];							inform_R[43][1] = r_cell_wire[43];							inform_R[44][1] = r_cell_wire[44];							inform_R[45][1] = r_cell_wire[45];							inform_R[46][1] = r_cell_wire[46];							inform_R[47][1] = r_cell_wire[47];							inform_R[48][1] = r_cell_wire[48];							inform_R[49][1] = r_cell_wire[49];							inform_R[50][1] = r_cell_wire[50];							inform_R[51][1] = r_cell_wire[51];							inform_R[52][1] = r_cell_wire[52];							inform_R[53][1] = r_cell_wire[53];							inform_R[54][1] = r_cell_wire[54];							inform_R[55][1] = r_cell_wire[55];							inform_R[56][1] = r_cell_wire[56];							inform_R[57][1] = r_cell_wire[57];							inform_R[58][1] = r_cell_wire[58];							inform_R[59][1] = r_cell_wire[59];							inform_R[60][1] = r_cell_wire[60];							inform_R[61][1] = r_cell_wire[61];							inform_R[62][1] = r_cell_wire[62];							inform_R[63][1] = r_cell_wire[63];							inform_R[64][1] = r_cell_wire[64];							inform_R[65][1] = r_cell_wire[65];							inform_R[66][1] = r_cell_wire[66];							inform_R[67][1] = r_cell_wire[67];							inform_R[68][1] = r_cell_wire[68];							inform_R[69][1] = r_cell_wire[69];							inform_R[70][1] = r_cell_wire[70];							inform_R[71][1] = r_cell_wire[71];							inform_R[72][1] = r_cell_wire[72];							inform_R[73][1] = r_cell_wire[73];							inform_R[74][1] = r_cell_wire[74];							inform_R[75][1] = r_cell_wire[75];							inform_R[76][1] = r_cell_wire[76];							inform_R[77][1] = r_cell_wire[77];							inform_R[78][1] = r_cell_wire[78];							inform_R[79][1] = r_cell_wire[79];							inform_R[80][1] = r_cell_wire[80];							inform_R[81][1] = r_cell_wire[81];							inform_R[82][1] = r_cell_wire[82];							inform_R[83][1] = r_cell_wire[83];							inform_R[84][1] = r_cell_wire[84];							inform_R[85][1] = r_cell_wire[85];							inform_R[86][1] = r_cell_wire[86];							inform_R[87][1] = r_cell_wire[87];							inform_R[88][1] = r_cell_wire[88];							inform_R[89][1] = r_cell_wire[89];							inform_R[90][1] = r_cell_wire[90];							inform_R[91][1] = r_cell_wire[91];							inform_R[92][1] = r_cell_wire[92];							inform_R[93][1] = r_cell_wire[93];							inform_R[94][1] = r_cell_wire[94];							inform_R[95][1] = r_cell_wire[95];							inform_R[96][1] = r_cell_wire[96];							inform_R[97][1] = r_cell_wire[97];							inform_R[98][1] = r_cell_wire[98];							inform_R[99][1] = r_cell_wire[99];							inform_R[100][1] = r_cell_wire[100];							inform_R[101][1] = r_cell_wire[101];							inform_R[102][1] = r_cell_wire[102];							inform_R[103][1] = r_cell_wire[103];							inform_R[104][1] = r_cell_wire[104];							inform_R[105][1] = r_cell_wire[105];							inform_R[106][1] = r_cell_wire[106];							inform_R[107][1] = r_cell_wire[107];							inform_R[108][1] = r_cell_wire[108];							inform_R[109][1] = r_cell_wire[109];							inform_R[110][1] = r_cell_wire[110];							inform_R[111][1] = r_cell_wire[111];							inform_R[112][1] = r_cell_wire[112];							inform_R[113][1] = r_cell_wire[113];							inform_R[114][1] = r_cell_wire[114];							inform_R[115][1] = r_cell_wire[115];							inform_R[116][1] = r_cell_wire[116];							inform_R[117][1] = r_cell_wire[117];							inform_R[118][1] = r_cell_wire[118];							inform_R[119][1] = r_cell_wire[119];							inform_R[120][1] = r_cell_wire[120];							inform_R[121][1] = r_cell_wire[121];							inform_R[122][1] = r_cell_wire[122];							inform_R[123][1] = r_cell_wire[123];							inform_R[124][1] = r_cell_wire[124];							inform_R[125][1] = r_cell_wire[125];							inform_R[126][1] = r_cell_wire[126];							inform_R[127][1] = r_cell_wire[127];							inform_R[128][1] = r_cell_wire[128];							inform_R[129][1] = r_cell_wire[129];							inform_R[130][1] = r_cell_wire[130];							inform_R[131][1] = r_cell_wire[131];							inform_R[132][1] = r_cell_wire[132];							inform_R[133][1] = r_cell_wire[133];							inform_R[134][1] = r_cell_wire[134];							inform_R[135][1] = r_cell_wire[135];							inform_R[136][1] = r_cell_wire[136];							inform_R[137][1] = r_cell_wire[137];							inform_R[138][1] = r_cell_wire[138];							inform_R[139][1] = r_cell_wire[139];							inform_R[140][1] = r_cell_wire[140];							inform_R[141][1] = r_cell_wire[141];							inform_R[142][1] = r_cell_wire[142];							inform_R[143][1] = r_cell_wire[143];							inform_R[144][1] = r_cell_wire[144];							inform_R[145][1] = r_cell_wire[145];							inform_R[146][1] = r_cell_wire[146];							inform_R[147][1] = r_cell_wire[147];							inform_R[148][1] = r_cell_wire[148];							inform_R[149][1] = r_cell_wire[149];							inform_R[150][1] = r_cell_wire[150];							inform_R[151][1] = r_cell_wire[151];							inform_R[152][1] = r_cell_wire[152];							inform_R[153][1] = r_cell_wire[153];							inform_R[154][1] = r_cell_wire[154];							inform_R[155][1] = r_cell_wire[155];							inform_R[156][1] = r_cell_wire[156];							inform_R[157][1] = r_cell_wire[157];							inform_R[158][1] = r_cell_wire[158];							inform_R[159][1] = r_cell_wire[159];							inform_R[160][1] = r_cell_wire[160];							inform_R[161][1] = r_cell_wire[161];							inform_R[162][1] = r_cell_wire[162];							inform_R[163][1] = r_cell_wire[163];							inform_R[164][1] = r_cell_wire[164];							inform_R[165][1] = r_cell_wire[165];							inform_R[166][1] = r_cell_wire[166];							inform_R[167][1] = r_cell_wire[167];							inform_R[168][1] = r_cell_wire[168];							inform_R[169][1] = r_cell_wire[169];							inform_R[170][1] = r_cell_wire[170];							inform_R[171][1] = r_cell_wire[171];							inform_R[172][1] = r_cell_wire[172];							inform_R[173][1] = r_cell_wire[173];							inform_R[174][1] = r_cell_wire[174];							inform_R[175][1] = r_cell_wire[175];							inform_R[176][1] = r_cell_wire[176];							inform_R[177][1] = r_cell_wire[177];							inform_R[178][1] = r_cell_wire[178];							inform_R[179][1] = r_cell_wire[179];							inform_R[180][1] = r_cell_wire[180];							inform_R[181][1] = r_cell_wire[181];							inform_R[182][1] = r_cell_wire[182];							inform_R[183][1] = r_cell_wire[183];							inform_R[184][1] = r_cell_wire[184];							inform_R[185][1] = r_cell_wire[185];							inform_R[186][1] = r_cell_wire[186];							inform_R[187][1] = r_cell_wire[187];							inform_R[188][1] = r_cell_wire[188];							inform_R[189][1] = r_cell_wire[189];							inform_R[190][1] = r_cell_wire[190];							inform_R[191][1] = r_cell_wire[191];							inform_R[192][1] = r_cell_wire[192];							inform_R[193][1] = r_cell_wire[193];							inform_R[194][1] = r_cell_wire[194];							inform_R[195][1] = r_cell_wire[195];							inform_R[196][1] = r_cell_wire[196];							inform_R[197][1] = r_cell_wire[197];							inform_R[198][1] = r_cell_wire[198];							inform_R[199][1] = r_cell_wire[199];							inform_R[200][1] = r_cell_wire[200];							inform_R[201][1] = r_cell_wire[201];							inform_R[202][1] = r_cell_wire[202];							inform_R[203][1] = r_cell_wire[203];							inform_R[204][1] = r_cell_wire[204];							inform_R[205][1] = r_cell_wire[205];							inform_R[206][1] = r_cell_wire[206];							inform_R[207][1] = r_cell_wire[207];							inform_R[208][1] = r_cell_wire[208];							inform_R[209][1] = r_cell_wire[209];							inform_R[210][1] = r_cell_wire[210];							inform_R[211][1] = r_cell_wire[211];							inform_R[212][1] = r_cell_wire[212];							inform_R[213][1] = r_cell_wire[213];							inform_R[214][1] = r_cell_wire[214];							inform_R[215][1] = r_cell_wire[215];							inform_R[216][1] = r_cell_wire[216];							inform_R[217][1] = r_cell_wire[217];							inform_R[218][1] = r_cell_wire[218];							inform_R[219][1] = r_cell_wire[219];							inform_R[220][1] = r_cell_wire[220];							inform_R[221][1] = r_cell_wire[221];							inform_R[222][1] = r_cell_wire[222];							inform_R[223][1] = r_cell_wire[223];							inform_R[224][1] = r_cell_wire[224];							inform_R[225][1] = r_cell_wire[225];							inform_R[226][1] = r_cell_wire[226];							inform_R[227][1] = r_cell_wire[227];							inform_R[228][1] = r_cell_wire[228];							inform_R[229][1] = r_cell_wire[229];							inform_R[230][1] = r_cell_wire[230];							inform_R[231][1] = r_cell_wire[231];							inform_R[232][1] = r_cell_wire[232];							inform_R[233][1] = r_cell_wire[233];							inform_R[234][1] = r_cell_wire[234];							inform_R[235][1] = r_cell_wire[235];							inform_R[236][1] = r_cell_wire[236];							inform_R[237][1] = r_cell_wire[237];							inform_R[238][1] = r_cell_wire[238];							inform_R[239][1] = r_cell_wire[239];							inform_R[240][1] = r_cell_wire[240];							inform_R[241][1] = r_cell_wire[241];							inform_R[242][1] = r_cell_wire[242];							inform_R[243][1] = r_cell_wire[243];							inform_R[244][1] = r_cell_wire[244];							inform_R[245][1] = r_cell_wire[245];							inform_R[246][1] = r_cell_wire[246];							inform_R[247][1] = r_cell_wire[247];							inform_R[248][1] = r_cell_wire[248];							inform_R[249][1] = r_cell_wire[249];							inform_R[250][1] = r_cell_wire[250];							inform_R[251][1] = r_cell_wire[251];							inform_R[252][1] = r_cell_wire[252];							inform_R[253][1] = r_cell_wire[253];							inform_R[254][1] = r_cell_wire[254];							inform_R[255][1] = r_cell_wire[255];							inform_R[256][1] = r_cell_wire[256];							inform_R[257][1] = r_cell_wire[257];							inform_R[258][1] = r_cell_wire[258];							inform_R[259][1] = r_cell_wire[259];							inform_R[260][1] = r_cell_wire[260];							inform_R[261][1] = r_cell_wire[261];							inform_R[262][1] = r_cell_wire[262];							inform_R[263][1] = r_cell_wire[263];							inform_R[264][1] = r_cell_wire[264];							inform_R[265][1] = r_cell_wire[265];							inform_R[266][1] = r_cell_wire[266];							inform_R[267][1] = r_cell_wire[267];							inform_R[268][1] = r_cell_wire[268];							inform_R[269][1] = r_cell_wire[269];							inform_R[270][1] = r_cell_wire[270];							inform_R[271][1] = r_cell_wire[271];							inform_R[272][1] = r_cell_wire[272];							inform_R[273][1] = r_cell_wire[273];							inform_R[274][1] = r_cell_wire[274];							inform_R[275][1] = r_cell_wire[275];							inform_R[276][1] = r_cell_wire[276];							inform_R[277][1] = r_cell_wire[277];							inform_R[278][1] = r_cell_wire[278];							inform_R[279][1] = r_cell_wire[279];							inform_R[280][1] = r_cell_wire[280];							inform_R[281][1] = r_cell_wire[281];							inform_R[282][1] = r_cell_wire[282];							inform_R[283][1] = r_cell_wire[283];							inform_R[284][1] = r_cell_wire[284];							inform_R[285][1] = r_cell_wire[285];							inform_R[286][1] = r_cell_wire[286];							inform_R[287][1] = r_cell_wire[287];							inform_R[288][1] = r_cell_wire[288];							inform_R[289][1] = r_cell_wire[289];							inform_R[290][1] = r_cell_wire[290];							inform_R[291][1] = r_cell_wire[291];							inform_R[292][1] = r_cell_wire[292];							inform_R[293][1] = r_cell_wire[293];							inform_R[294][1] = r_cell_wire[294];							inform_R[295][1] = r_cell_wire[295];							inform_R[296][1] = r_cell_wire[296];							inform_R[297][1] = r_cell_wire[297];							inform_R[298][1] = r_cell_wire[298];							inform_R[299][1] = r_cell_wire[299];							inform_R[300][1] = r_cell_wire[300];							inform_R[301][1] = r_cell_wire[301];							inform_R[302][1] = r_cell_wire[302];							inform_R[303][1] = r_cell_wire[303];							inform_R[304][1] = r_cell_wire[304];							inform_R[305][1] = r_cell_wire[305];							inform_R[306][1] = r_cell_wire[306];							inform_R[307][1] = r_cell_wire[307];							inform_R[308][1] = r_cell_wire[308];							inform_R[309][1] = r_cell_wire[309];							inform_R[310][1] = r_cell_wire[310];							inform_R[311][1] = r_cell_wire[311];							inform_R[312][1] = r_cell_wire[312];							inform_R[313][1] = r_cell_wire[313];							inform_R[314][1] = r_cell_wire[314];							inform_R[315][1] = r_cell_wire[315];							inform_R[316][1] = r_cell_wire[316];							inform_R[317][1] = r_cell_wire[317];							inform_R[318][1] = r_cell_wire[318];							inform_R[319][1] = r_cell_wire[319];							inform_R[320][1] = r_cell_wire[320];							inform_R[321][1] = r_cell_wire[321];							inform_R[322][1] = r_cell_wire[322];							inform_R[323][1] = r_cell_wire[323];							inform_R[324][1] = r_cell_wire[324];							inform_R[325][1] = r_cell_wire[325];							inform_R[326][1] = r_cell_wire[326];							inform_R[327][1] = r_cell_wire[327];							inform_R[328][1] = r_cell_wire[328];							inform_R[329][1] = r_cell_wire[329];							inform_R[330][1] = r_cell_wire[330];							inform_R[331][1] = r_cell_wire[331];							inform_R[332][1] = r_cell_wire[332];							inform_R[333][1] = r_cell_wire[333];							inform_R[334][1] = r_cell_wire[334];							inform_R[335][1] = r_cell_wire[335];							inform_R[336][1] = r_cell_wire[336];							inform_R[337][1] = r_cell_wire[337];							inform_R[338][1] = r_cell_wire[338];							inform_R[339][1] = r_cell_wire[339];							inform_R[340][1] = r_cell_wire[340];							inform_R[341][1] = r_cell_wire[341];							inform_R[342][1] = r_cell_wire[342];							inform_R[343][1] = r_cell_wire[343];							inform_R[344][1] = r_cell_wire[344];							inform_R[345][1] = r_cell_wire[345];							inform_R[346][1] = r_cell_wire[346];							inform_R[347][1] = r_cell_wire[347];							inform_R[348][1] = r_cell_wire[348];							inform_R[349][1] = r_cell_wire[349];							inform_R[350][1] = r_cell_wire[350];							inform_R[351][1] = r_cell_wire[351];							inform_R[352][1] = r_cell_wire[352];							inform_R[353][1] = r_cell_wire[353];							inform_R[354][1] = r_cell_wire[354];							inform_R[355][1] = r_cell_wire[355];							inform_R[356][1] = r_cell_wire[356];							inform_R[357][1] = r_cell_wire[357];							inform_R[358][1] = r_cell_wire[358];							inform_R[359][1] = r_cell_wire[359];							inform_R[360][1] = r_cell_wire[360];							inform_R[361][1] = r_cell_wire[361];							inform_R[362][1] = r_cell_wire[362];							inform_R[363][1] = r_cell_wire[363];							inform_R[364][1] = r_cell_wire[364];							inform_R[365][1] = r_cell_wire[365];							inform_R[366][1] = r_cell_wire[366];							inform_R[367][1] = r_cell_wire[367];							inform_R[368][1] = r_cell_wire[368];							inform_R[369][1] = r_cell_wire[369];							inform_R[370][1] = r_cell_wire[370];							inform_R[371][1] = r_cell_wire[371];							inform_R[372][1] = r_cell_wire[372];							inform_R[373][1] = r_cell_wire[373];							inform_R[374][1] = r_cell_wire[374];							inform_R[375][1] = r_cell_wire[375];							inform_R[376][1] = r_cell_wire[376];							inform_R[377][1] = r_cell_wire[377];							inform_R[378][1] = r_cell_wire[378];							inform_R[379][1] = r_cell_wire[379];							inform_R[380][1] = r_cell_wire[380];							inform_R[381][1] = r_cell_wire[381];							inform_R[382][1] = r_cell_wire[382];							inform_R[383][1] = r_cell_wire[383];							inform_R[384][1] = r_cell_wire[384];							inform_R[385][1] = r_cell_wire[385];							inform_R[386][1] = r_cell_wire[386];							inform_R[387][1] = r_cell_wire[387];							inform_R[388][1] = r_cell_wire[388];							inform_R[389][1] = r_cell_wire[389];							inform_R[390][1] = r_cell_wire[390];							inform_R[391][1] = r_cell_wire[391];							inform_R[392][1] = r_cell_wire[392];							inform_R[393][1] = r_cell_wire[393];							inform_R[394][1] = r_cell_wire[394];							inform_R[395][1] = r_cell_wire[395];							inform_R[396][1] = r_cell_wire[396];							inform_R[397][1] = r_cell_wire[397];							inform_R[398][1] = r_cell_wire[398];							inform_R[399][1] = r_cell_wire[399];							inform_R[400][1] = r_cell_wire[400];							inform_R[401][1] = r_cell_wire[401];							inform_R[402][1] = r_cell_wire[402];							inform_R[403][1] = r_cell_wire[403];							inform_R[404][1] = r_cell_wire[404];							inform_R[405][1] = r_cell_wire[405];							inform_R[406][1] = r_cell_wire[406];							inform_R[407][1] = r_cell_wire[407];							inform_R[408][1] = r_cell_wire[408];							inform_R[409][1] = r_cell_wire[409];							inform_R[410][1] = r_cell_wire[410];							inform_R[411][1] = r_cell_wire[411];							inform_R[412][1] = r_cell_wire[412];							inform_R[413][1] = r_cell_wire[413];							inform_R[414][1] = r_cell_wire[414];							inform_R[415][1] = r_cell_wire[415];							inform_R[416][1] = r_cell_wire[416];							inform_R[417][1] = r_cell_wire[417];							inform_R[418][1] = r_cell_wire[418];							inform_R[419][1] = r_cell_wire[419];							inform_R[420][1] = r_cell_wire[420];							inform_R[421][1] = r_cell_wire[421];							inform_R[422][1] = r_cell_wire[422];							inform_R[423][1] = r_cell_wire[423];							inform_R[424][1] = r_cell_wire[424];							inform_R[425][1] = r_cell_wire[425];							inform_R[426][1] = r_cell_wire[426];							inform_R[427][1] = r_cell_wire[427];							inform_R[428][1] = r_cell_wire[428];							inform_R[429][1] = r_cell_wire[429];							inform_R[430][1] = r_cell_wire[430];							inform_R[431][1] = r_cell_wire[431];							inform_R[432][1] = r_cell_wire[432];							inform_R[433][1] = r_cell_wire[433];							inform_R[434][1] = r_cell_wire[434];							inform_R[435][1] = r_cell_wire[435];							inform_R[436][1] = r_cell_wire[436];							inform_R[437][1] = r_cell_wire[437];							inform_R[438][1] = r_cell_wire[438];							inform_R[439][1] = r_cell_wire[439];							inform_R[440][1] = r_cell_wire[440];							inform_R[441][1] = r_cell_wire[441];							inform_R[442][1] = r_cell_wire[442];							inform_R[443][1] = r_cell_wire[443];							inform_R[444][1] = r_cell_wire[444];							inform_R[445][1] = r_cell_wire[445];							inform_R[446][1] = r_cell_wire[446];							inform_R[447][1] = r_cell_wire[447];							inform_R[448][1] = r_cell_wire[448];							inform_R[449][1] = r_cell_wire[449];							inform_R[450][1] = r_cell_wire[450];							inform_R[451][1] = r_cell_wire[451];							inform_R[452][1] = r_cell_wire[452];							inform_R[453][1] = r_cell_wire[453];							inform_R[454][1] = r_cell_wire[454];							inform_R[455][1] = r_cell_wire[455];							inform_R[456][1] = r_cell_wire[456];							inform_R[457][1] = r_cell_wire[457];							inform_R[458][1] = r_cell_wire[458];							inform_R[459][1] = r_cell_wire[459];							inform_R[460][1] = r_cell_wire[460];							inform_R[461][1] = r_cell_wire[461];							inform_R[462][1] = r_cell_wire[462];							inform_R[463][1] = r_cell_wire[463];							inform_R[464][1] = r_cell_wire[464];							inform_R[465][1] = r_cell_wire[465];							inform_R[466][1] = r_cell_wire[466];							inform_R[467][1] = r_cell_wire[467];							inform_R[468][1] = r_cell_wire[468];							inform_R[469][1] = r_cell_wire[469];							inform_R[470][1] = r_cell_wire[470];							inform_R[471][1] = r_cell_wire[471];							inform_R[472][1] = r_cell_wire[472];							inform_R[473][1] = r_cell_wire[473];							inform_R[474][1] = r_cell_wire[474];							inform_R[475][1] = r_cell_wire[475];							inform_R[476][1] = r_cell_wire[476];							inform_R[477][1] = r_cell_wire[477];							inform_R[478][1] = r_cell_wire[478];							inform_R[479][1] = r_cell_wire[479];							inform_R[480][1] = r_cell_wire[480];							inform_R[481][1] = r_cell_wire[481];							inform_R[482][1] = r_cell_wire[482];							inform_R[483][1] = r_cell_wire[483];							inform_R[484][1] = r_cell_wire[484];							inform_R[485][1] = r_cell_wire[485];							inform_R[486][1] = r_cell_wire[486];							inform_R[487][1] = r_cell_wire[487];							inform_R[488][1] = r_cell_wire[488];							inform_R[489][1] = r_cell_wire[489];							inform_R[490][1] = r_cell_wire[490];							inform_R[491][1] = r_cell_wire[491];							inform_R[492][1] = r_cell_wire[492];							inform_R[493][1] = r_cell_wire[493];							inform_R[494][1] = r_cell_wire[494];							inform_R[495][1] = r_cell_wire[495];							inform_R[496][1] = r_cell_wire[496];							inform_R[497][1] = r_cell_wire[497];							inform_R[498][1] = r_cell_wire[498];							inform_R[499][1] = r_cell_wire[499];							inform_R[500][1] = r_cell_wire[500];							inform_R[501][1] = r_cell_wire[501];							inform_R[502][1] = r_cell_wire[502];							inform_R[503][1] = r_cell_wire[503];							inform_R[504][1] = r_cell_wire[504];							inform_R[505][1] = r_cell_wire[505];							inform_R[506][1] = r_cell_wire[506];							inform_R[507][1] = r_cell_wire[507];							inform_R[508][1] = r_cell_wire[508];							inform_R[509][1] = r_cell_wire[509];							inform_R[510][1] = r_cell_wire[510];							inform_R[511][1] = r_cell_wire[511];							inform_R[512][1] = r_cell_wire[512];							inform_R[513][1] = r_cell_wire[513];							inform_R[514][1] = r_cell_wire[514];							inform_R[515][1] = r_cell_wire[515];							inform_R[516][1] = r_cell_wire[516];							inform_R[517][1] = r_cell_wire[517];							inform_R[518][1] = r_cell_wire[518];							inform_R[519][1] = r_cell_wire[519];							inform_R[520][1] = r_cell_wire[520];							inform_R[521][1] = r_cell_wire[521];							inform_R[522][1] = r_cell_wire[522];							inform_R[523][1] = r_cell_wire[523];							inform_R[524][1] = r_cell_wire[524];							inform_R[525][1] = r_cell_wire[525];							inform_R[526][1] = r_cell_wire[526];							inform_R[527][1] = r_cell_wire[527];							inform_R[528][1] = r_cell_wire[528];							inform_R[529][1] = r_cell_wire[529];							inform_R[530][1] = r_cell_wire[530];							inform_R[531][1] = r_cell_wire[531];							inform_R[532][1] = r_cell_wire[532];							inform_R[533][1] = r_cell_wire[533];							inform_R[534][1] = r_cell_wire[534];							inform_R[535][1] = r_cell_wire[535];							inform_R[536][1] = r_cell_wire[536];							inform_R[537][1] = r_cell_wire[537];							inform_R[538][1] = r_cell_wire[538];							inform_R[539][1] = r_cell_wire[539];							inform_R[540][1] = r_cell_wire[540];							inform_R[541][1] = r_cell_wire[541];							inform_R[542][1] = r_cell_wire[542];							inform_R[543][1] = r_cell_wire[543];							inform_R[544][1] = r_cell_wire[544];							inform_R[545][1] = r_cell_wire[545];							inform_R[546][1] = r_cell_wire[546];							inform_R[547][1] = r_cell_wire[547];							inform_R[548][1] = r_cell_wire[548];							inform_R[549][1] = r_cell_wire[549];							inform_R[550][1] = r_cell_wire[550];							inform_R[551][1] = r_cell_wire[551];							inform_R[552][1] = r_cell_wire[552];							inform_R[553][1] = r_cell_wire[553];							inform_R[554][1] = r_cell_wire[554];							inform_R[555][1] = r_cell_wire[555];							inform_R[556][1] = r_cell_wire[556];							inform_R[557][1] = r_cell_wire[557];							inform_R[558][1] = r_cell_wire[558];							inform_R[559][1] = r_cell_wire[559];							inform_R[560][1] = r_cell_wire[560];							inform_R[561][1] = r_cell_wire[561];							inform_R[562][1] = r_cell_wire[562];							inform_R[563][1] = r_cell_wire[563];							inform_R[564][1] = r_cell_wire[564];							inform_R[565][1] = r_cell_wire[565];							inform_R[566][1] = r_cell_wire[566];							inform_R[567][1] = r_cell_wire[567];							inform_R[568][1] = r_cell_wire[568];							inform_R[569][1] = r_cell_wire[569];							inform_R[570][1] = r_cell_wire[570];							inform_R[571][1] = r_cell_wire[571];							inform_R[572][1] = r_cell_wire[572];							inform_R[573][1] = r_cell_wire[573];							inform_R[574][1] = r_cell_wire[574];							inform_R[575][1] = r_cell_wire[575];							inform_R[576][1] = r_cell_wire[576];							inform_R[577][1] = r_cell_wire[577];							inform_R[578][1] = r_cell_wire[578];							inform_R[579][1] = r_cell_wire[579];							inform_R[580][1] = r_cell_wire[580];							inform_R[581][1] = r_cell_wire[581];							inform_R[582][1] = r_cell_wire[582];							inform_R[583][1] = r_cell_wire[583];							inform_R[584][1] = r_cell_wire[584];							inform_R[585][1] = r_cell_wire[585];							inform_R[586][1] = r_cell_wire[586];							inform_R[587][1] = r_cell_wire[587];							inform_R[588][1] = r_cell_wire[588];							inform_R[589][1] = r_cell_wire[589];							inform_R[590][1] = r_cell_wire[590];							inform_R[591][1] = r_cell_wire[591];							inform_R[592][1] = r_cell_wire[592];							inform_R[593][1] = r_cell_wire[593];							inform_R[594][1] = r_cell_wire[594];							inform_R[595][1] = r_cell_wire[595];							inform_R[596][1] = r_cell_wire[596];							inform_R[597][1] = r_cell_wire[597];							inform_R[598][1] = r_cell_wire[598];							inform_R[599][1] = r_cell_wire[599];							inform_R[600][1] = r_cell_wire[600];							inform_R[601][1] = r_cell_wire[601];							inform_R[602][1] = r_cell_wire[602];							inform_R[603][1] = r_cell_wire[603];							inform_R[604][1] = r_cell_wire[604];							inform_R[605][1] = r_cell_wire[605];							inform_R[606][1] = r_cell_wire[606];							inform_R[607][1] = r_cell_wire[607];							inform_R[608][1] = r_cell_wire[608];							inform_R[609][1] = r_cell_wire[609];							inform_R[610][1] = r_cell_wire[610];							inform_R[611][1] = r_cell_wire[611];							inform_R[612][1] = r_cell_wire[612];							inform_R[613][1] = r_cell_wire[613];							inform_R[614][1] = r_cell_wire[614];							inform_R[615][1] = r_cell_wire[615];							inform_R[616][1] = r_cell_wire[616];							inform_R[617][1] = r_cell_wire[617];							inform_R[618][1] = r_cell_wire[618];							inform_R[619][1] = r_cell_wire[619];							inform_R[620][1] = r_cell_wire[620];							inform_R[621][1] = r_cell_wire[621];							inform_R[622][1] = r_cell_wire[622];							inform_R[623][1] = r_cell_wire[623];							inform_R[624][1] = r_cell_wire[624];							inform_R[625][1] = r_cell_wire[625];							inform_R[626][1] = r_cell_wire[626];							inform_R[627][1] = r_cell_wire[627];							inform_R[628][1] = r_cell_wire[628];							inform_R[629][1] = r_cell_wire[629];							inform_R[630][1] = r_cell_wire[630];							inform_R[631][1] = r_cell_wire[631];							inform_R[632][1] = r_cell_wire[632];							inform_R[633][1] = r_cell_wire[633];							inform_R[634][1] = r_cell_wire[634];							inform_R[635][1] = r_cell_wire[635];							inform_R[636][1] = r_cell_wire[636];							inform_R[637][1] = r_cell_wire[637];							inform_R[638][1] = r_cell_wire[638];							inform_R[639][1] = r_cell_wire[639];							inform_R[640][1] = r_cell_wire[640];							inform_R[641][1] = r_cell_wire[641];							inform_R[642][1] = r_cell_wire[642];							inform_R[643][1] = r_cell_wire[643];							inform_R[644][1] = r_cell_wire[644];							inform_R[645][1] = r_cell_wire[645];							inform_R[646][1] = r_cell_wire[646];							inform_R[647][1] = r_cell_wire[647];							inform_R[648][1] = r_cell_wire[648];							inform_R[649][1] = r_cell_wire[649];							inform_R[650][1] = r_cell_wire[650];							inform_R[651][1] = r_cell_wire[651];							inform_R[652][1] = r_cell_wire[652];							inform_R[653][1] = r_cell_wire[653];							inform_R[654][1] = r_cell_wire[654];							inform_R[655][1] = r_cell_wire[655];							inform_R[656][1] = r_cell_wire[656];							inform_R[657][1] = r_cell_wire[657];							inform_R[658][1] = r_cell_wire[658];							inform_R[659][1] = r_cell_wire[659];							inform_R[660][1] = r_cell_wire[660];							inform_R[661][1] = r_cell_wire[661];							inform_R[662][1] = r_cell_wire[662];							inform_R[663][1] = r_cell_wire[663];							inform_R[664][1] = r_cell_wire[664];							inform_R[665][1] = r_cell_wire[665];							inform_R[666][1] = r_cell_wire[666];							inform_R[667][1] = r_cell_wire[667];							inform_R[668][1] = r_cell_wire[668];							inform_R[669][1] = r_cell_wire[669];							inform_R[670][1] = r_cell_wire[670];							inform_R[671][1] = r_cell_wire[671];							inform_R[672][1] = r_cell_wire[672];							inform_R[673][1] = r_cell_wire[673];							inform_R[674][1] = r_cell_wire[674];							inform_R[675][1] = r_cell_wire[675];							inform_R[676][1] = r_cell_wire[676];							inform_R[677][1] = r_cell_wire[677];							inform_R[678][1] = r_cell_wire[678];							inform_R[679][1] = r_cell_wire[679];							inform_R[680][1] = r_cell_wire[680];							inform_R[681][1] = r_cell_wire[681];							inform_R[682][1] = r_cell_wire[682];							inform_R[683][1] = r_cell_wire[683];							inform_R[684][1] = r_cell_wire[684];							inform_R[685][1] = r_cell_wire[685];							inform_R[686][1] = r_cell_wire[686];							inform_R[687][1] = r_cell_wire[687];							inform_R[688][1] = r_cell_wire[688];							inform_R[689][1] = r_cell_wire[689];							inform_R[690][1] = r_cell_wire[690];							inform_R[691][1] = r_cell_wire[691];							inform_R[692][1] = r_cell_wire[692];							inform_R[693][1] = r_cell_wire[693];							inform_R[694][1] = r_cell_wire[694];							inform_R[695][1] = r_cell_wire[695];							inform_R[696][1] = r_cell_wire[696];							inform_R[697][1] = r_cell_wire[697];							inform_R[698][1] = r_cell_wire[698];							inform_R[699][1] = r_cell_wire[699];							inform_R[700][1] = r_cell_wire[700];							inform_R[701][1] = r_cell_wire[701];							inform_R[702][1] = r_cell_wire[702];							inform_R[703][1] = r_cell_wire[703];							inform_R[704][1] = r_cell_wire[704];							inform_R[705][1] = r_cell_wire[705];							inform_R[706][1] = r_cell_wire[706];							inform_R[707][1] = r_cell_wire[707];							inform_R[708][1] = r_cell_wire[708];							inform_R[709][1] = r_cell_wire[709];							inform_R[710][1] = r_cell_wire[710];							inform_R[711][1] = r_cell_wire[711];							inform_R[712][1] = r_cell_wire[712];							inform_R[713][1] = r_cell_wire[713];							inform_R[714][1] = r_cell_wire[714];							inform_R[715][1] = r_cell_wire[715];							inform_R[716][1] = r_cell_wire[716];							inform_R[717][1] = r_cell_wire[717];							inform_R[718][1] = r_cell_wire[718];							inform_R[719][1] = r_cell_wire[719];							inform_R[720][1] = r_cell_wire[720];							inform_R[721][1] = r_cell_wire[721];							inform_R[722][1] = r_cell_wire[722];							inform_R[723][1] = r_cell_wire[723];							inform_R[724][1] = r_cell_wire[724];							inform_R[725][1] = r_cell_wire[725];							inform_R[726][1] = r_cell_wire[726];							inform_R[727][1] = r_cell_wire[727];							inform_R[728][1] = r_cell_wire[728];							inform_R[729][1] = r_cell_wire[729];							inform_R[730][1] = r_cell_wire[730];							inform_R[731][1] = r_cell_wire[731];							inform_R[732][1] = r_cell_wire[732];							inform_R[733][1] = r_cell_wire[733];							inform_R[734][1] = r_cell_wire[734];							inform_R[735][1] = r_cell_wire[735];							inform_R[736][1] = r_cell_wire[736];							inform_R[737][1] = r_cell_wire[737];							inform_R[738][1] = r_cell_wire[738];							inform_R[739][1] = r_cell_wire[739];							inform_R[740][1] = r_cell_wire[740];							inform_R[741][1] = r_cell_wire[741];							inform_R[742][1] = r_cell_wire[742];							inform_R[743][1] = r_cell_wire[743];							inform_R[744][1] = r_cell_wire[744];							inform_R[745][1] = r_cell_wire[745];							inform_R[746][1] = r_cell_wire[746];							inform_R[747][1] = r_cell_wire[747];							inform_R[748][1] = r_cell_wire[748];							inform_R[749][1] = r_cell_wire[749];							inform_R[750][1] = r_cell_wire[750];							inform_R[751][1] = r_cell_wire[751];							inform_R[752][1] = r_cell_wire[752];							inform_R[753][1] = r_cell_wire[753];							inform_R[754][1] = r_cell_wire[754];							inform_R[755][1] = r_cell_wire[755];							inform_R[756][1] = r_cell_wire[756];							inform_R[757][1] = r_cell_wire[757];							inform_R[758][1] = r_cell_wire[758];							inform_R[759][1] = r_cell_wire[759];							inform_R[760][1] = r_cell_wire[760];							inform_R[761][1] = r_cell_wire[761];							inform_R[762][1] = r_cell_wire[762];							inform_R[763][1] = r_cell_wire[763];							inform_R[764][1] = r_cell_wire[764];							inform_R[765][1] = r_cell_wire[765];							inform_R[766][1] = r_cell_wire[766];							inform_R[767][1] = r_cell_wire[767];							inform_R[768][1] = r_cell_wire[768];							inform_R[769][1] = r_cell_wire[769];							inform_R[770][1] = r_cell_wire[770];							inform_R[771][1] = r_cell_wire[771];							inform_R[772][1] = r_cell_wire[772];							inform_R[773][1] = r_cell_wire[773];							inform_R[774][1] = r_cell_wire[774];							inform_R[775][1] = r_cell_wire[775];							inform_R[776][1] = r_cell_wire[776];							inform_R[777][1] = r_cell_wire[777];							inform_R[778][1] = r_cell_wire[778];							inform_R[779][1] = r_cell_wire[779];							inform_R[780][1] = r_cell_wire[780];							inform_R[781][1] = r_cell_wire[781];							inform_R[782][1] = r_cell_wire[782];							inform_R[783][1] = r_cell_wire[783];							inform_R[784][1] = r_cell_wire[784];							inform_R[785][1] = r_cell_wire[785];							inform_R[786][1] = r_cell_wire[786];							inform_R[787][1] = r_cell_wire[787];							inform_R[788][1] = r_cell_wire[788];							inform_R[789][1] = r_cell_wire[789];							inform_R[790][1] = r_cell_wire[790];							inform_R[791][1] = r_cell_wire[791];							inform_R[792][1] = r_cell_wire[792];							inform_R[793][1] = r_cell_wire[793];							inform_R[794][1] = r_cell_wire[794];							inform_R[795][1] = r_cell_wire[795];							inform_R[796][1] = r_cell_wire[796];							inform_R[797][1] = r_cell_wire[797];							inform_R[798][1] = r_cell_wire[798];							inform_R[799][1] = r_cell_wire[799];							inform_R[800][1] = r_cell_wire[800];							inform_R[801][1] = r_cell_wire[801];							inform_R[802][1] = r_cell_wire[802];							inform_R[803][1] = r_cell_wire[803];							inform_R[804][1] = r_cell_wire[804];							inform_R[805][1] = r_cell_wire[805];							inform_R[806][1] = r_cell_wire[806];							inform_R[807][1] = r_cell_wire[807];							inform_R[808][1] = r_cell_wire[808];							inform_R[809][1] = r_cell_wire[809];							inform_R[810][1] = r_cell_wire[810];							inform_R[811][1] = r_cell_wire[811];							inform_R[812][1] = r_cell_wire[812];							inform_R[813][1] = r_cell_wire[813];							inform_R[814][1] = r_cell_wire[814];							inform_R[815][1] = r_cell_wire[815];							inform_R[816][1] = r_cell_wire[816];							inform_R[817][1] = r_cell_wire[817];							inform_R[818][1] = r_cell_wire[818];							inform_R[819][1] = r_cell_wire[819];							inform_R[820][1] = r_cell_wire[820];							inform_R[821][1] = r_cell_wire[821];							inform_R[822][1] = r_cell_wire[822];							inform_R[823][1] = r_cell_wire[823];							inform_R[824][1] = r_cell_wire[824];							inform_R[825][1] = r_cell_wire[825];							inform_R[826][1] = r_cell_wire[826];							inform_R[827][1] = r_cell_wire[827];							inform_R[828][1] = r_cell_wire[828];							inform_R[829][1] = r_cell_wire[829];							inform_R[830][1] = r_cell_wire[830];							inform_R[831][1] = r_cell_wire[831];							inform_R[832][1] = r_cell_wire[832];							inform_R[833][1] = r_cell_wire[833];							inform_R[834][1] = r_cell_wire[834];							inform_R[835][1] = r_cell_wire[835];							inform_R[836][1] = r_cell_wire[836];							inform_R[837][1] = r_cell_wire[837];							inform_R[838][1] = r_cell_wire[838];							inform_R[839][1] = r_cell_wire[839];							inform_R[840][1] = r_cell_wire[840];							inform_R[841][1] = r_cell_wire[841];							inform_R[842][1] = r_cell_wire[842];							inform_R[843][1] = r_cell_wire[843];							inform_R[844][1] = r_cell_wire[844];							inform_R[845][1] = r_cell_wire[845];							inform_R[846][1] = r_cell_wire[846];							inform_R[847][1] = r_cell_wire[847];							inform_R[848][1] = r_cell_wire[848];							inform_R[849][1] = r_cell_wire[849];							inform_R[850][1] = r_cell_wire[850];							inform_R[851][1] = r_cell_wire[851];							inform_R[852][1] = r_cell_wire[852];							inform_R[853][1] = r_cell_wire[853];							inform_R[854][1] = r_cell_wire[854];							inform_R[855][1] = r_cell_wire[855];							inform_R[856][1] = r_cell_wire[856];							inform_R[857][1] = r_cell_wire[857];							inform_R[858][1] = r_cell_wire[858];							inform_R[859][1] = r_cell_wire[859];							inform_R[860][1] = r_cell_wire[860];							inform_R[861][1] = r_cell_wire[861];							inform_R[862][1] = r_cell_wire[862];							inform_R[863][1] = r_cell_wire[863];							inform_R[864][1] = r_cell_wire[864];							inform_R[865][1] = r_cell_wire[865];							inform_R[866][1] = r_cell_wire[866];							inform_R[867][1] = r_cell_wire[867];							inform_R[868][1] = r_cell_wire[868];							inform_R[869][1] = r_cell_wire[869];							inform_R[870][1] = r_cell_wire[870];							inform_R[871][1] = r_cell_wire[871];							inform_R[872][1] = r_cell_wire[872];							inform_R[873][1] = r_cell_wire[873];							inform_R[874][1] = r_cell_wire[874];							inform_R[875][1] = r_cell_wire[875];							inform_R[876][1] = r_cell_wire[876];							inform_R[877][1] = r_cell_wire[877];							inform_R[878][1] = r_cell_wire[878];							inform_R[879][1] = r_cell_wire[879];							inform_R[880][1] = r_cell_wire[880];							inform_R[881][1] = r_cell_wire[881];							inform_R[882][1] = r_cell_wire[882];							inform_R[883][1] = r_cell_wire[883];							inform_R[884][1] = r_cell_wire[884];							inform_R[885][1] = r_cell_wire[885];							inform_R[886][1] = r_cell_wire[886];							inform_R[887][1] = r_cell_wire[887];							inform_R[888][1] = r_cell_wire[888];							inform_R[889][1] = r_cell_wire[889];							inform_R[890][1] = r_cell_wire[890];							inform_R[891][1] = r_cell_wire[891];							inform_R[892][1] = r_cell_wire[892];							inform_R[893][1] = r_cell_wire[893];							inform_R[894][1] = r_cell_wire[894];							inform_R[895][1] = r_cell_wire[895];							inform_R[896][1] = r_cell_wire[896];							inform_R[897][1] = r_cell_wire[897];							inform_R[898][1] = r_cell_wire[898];							inform_R[899][1] = r_cell_wire[899];							inform_R[900][1] = r_cell_wire[900];							inform_R[901][1] = r_cell_wire[901];							inform_R[902][1] = r_cell_wire[902];							inform_R[903][1] = r_cell_wire[903];							inform_R[904][1] = r_cell_wire[904];							inform_R[905][1] = r_cell_wire[905];							inform_R[906][1] = r_cell_wire[906];							inform_R[907][1] = r_cell_wire[907];							inform_R[908][1] = r_cell_wire[908];							inform_R[909][1] = r_cell_wire[909];							inform_R[910][1] = r_cell_wire[910];							inform_R[911][1] = r_cell_wire[911];							inform_R[912][1] = r_cell_wire[912];							inform_R[913][1] = r_cell_wire[913];							inform_R[914][1] = r_cell_wire[914];							inform_R[915][1] = r_cell_wire[915];							inform_R[916][1] = r_cell_wire[916];							inform_R[917][1] = r_cell_wire[917];							inform_R[918][1] = r_cell_wire[918];							inform_R[919][1] = r_cell_wire[919];							inform_R[920][1] = r_cell_wire[920];							inform_R[921][1] = r_cell_wire[921];							inform_R[922][1] = r_cell_wire[922];							inform_R[923][1] = r_cell_wire[923];							inform_R[924][1] = r_cell_wire[924];							inform_R[925][1] = r_cell_wire[925];							inform_R[926][1] = r_cell_wire[926];							inform_R[927][1] = r_cell_wire[927];							inform_R[928][1] = r_cell_wire[928];							inform_R[929][1] = r_cell_wire[929];							inform_R[930][1] = r_cell_wire[930];							inform_R[931][1] = r_cell_wire[931];							inform_R[932][1] = r_cell_wire[932];							inform_R[933][1] = r_cell_wire[933];							inform_R[934][1] = r_cell_wire[934];							inform_R[935][1] = r_cell_wire[935];							inform_R[936][1] = r_cell_wire[936];							inform_R[937][1] = r_cell_wire[937];							inform_R[938][1] = r_cell_wire[938];							inform_R[939][1] = r_cell_wire[939];							inform_R[940][1] = r_cell_wire[940];							inform_R[941][1] = r_cell_wire[941];							inform_R[942][1] = r_cell_wire[942];							inform_R[943][1] = r_cell_wire[943];							inform_R[944][1] = r_cell_wire[944];							inform_R[945][1] = r_cell_wire[945];							inform_R[946][1] = r_cell_wire[946];							inform_R[947][1] = r_cell_wire[947];							inform_R[948][1] = r_cell_wire[948];							inform_R[949][1] = r_cell_wire[949];							inform_R[950][1] = r_cell_wire[950];							inform_R[951][1] = r_cell_wire[951];							inform_R[952][1] = r_cell_wire[952];							inform_R[953][1] = r_cell_wire[953];							inform_R[954][1] = r_cell_wire[954];							inform_R[955][1] = r_cell_wire[955];							inform_R[956][1] = r_cell_wire[956];							inform_R[957][1] = r_cell_wire[957];							inform_R[958][1] = r_cell_wire[958];							inform_R[959][1] = r_cell_wire[959];							inform_R[960][1] = r_cell_wire[960];							inform_R[961][1] = r_cell_wire[961];							inform_R[962][1] = r_cell_wire[962];							inform_R[963][1] = r_cell_wire[963];							inform_R[964][1] = r_cell_wire[964];							inform_R[965][1] = r_cell_wire[965];							inform_R[966][1] = r_cell_wire[966];							inform_R[967][1] = r_cell_wire[967];							inform_R[968][1] = r_cell_wire[968];							inform_R[969][1] = r_cell_wire[969];							inform_R[970][1] = r_cell_wire[970];							inform_R[971][1] = r_cell_wire[971];							inform_R[972][1] = r_cell_wire[972];							inform_R[973][1] = r_cell_wire[973];							inform_R[974][1] = r_cell_wire[974];							inform_R[975][1] = r_cell_wire[975];							inform_R[976][1] = r_cell_wire[976];							inform_R[977][1] = r_cell_wire[977];							inform_R[978][1] = r_cell_wire[978];							inform_R[979][1] = r_cell_wire[979];							inform_R[980][1] = r_cell_wire[980];							inform_R[981][1] = r_cell_wire[981];							inform_R[982][1] = r_cell_wire[982];							inform_R[983][1] = r_cell_wire[983];							inform_R[984][1] = r_cell_wire[984];							inform_R[985][1] = r_cell_wire[985];							inform_R[986][1] = r_cell_wire[986];							inform_R[987][1] = r_cell_wire[987];							inform_R[988][1] = r_cell_wire[988];							inform_R[989][1] = r_cell_wire[989];							inform_R[990][1] = r_cell_wire[990];							inform_R[991][1] = r_cell_wire[991];							inform_R[992][1] = r_cell_wire[992];							inform_R[993][1] = r_cell_wire[993];							inform_R[994][1] = r_cell_wire[994];							inform_R[995][1] = r_cell_wire[995];							inform_R[996][1] = r_cell_wire[996];							inform_R[997][1] = r_cell_wire[997];							inform_R[998][1] = r_cell_wire[998];							inform_R[999][1] = r_cell_wire[999];							inform_R[1000][1] = r_cell_wire[1000];							inform_R[1001][1] = r_cell_wire[1001];							inform_R[1002][1] = r_cell_wire[1002];							inform_R[1003][1] = r_cell_wire[1003];							inform_R[1004][1] = r_cell_wire[1004];							inform_R[1005][1] = r_cell_wire[1005];							inform_R[1006][1] = r_cell_wire[1006];							inform_R[1007][1] = r_cell_wire[1007];							inform_R[1008][1] = r_cell_wire[1008];							inform_R[1009][1] = r_cell_wire[1009];							inform_R[1010][1] = r_cell_wire[1010];							inform_R[1011][1] = r_cell_wire[1011];							inform_R[1012][1] = r_cell_wire[1012];							inform_R[1013][1] = r_cell_wire[1013];							inform_R[1014][1] = r_cell_wire[1014];							inform_R[1015][1] = r_cell_wire[1015];							inform_R[1016][1] = r_cell_wire[1016];							inform_R[1017][1] = r_cell_wire[1017];							inform_R[1018][1] = r_cell_wire[1018];							inform_R[1019][1] = r_cell_wire[1019];							inform_R[1020][1] = r_cell_wire[1020];							inform_R[1021][1] = r_cell_wire[1021];							inform_R[1022][1] = r_cell_wire[1022];							inform_R[1023][1] = r_cell_wire[1023];							inform_L[0][0] = l_cell_wire[0];							inform_L[1][0] = l_cell_wire[1];							inform_L[2][0] = l_cell_wire[2];							inform_L[3][0] = l_cell_wire[3];							inform_L[4][0] = l_cell_wire[4];							inform_L[5][0] = l_cell_wire[5];							inform_L[6][0] = l_cell_wire[6];							inform_L[7][0] = l_cell_wire[7];							inform_L[8][0] = l_cell_wire[8];							inform_L[9][0] = l_cell_wire[9];							inform_L[10][0] = l_cell_wire[10];							inform_L[11][0] = l_cell_wire[11];							inform_L[12][0] = l_cell_wire[12];							inform_L[13][0] = l_cell_wire[13];							inform_L[14][0] = l_cell_wire[14];							inform_L[15][0] = l_cell_wire[15];							inform_L[16][0] = l_cell_wire[16];							inform_L[17][0] = l_cell_wire[17];							inform_L[18][0] = l_cell_wire[18];							inform_L[19][0] = l_cell_wire[19];							inform_L[20][0] = l_cell_wire[20];							inform_L[21][0] = l_cell_wire[21];							inform_L[22][0] = l_cell_wire[22];							inform_L[23][0] = l_cell_wire[23];							inform_L[24][0] = l_cell_wire[24];							inform_L[25][0] = l_cell_wire[25];							inform_L[26][0] = l_cell_wire[26];							inform_L[27][0] = l_cell_wire[27];							inform_L[28][0] = l_cell_wire[28];							inform_L[29][0] = l_cell_wire[29];							inform_L[30][0] = l_cell_wire[30];							inform_L[31][0] = l_cell_wire[31];							inform_L[32][0] = l_cell_wire[32];							inform_L[33][0] = l_cell_wire[33];							inform_L[34][0] = l_cell_wire[34];							inform_L[35][0] = l_cell_wire[35];							inform_L[36][0] = l_cell_wire[36];							inform_L[37][0] = l_cell_wire[37];							inform_L[38][0] = l_cell_wire[38];							inform_L[39][0] = l_cell_wire[39];							inform_L[40][0] = l_cell_wire[40];							inform_L[41][0] = l_cell_wire[41];							inform_L[42][0] = l_cell_wire[42];							inform_L[43][0] = l_cell_wire[43];							inform_L[44][0] = l_cell_wire[44];							inform_L[45][0] = l_cell_wire[45];							inform_L[46][0] = l_cell_wire[46];							inform_L[47][0] = l_cell_wire[47];							inform_L[48][0] = l_cell_wire[48];							inform_L[49][0] = l_cell_wire[49];							inform_L[50][0] = l_cell_wire[50];							inform_L[51][0] = l_cell_wire[51];							inform_L[52][0] = l_cell_wire[52];							inform_L[53][0] = l_cell_wire[53];							inform_L[54][0] = l_cell_wire[54];							inform_L[55][0] = l_cell_wire[55];							inform_L[56][0] = l_cell_wire[56];							inform_L[57][0] = l_cell_wire[57];							inform_L[58][0] = l_cell_wire[58];							inform_L[59][0] = l_cell_wire[59];							inform_L[60][0] = l_cell_wire[60];							inform_L[61][0] = l_cell_wire[61];							inform_L[62][0] = l_cell_wire[62];							inform_L[63][0] = l_cell_wire[63];							inform_L[64][0] = l_cell_wire[64];							inform_L[65][0] = l_cell_wire[65];							inform_L[66][0] = l_cell_wire[66];							inform_L[67][0] = l_cell_wire[67];							inform_L[68][0] = l_cell_wire[68];							inform_L[69][0] = l_cell_wire[69];							inform_L[70][0] = l_cell_wire[70];							inform_L[71][0] = l_cell_wire[71];							inform_L[72][0] = l_cell_wire[72];							inform_L[73][0] = l_cell_wire[73];							inform_L[74][0] = l_cell_wire[74];							inform_L[75][0] = l_cell_wire[75];							inform_L[76][0] = l_cell_wire[76];							inform_L[77][0] = l_cell_wire[77];							inform_L[78][0] = l_cell_wire[78];							inform_L[79][0] = l_cell_wire[79];							inform_L[80][0] = l_cell_wire[80];							inform_L[81][0] = l_cell_wire[81];							inform_L[82][0] = l_cell_wire[82];							inform_L[83][0] = l_cell_wire[83];							inform_L[84][0] = l_cell_wire[84];							inform_L[85][0] = l_cell_wire[85];							inform_L[86][0] = l_cell_wire[86];							inform_L[87][0] = l_cell_wire[87];							inform_L[88][0] = l_cell_wire[88];							inform_L[89][0] = l_cell_wire[89];							inform_L[90][0] = l_cell_wire[90];							inform_L[91][0] = l_cell_wire[91];							inform_L[92][0] = l_cell_wire[92];							inform_L[93][0] = l_cell_wire[93];							inform_L[94][0] = l_cell_wire[94];							inform_L[95][0] = l_cell_wire[95];							inform_L[96][0] = l_cell_wire[96];							inform_L[97][0] = l_cell_wire[97];							inform_L[98][0] = l_cell_wire[98];							inform_L[99][0] = l_cell_wire[99];							inform_L[100][0] = l_cell_wire[100];							inform_L[101][0] = l_cell_wire[101];							inform_L[102][0] = l_cell_wire[102];							inform_L[103][0] = l_cell_wire[103];							inform_L[104][0] = l_cell_wire[104];							inform_L[105][0] = l_cell_wire[105];							inform_L[106][0] = l_cell_wire[106];							inform_L[107][0] = l_cell_wire[107];							inform_L[108][0] = l_cell_wire[108];							inform_L[109][0] = l_cell_wire[109];							inform_L[110][0] = l_cell_wire[110];							inform_L[111][0] = l_cell_wire[111];							inform_L[112][0] = l_cell_wire[112];							inform_L[113][0] = l_cell_wire[113];							inform_L[114][0] = l_cell_wire[114];							inform_L[115][0] = l_cell_wire[115];							inform_L[116][0] = l_cell_wire[116];							inform_L[117][0] = l_cell_wire[117];							inform_L[118][0] = l_cell_wire[118];							inform_L[119][0] = l_cell_wire[119];							inform_L[120][0] = l_cell_wire[120];							inform_L[121][0] = l_cell_wire[121];							inform_L[122][0] = l_cell_wire[122];							inform_L[123][0] = l_cell_wire[123];							inform_L[124][0] = l_cell_wire[124];							inform_L[125][0] = l_cell_wire[125];							inform_L[126][0] = l_cell_wire[126];							inform_L[127][0] = l_cell_wire[127];							inform_L[128][0] = l_cell_wire[128];							inform_L[129][0] = l_cell_wire[129];							inform_L[130][0] = l_cell_wire[130];							inform_L[131][0] = l_cell_wire[131];							inform_L[132][0] = l_cell_wire[132];							inform_L[133][0] = l_cell_wire[133];							inform_L[134][0] = l_cell_wire[134];							inform_L[135][0] = l_cell_wire[135];							inform_L[136][0] = l_cell_wire[136];							inform_L[137][0] = l_cell_wire[137];							inform_L[138][0] = l_cell_wire[138];							inform_L[139][0] = l_cell_wire[139];							inform_L[140][0] = l_cell_wire[140];							inform_L[141][0] = l_cell_wire[141];							inform_L[142][0] = l_cell_wire[142];							inform_L[143][0] = l_cell_wire[143];							inform_L[144][0] = l_cell_wire[144];							inform_L[145][0] = l_cell_wire[145];							inform_L[146][0] = l_cell_wire[146];							inform_L[147][0] = l_cell_wire[147];							inform_L[148][0] = l_cell_wire[148];							inform_L[149][0] = l_cell_wire[149];							inform_L[150][0] = l_cell_wire[150];							inform_L[151][0] = l_cell_wire[151];							inform_L[152][0] = l_cell_wire[152];							inform_L[153][0] = l_cell_wire[153];							inform_L[154][0] = l_cell_wire[154];							inform_L[155][0] = l_cell_wire[155];							inform_L[156][0] = l_cell_wire[156];							inform_L[157][0] = l_cell_wire[157];							inform_L[158][0] = l_cell_wire[158];							inform_L[159][0] = l_cell_wire[159];							inform_L[160][0] = l_cell_wire[160];							inform_L[161][0] = l_cell_wire[161];							inform_L[162][0] = l_cell_wire[162];							inform_L[163][0] = l_cell_wire[163];							inform_L[164][0] = l_cell_wire[164];							inform_L[165][0] = l_cell_wire[165];							inform_L[166][0] = l_cell_wire[166];							inform_L[167][0] = l_cell_wire[167];							inform_L[168][0] = l_cell_wire[168];							inform_L[169][0] = l_cell_wire[169];							inform_L[170][0] = l_cell_wire[170];							inform_L[171][0] = l_cell_wire[171];							inform_L[172][0] = l_cell_wire[172];							inform_L[173][0] = l_cell_wire[173];							inform_L[174][0] = l_cell_wire[174];							inform_L[175][0] = l_cell_wire[175];							inform_L[176][0] = l_cell_wire[176];							inform_L[177][0] = l_cell_wire[177];							inform_L[178][0] = l_cell_wire[178];							inform_L[179][0] = l_cell_wire[179];							inform_L[180][0] = l_cell_wire[180];							inform_L[181][0] = l_cell_wire[181];							inform_L[182][0] = l_cell_wire[182];							inform_L[183][0] = l_cell_wire[183];							inform_L[184][0] = l_cell_wire[184];							inform_L[185][0] = l_cell_wire[185];							inform_L[186][0] = l_cell_wire[186];							inform_L[187][0] = l_cell_wire[187];							inform_L[188][0] = l_cell_wire[188];							inform_L[189][0] = l_cell_wire[189];							inform_L[190][0] = l_cell_wire[190];							inform_L[191][0] = l_cell_wire[191];							inform_L[192][0] = l_cell_wire[192];							inform_L[193][0] = l_cell_wire[193];							inform_L[194][0] = l_cell_wire[194];							inform_L[195][0] = l_cell_wire[195];							inform_L[196][0] = l_cell_wire[196];							inform_L[197][0] = l_cell_wire[197];							inform_L[198][0] = l_cell_wire[198];							inform_L[199][0] = l_cell_wire[199];							inform_L[200][0] = l_cell_wire[200];							inform_L[201][0] = l_cell_wire[201];							inform_L[202][0] = l_cell_wire[202];							inform_L[203][0] = l_cell_wire[203];							inform_L[204][0] = l_cell_wire[204];							inform_L[205][0] = l_cell_wire[205];							inform_L[206][0] = l_cell_wire[206];							inform_L[207][0] = l_cell_wire[207];							inform_L[208][0] = l_cell_wire[208];							inform_L[209][0] = l_cell_wire[209];							inform_L[210][0] = l_cell_wire[210];							inform_L[211][0] = l_cell_wire[211];							inform_L[212][0] = l_cell_wire[212];							inform_L[213][0] = l_cell_wire[213];							inform_L[214][0] = l_cell_wire[214];							inform_L[215][0] = l_cell_wire[215];							inform_L[216][0] = l_cell_wire[216];							inform_L[217][0] = l_cell_wire[217];							inform_L[218][0] = l_cell_wire[218];							inform_L[219][0] = l_cell_wire[219];							inform_L[220][0] = l_cell_wire[220];							inform_L[221][0] = l_cell_wire[221];							inform_L[222][0] = l_cell_wire[222];							inform_L[223][0] = l_cell_wire[223];							inform_L[224][0] = l_cell_wire[224];							inform_L[225][0] = l_cell_wire[225];							inform_L[226][0] = l_cell_wire[226];							inform_L[227][0] = l_cell_wire[227];							inform_L[228][0] = l_cell_wire[228];							inform_L[229][0] = l_cell_wire[229];							inform_L[230][0] = l_cell_wire[230];							inform_L[231][0] = l_cell_wire[231];							inform_L[232][0] = l_cell_wire[232];							inform_L[233][0] = l_cell_wire[233];							inform_L[234][0] = l_cell_wire[234];							inform_L[235][0] = l_cell_wire[235];							inform_L[236][0] = l_cell_wire[236];							inform_L[237][0] = l_cell_wire[237];							inform_L[238][0] = l_cell_wire[238];							inform_L[239][0] = l_cell_wire[239];							inform_L[240][0] = l_cell_wire[240];							inform_L[241][0] = l_cell_wire[241];							inform_L[242][0] = l_cell_wire[242];							inform_L[243][0] = l_cell_wire[243];							inform_L[244][0] = l_cell_wire[244];							inform_L[245][0] = l_cell_wire[245];							inform_L[246][0] = l_cell_wire[246];							inform_L[247][0] = l_cell_wire[247];							inform_L[248][0] = l_cell_wire[248];							inform_L[249][0] = l_cell_wire[249];							inform_L[250][0] = l_cell_wire[250];							inform_L[251][0] = l_cell_wire[251];							inform_L[252][0] = l_cell_wire[252];							inform_L[253][0] = l_cell_wire[253];							inform_L[254][0] = l_cell_wire[254];							inform_L[255][0] = l_cell_wire[255];							inform_L[256][0] = l_cell_wire[256];							inform_L[257][0] = l_cell_wire[257];							inform_L[258][0] = l_cell_wire[258];							inform_L[259][0] = l_cell_wire[259];							inform_L[260][0] = l_cell_wire[260];							inform_L[261][0] = l_cell_wire[261];							inform_L[262][0] = l_cell_wire[262];							inform_L[263][0] = l_cell_wire[263];							inform_L[264][0] = l_cell_wire[264];							inform_L[265][0] = l_cell_wire[265];							inform_L[266][0] = l_cell_wire[266];							inform_L[267][0] = l_cell_wire[267];							inform_L[268][0] = l_cell_wire[268];							inform_L[269][0] = l_cell_wire[269];							inform_L[270][0] = l_cell_wire[270];							inform_L[271][0] = l_cell_wire[271];							inform_L[272][0] = l_cell_wire[272];							inform_L[273][0] = l_cell_wire[273];							inform_L[274][0] = l_cell_wire[274];							inform_L[275][0] = l_cell_wire[275];							inform_L[276][0] = l_cell_wire[276];							inform_L[277][0] = l_cell_wire[277];							inform_L[278][0] = l_cell_wire[278];							inform_L[279][0] = l_cell_wire[279];							inform_L[280][0] = l_cell_wire[280];							inform_L[281][0] = l_cell_wire[281];							inform_L[282][0] = l_cell_wire[282];							inform_L[283][0] = l_cell_wire[283];							inform_L[284][0] = l_cell_wire[284];							inform_L[285][0] = l_cell_wire[285];							inform_L[286][0] = l_cell_wire[286];							inform_L[287][0] = l_cell_wire[287];							inform_L[288][0] = l_cell_wire[288];							inform_L[289][0] = l_cell_wire[289];							inform_L[290][0] = l_cell_wire[290];							inform_L[291][0] = l_cell_wire[291];							inform_L[292][0] = l_cell_wire[292];							inform_L[293][0] = l_cell_wire[293];							inform_L[294][0] = l_cell_wire[294];							inform_L[295][0] = l_cell_wire[295];							inform_L[296][0] = l_cell_wire[296];							inform_L[297][0] = l_cell_wire[297];							inform_L[298][0] = l_cell_wire[298];							inform_L[299][0] = l_cell_wire[299];							inform_L[300][0] = l_cell_wire[300];							inform_L[301][0] = l_cell_wire[301];							inform_L[302][0] = l_cell_wire[302];							inform_L[303][0] = l_cell_wire[303];							inform_L[304][0] = l_cell_wire[304];							inform_L[305][0] = l_cell_wire[305];							inform_L[306][0] = l_cell_wire[306];							inform_L[307][0] = l_cell_wire[307];							inform_L[308][0] = l_cell_wire[308];							inform_L[309][0] = l_cell_wire[309];							inform_L[310][0] = l_cell_wire[310];							inform_L[311][0] = l_cell_wire[311];							inform_L[312][0] = l_cell_wire[312];							inform_L[313][0] = l_cell_wire[313];							inform_L[314][0] = l_cell_wire[314];							inform_L[315][0] = l_cell_wire[315];							inform_L[316][0] = l_cell_wire[316];							inform_L[317][0] = l_cell_wire[317];							inform_L[318][0] = l_cell_wire[318];							inform_L[319][0] = l_cell_wire[319];							inform_L[320][0] = l_cell_wire[320];							inform_L[321][0] = l_cell_wire[321];							inform_L[322][0] = l_cell_wire[322];							inform_L[323][0] = l_cell_wire[323];							inform_L[324][0] = l_cell_wire[324];							inform_L[325][0] = l_cell_wire[325];							inform_L[326][0] = l_cell_wire[326];							inform_L[327][0] = l_cell_wire[327];							inform_L[328][0] = l_cell_wire[328];							inform_L[329][0] = l_cell_wire[329];							inform_L[330][0] = l_cell_wire[330];							inform_L[331][0] = l_cell_wire[331];							inform_L[332][0] = l_cell_wire[332];							inform_L[333][0] = l_cell_wire[333];							inform_L[334][0] = l_cell_wire[334];							inform_L[335][0] = l_cell_wire[335];							inform_L[336][0] = l_cell_wire[336];							inform_L[337][0] = l_cell_wire[337];							inform_L[338][0] = l_cell_wire[338];							inform_L[339][0] = l_cell_wire[339];							inform_L[340][0] = l_cell_wire[340];							inform_L[341][0] = l_cell_wire[341];							inform_L[342][0] = l_cell_wire[342];							inform_L[343][0] = l_cell_wire[343];							inform_L[344][0] = l_cell_wire[344];							inform_L[345][0] = l_cell_wire[345];							inform_L[346][0] = l_cell_wire[346];							inform_L[347][0] = l_cell_wire[347];							inform_L[348][0] = l_cell_wire[348];							inform_L[349][0] = l_cell_wire[349];							inform_L[350][0] = l_cell_wire[350];							inform_L[351][0] = l_cell_wire[351];							inform_L[352][0] = l_cell_wire[352];							inform_L[353][0] = l_cell_wire[353];							inform_L[354][0] = l_cell_wire[354];							inform_L[355][0] = l_cell_wire[355];							inform_L[356][0] = l_cell_wire[356];							inform_L[357][0] = l_cell_wire[357];							inform_L[358][0] = l_cell_wire[358];							inform_L[359][0] = l_cell_wire[359];							inform_L[360][0] = l_cell_wire[360];							inform_L[361][0] = l_cell_wire[361];							inform_L[362][0] = l_cell_wire[362];							inform_L[363][0] = l_cell_wire[363];							inform_L[364][0] = l_cell_wire[364];							inform_L[365][0] = l_cell_wire[365];							inform_L[366][0] = l_cell_wire[366];							inform_L[367][0] = l_cell_wire[367];							inform_L[368][0] = l_cell_wire[368];							inform_L[369][0] = l_cell_wire[369];							inform_L[370][0] = l_cell_wire[370];							inform_L[371][0] = l_cell_wire[371];							inform_L[372][0] = l_cell_wire[372];							inform_L[373][0] = l_cell_wire[373];							inform_L[374][0] = l_cell_wire[374];							inform_L[375][0] = l_cell_wire[375];							inform_L[376][0] = l_cell_wire[376];							inform_L[377][0] = l_cell_wire[377];							inform_L[378][0] = l_cell_wire[378];							inform_L[379][0] = l_cell_wire[379];							inform_L[380][0] = l_cell_wire[380];							inform_L[381][0] = l_cell_wire[381];							inform_L[382][0] = l_cell_wire[382];							inform_L[383][0] = l_cell_wire[383];							inform_L[384][0] = l_cell_wire[384];							inform_L[385][0] = l_cell_wire[385];							inform_L[386][0] = l_cell_wire[386];							inform_L[387][0] = l_cell_wire[387];							inform_L[388][0] = l_cell_wire[388];							inform_L[389][0] = l_cell_wire[389];							inform_L[390][0] = l_cell_wire[390];							inform_L[391][0] = l_cell_wire[391];							inform_L[392][0] = l_cell_wire[392];							inform_L[393][0] = l_cell_wire[393];							inform_L[394][0] = l_cell_wire[394];							inform_L[395][0] = l_cell_wire[395];							inform_L[396][0] = l_cell_wire[396];							inform_L[397][0] = l_cell_wire[397];							inform_L[398][0] = l_cell_wire[398];							inform_L[399][0] = l_cell_wire[399];							inform_L[400][0] = l_cell_wire[400];							inform_L[401][0] = l_cell_wire[401];							inform_L[402][0] = l_cell_wire[402];							inform_L[403][0] = l_cell_wire[403];							inform_L[404][0] = l_cell_wire[404];							inform_L[405][0] = l_cell_wire[405];							inform_L[406][0] = l_cell_wire[406];							inform_L[407][0] = l_cell_wire[407];							inform_L[408][0] = l_cell_wire[408];							inform_L[409][0] = l_cell_wire[409];							inform_L[410][0] = l_cell_wire[410];							inform_L[411][0] = l_cell_wire[411];							inform_L[412][0] = l_cell_wire[412];							inform_L[413][0] = l_cell_wire[413];							inform_L[414][0] = l_cell_wire[414];							inform_L[415][0] = l_cell_wire[415];							inform_L[416][0] = l_cell_wire[416];							inform_L[417][0] = l_cell_wire[417];							inform_L[418][0] = l_cell_wire[418];							inform_L[419][0] = l_cell_wire[419];							inform_L[420][0] = l_cell_wire[420];							inform_L[421][0] = l_cell_wire[421];							inform_L[422][0] = l_cell_wire[422];							inform_L[423][0] = l_cell_wire[423];							inform_L[424][0] = l_cell_wire[424];							inform_L[425][0] = l_cell_wire[425];							inform_L[426][0] = l_cell_wire[426];							inform_L[427][0] = l_cell_wire[427];							inform_L[428][0] = l_cell_wire[428];							inform_L[429][0] = l_cell_wire[429];							inform_L[430][0] = l_cell_wire[430];							inform_L[431][0] = l_cell_wire[431];							inform_L[432][0] = l_cell_wire[432];							inform_L[433][0] = l_cell_wire[433];							inform_L[434][0] = l_cell_wire[434];							inform_L[435][0] = l_cell_wire[435];							inform_L[436][0] = l_cell_wire[436];							inform_L[437][0] = l_cell_wire[437];							inform_L[438][0] = l_cell_wire[438];							inform_L[439][0] = l_cell_wire[439];							inform_L[440][0] = l_cell_wire[440];							inform_L[441][0] = l_cell_wire[441];							inform_L[442][0] = l_cell_wire[442];							inform_L[443][0] = l_cell_wire[443];							inform_L[444][0] = l_cell_wire[444];							inform_L[445][0] = l_cell_wire[445];							inform_L[446][0] = l_cell_wire[446];							inform_L[447][0] = l_cell_wire[447];							inform_L[448][0] = l_cell_wire[448];							inform_L[449][0] = l_cell_wire[449];							inform_L[450][0] = l_cell_wire[450];							inform_L[451][0] = l_cell_wire[451];							inform_L[452][0] = l_cell_wire[452];							inform_L[453][0] = l_cell_wire[453];							inform_L[454][0] = l_cell_wire[454];							inform_L[455][0] = l_cell_wire[455];							inform_L[456][0] = l_cell_wire[456];							inform_L[457][0] = l_cell_wire[457];							inform_L[458][0] = l_cell_wire[458];							inform_L[459][0] = l_cell_wire[459];							inform_L[460][0] = l_cell_wire[460];							inform_L[461][0] = l_cell_wire[461];							inform_L[462][0] = l_cell_wire[462];							inform_L[463][0] = l_cell_wire[463];							inform_L[464][0] = l_cell_wire[464];							inform_L[465][0] = l_cell_wire[465];							inform_L[466][0] = l_cell_wire[466];							inform_L[467][0] = l_cell_wire[467];							inform_L[468][0] = l_cell_wire[468];							inform_L[469][0] = l_cell_wire[469];							inform_L[470][0] = l_cell_wire[470];							inform_L[471][0] = l_cell_wire[471];							inform_L[472][0] = l_cell_wire[472];							inform_L[473][0] = l_cell_wire[473];							inform_L[474][0] = l_cell_wire[474];							inform_L[475][0] = l_cell_wire[475];							inform_L[476][0] = l_cell_wire[476];							inform_L[477][0] = l_cell_wire[477];							inform_L[478][0] = l_cell_wire[478];							inform_L[479][0] = l_cell_wire[479];							inform_L[480][0] = l_cell_wire[480];							inform_L[481][0] = l_cell_wire[481];							inform_L[482][0] = l_cell_wire[482];							inform_L[483][0] = l_cell_wire[483];							inform_L[484][0] = l_cell_wire[484];							inform_L[485][0] = l_cell_wire[485];							inform_L[486][0] = l_cell_wire[486];							inform_L[487][0] = l_cell_wire[487];							inform_L[488][0] = l_cell_wire[488];							inform_L[489][0] = l_cell_wire[489];							inform_L[490][0] = l_cell_wire[490];							inform_L[491][0] = l_cell_wire[491];							inform_L[492][0] = l_cell_wire[492];							inform_L[493][0] = l_cell_wire[493];							inform_L[494][0] = l_cell_wire[494];							inform_L[495][0] = l_cell_wire[495];							inform_L[496][0] = l_cell_wire[496];							inform_L[497][0] = l_cell_wire[497];							inform_L[498][0] = l_cell_wire[498];							inform_L[499][0] = l_cell_wire[499];							inform_L[500][0] = l_cell_wire[500];							inform_L[501][0] = l_cell_wire[501];							inform_L[502][0] = l_cell_wire[502];							inform_L[503][0] = l_cell_wire[503];							inform_L[504][0] = l_cell_wire[504];							inform_L[505][0] = l_cell_wire[505];							inform_L[506][0] = l_cell_wire[506];							inform_L[507][0] = l_cell_wire[507];							inform_L[508][0] = l_cell_wire[508];							inform_L[509][0] = l_cell_wire[509];							inform_L[510][0] = l_cell_wire[510];							inform_L[511][0] = l_cell_wire[511];							inform_L[512][0] = l_cell_wire[512];							inform_L[513][0] = l_cell_wire[513];							inform_L[514][0] = l_cell_wire[514];							inform_L[515][0] = l_cell_wire[515];							inform_L[516][0] = l_cell_wire[516];							inform_L[517][0] = l_cell_wire[517];							inform_L[518][0] = l_cell_wire[518];							inform_L[519][0] = l_cell_wire[519];							inform_L[520][0] = l_cell_wire[520];							inform_L[521][0] = l_cell_wire[521];							inform_L[522][0] = l_cell_wire[522];							inform_L[523][0] = l_cell_wire[523];							inform_L[524][0] = l_cell_wire[524];							inform_L[525][0] = l_cell_wire[525];							inform_L[526][0] = l_cell_wire[526];							inform_L[527][0] = l_cell_wire[527];							inform_L[528][0] = l_cell_wire[528];							inform_L[529][0] = l_cell_wire[529];							inform_L[530][0] = l_cell_wire[530];							inform_L[531][0] = l_cell_wire[531];							inform_L[532][0] = l_cell_wire[532];							inform_L[533][0] = l_cell_wire[533];							inform_L[534][0] = l_cell_wire[534];							inform_L[535][0] = l_cell_wire[535];							inform_L[536][0] = l_cell_wire[536];							inform_L[537][0] = l_cell_wire[537];							inform_L[538][0] = l_cell_wire[538];							inform_L[539][0] = l_cell_wire[539];							inform_L[540][0] = l_cell_wire[540];							inform_L[541][0] = l_cell_wire[541];							inform_L[542][0] = l_cell_wire[542];							inform_L[543][0] = l_cell_wire[543];							inform_L[544][0] = l_cell_wire[544];							inform_L[545][0] = l_cell_wire[545];							inform_L[546][0] = l_cell_wire[546];							inform_L[547][0] = l_cell_wire[547];							inform_L[548][0] = l_cell_wire[548];							inform_L[549][0] = l_cell_wire[549];							inform_L[550][0] = l_cell_wire[550];							inform_L[551][0] = l_cell_wire[551];							inform_L[552][0] = l_cell_wire[552];							inform_L[553][0] = l_cell_wire[553];							inform_L[554][0] = l_cell_wire[554];							inform_L[555][0] = l_cell_wire[555];							inform_L[556][0] = l_cell_wire[556];							inform_L[557][0] = l_cell_wire[557];							inform_L[558][0] = l_cell_wire[558];							inform_L[559][0] = l_cell_wire[559];							inform_L[560][0] = l_cell_wire[560];							inform_L[561][0] = l_cell_wire[561];							inform_L[562][0] = l_cell_wire[562];							inform_L[563][0] = l_cell_wire[563];							inform_L[564][0] = l_cell_wire[564];							inform_L[565][0] = l_cell_wire[565];							inform_L[566][0] = l_cell_wire[566];							inform_L[567][0] = l_cell_wire[567];							inform_L[568][0] = l_cell_wire[568];							inform_L[569][0] = l_cell_wire[569];							inform_L[570][0] = l_cell_wire[570];							inform_L[571][0] = l_cell_wire[571];							inform_L[572][0] = l_cell_wire[572];							inform_L[573][0] = l_cell_wire[573];							inform_L[574][0] = l_cell_wire[574];							inform_L[575][0] = l_cell_wire[575];							inform_L[576][0] = l_cell_wire[576];							inform_L[577][0] = l_cell_wire[577];							inform_L[578][0] = l_cell_wire[578];							inform_L[579][0] = l_cell_wire[579];							inform_L[580][0] = l_cell_wire[580];							inform_L[581][0] = l_cell_wire[581];							inform_L[582][0] = l_cell_wire[582];							inform_L[583][0] = l_cell_wire[583];							inform_L[584][0] = l_cell_wire[584];							inform_L[585][0] = l_cell_wire[585];							inform_L[586][0] = l_cell_wire[586];							inform_L[587][0] = l_cell_wire[587];							inform_L[588][0] = l_cell_wire[588];							inform_L[589][0] = l_cell_wire[589];							inform_L[590][0] = l_cell_wire[590];							inform_L[591][0] = l_cell_wire[591];							inform_L[592][0] = l_cell_wire[592];							inform_L[593][0] = l_cell_wire[593];							inform_L[594][0] = l_cell_wire[594];							inform_L[595][0] = l_cell_wire[595];							inform_L[596][0] = l_cell_wire[596];							inform_L[597][0] = l_cell_wire[597];							inform_L[598][0] = l_cell_wire[598];							inform_L[599][0] = l_cell_wire[599];							inform_L[600][0] = l_cell_wire[600];							inform_L[601][0] = l_cell_wire[601];							inform_L[602][0] = l_cell_wire[602];							inform_L[603][0] = l_cell_wire[603];							inform_L[604][0] = l_cell_wire[604];							inform_L[605][0] = l_cell_wire[605];							inform_L[606][0] = l_cell_wire[606];							inform_L[607][0] = l_cell_wire[607];							inform_L[608][0] = l_cell_wire[608];							inform_L[609][0] = l_cell_wire[609];							inform_L[610][0] = l_cell_wire[610];							inform_L[611][0] = l_cell_wire[611];							inform_L[612][0] = l_cell_wire[612];							inform_L[613][0] = l_cell_wire[613];							inform_L[614][0] = l_cell_wire[614];							inform_L[615][0] = l_cell_wire[615];							inform_L[616][0] = l_cell_wire[616];							inform_L[617][0] = l_cell_wire[617];							inform_L[618][0] = l_cell_wire[618];							inform_L[619][0] = l_cell_wire[619];							inform_L[620][0] = l_cell_wire[620];							inform_L[621][0] = l_cell_wire[621];							inform_L[622][0] = l_cell_wire[622];							inform_L[623][0] = l_cell_wire[623];							inform_L[624][0] = l_cell_wire[624];							inform_L[625][0] = l_cell_wire[625];							inform_L[626][0] = l_cell_wire[626];							inform_L[627][0] = l_cell_wire[627];							inform_L[628][0] = l_cell_wire[628];							inform_L[629][0] = l_cell_wire[629];							inform_L[630][0] = l_cell_wire[630];							inform_L[631][0] = l_cell_wire[631];							inform_L[632][0] = l_cell_wire[632];							inform_L[633][0] = l_cell_wire[633];							inform_L[634][0] = l_cell_wire[634];							inform_L[635][0] = l_cell_wire[635];							inform_L[636][0] = l_cell_wire[636];							inform_L[637][0] = l_cell_wire[637];							inform_L[638][0] = l_cell_wire[638];							inform_L[639][0] = l_cell_wire[639];							inform_L[640][0] = l_cell_wire[640];							inform_L[641][0] = l_cell_wire[641];							inform_L[642][0] = l_cell_wire[642];							inform_L[643][0] = l_cell_wire[643];							inform_L[644][0] = l_cell_wire[644];							inform_L[645][0] = l_cell_wire[645];							inform_L[646][0] = l_cell_wire[646];							inform_L[647][0] = l_cell_wire[647];							inform_L[648][0] = l_cell_wire[648];							inform_L[649][0] = l_cell_wire[649];							inform_L[650][0] = l_cell_wire[650];							inform_L[651][0] = l_cell_wire[651];							inform_L[652][0] = l_cell_wire[652];							inform_L[653][0] = l_cell_wire[653];							inform_L[654][0] = l_cell_wire[654];							inform_L[655][0] = l_cell_wire[655];							inform_L[656][0] = l_cell_wire[656];							inform_L[657][0] = l_cell_wire[657];							inform_L[658][0] = l_cell_wire[658];							inform_L[659][0] = l_cell_wire[659];							inform_L[660][0] = l_cell_wire[660];							inform_L[661][0] = l_cell_wire[661];							inform_L[662][0] = l_cell_wire[662];							inform_L[663][0] = l_cell_wire[663];							inform_L[664][0] = l_cell_wire[664];							inform_L[665][0] = l_cell_wire[665];							inform_L[666][0] = l_cell_wire[666];							inform_L[667][0] = l_cell_wire[667];							inform_L[668][0] = l_cell_wire[668];							inform_L[669][0] = l_cell_wire[669];							inform_L[670][0] = l_cell_wire[670];							inform_L[671][0] = l_cell_wire[671];							inform_L[672][0] = l_cell_wire[672];							inform_L[673][0] = l_cell_wire[673];							inform_L[674][0] = l_cell_wire[674];							inform_L[675][0] = l_cell_wire[675];							inform_L[676][0] = l_cell_wire[676];							inform_L[677][0] = l_cell_wire[677];							inform_L[678][0] = l_cell_wire[678];							inform_L[679][0] = l_cell_wire[679];							inform_L[680][0] = l_cell_wire[680];							inform_L[681][0] = l_cell_wire[681];							inform_L[682][0] = l_cell_wire[682];							inform_L[683][0] = l_cell_wire[683];							inform_L[684][0] = l_cell_wire[684];							inform_L[685][0] = l_cell_wire[685];							inform_L[686][0] = l_cell_wire[686];							inform_L[687][0] = l_cell_wire[687];							inform_L[688][0] = l_cell_wire[688];							inform_L[689][0] = l_cell_wire[689];							inform_L[690][0] = l_cell_wire[690];							inform_L[691][0] = l_cell_wire[691];							inform_L[692][0] = l_cell_wire[692];							inform_L[693][0] = l_cell_wire[693];							inform_L[694][0] = l_cell_wire[694];							inform_L[695][0] = l_cell_wire[695];							inform_L[696][0] = l_cell_wire[696];							inform_L[697][0] = l_cell_wire[697];							inform_L[698][0] = l_cell_wire[698];							inform_L[699][0] = l_cell_wire[699];							inform_L[700][0] = l_cell_wire[700];							inform_L[701][0] = l_cell_wire[701];							inform_L[702][0] = l_cell_wire[702];							inform_L[703][0] = l_cell_wire[703];							inform_L[704][0] = l_cell_wire[704];							inform_L[705][0] = l_cell_wire[705];							inform_L[706][0] = l_cell_wire[706];							inform_L[707][0] = l_cell_wire[707];							inform_L[708][0] = l_cell_wire[708];							inform_L[709][0] = l_cell_wire[709];							inform_L[710][0] = l_cell_wire[710];							inform_L[711][0] = l_cell_wire[711];							inform_L[712][0] = l_cell_wire[712];							inform_L[713][0] = l_cell_wire[713];							inform_L[714][0] = l_cell_wire[714];							inform_L[715][0] = l_cell_wire[715];							inform_L[716][0] = l_cell_wire[716];							inform_L[717][0] = l_cell_wire[717];							inform_L[718][0] = l_cell_wire[718];							inform_L[719][0] = l_cell_wire[719];							inform_L[720][0] = l_cell_wire[720];							inform_L[721][0] = l_cell_wire[721];							inform_L[722][0] = l_cell_wire[722];							inform_L[723][0] = l_cell_wire[723];							inform_L[724][0] = l_cell_wire[724];							inform_L[725][0] = l_cell_wire[725];							inform_L[726][0] = l_cell_wire[726];							inform_L[727][0] = l_cell_wire[727];							inform_L[728][0] = l_cell_wire[728];							inform_L[729][0] = l_cell_wire[729];							inform_L[730][0] = l_cell_wire[730];							inform_L[731][0] = l_cell_wire[731];							inform_L[732][0] = l_cell_wire[732];							inform_L[733][0] = l_cell_wire[733];							inform_L[734][0] = l_cell_wire[734];							inform_L[735][0] = l_cell_wire[735];							inform_L[736][0] = l_cell_wire[736];							inform_L[737][0] = l_cell_wire[737];							inform_L[738][0] = l_cell_wire[738];							inform_L[739][0] = l_cell_wire[739];							inform_L[740][0] = l_cell_wire[740];							inform_L[741][0] = l_cell_wire[741];							inform_L[742][0] = l_cell_wire[742];							inform_L[743][0] = l_cell_wire[743];							inform_L[744][0] = l_cell_wire[744];							inform_L[745][0] = l_cell_wire[745];							inform_L[746][0] = l_cell_wire[746];							inform_L[747][0] = l_cell_wire[747];							inform_L[748][0] = l_cell_wire[748];							inform_L[749][0] = l_cell_wire[749];							inform_L[750][0] = l_cell_wire[750];							inform_L[751][0] = l_cell_wire[751];							inform_L[752][0] = l_cell_wire[752];							inform_L[753][0] = l_cell_wire[753];							inform_L[754][0] = l_cell_wire[754];							inform_L[755][0] = l_cell_wire[755];							inform_L[756][0] = l_cell_wire[756];							inform_L[757][0] = l_cell_wire[757];							inform_L[758][0] = l_cell_wire[758];							inform_L[759][0] = l_cell_wire[759];							inform_L[760][0] = l_cell_wire[760];							inform_L[761][0] = l_cell_wire[761];							inform_L[762][0] = l_cell_wire[762];							inform_L[763][0] = l_cell_wire[763];							inform_L[764][0] = l_cell_wire[764];							inform_L[765][0] = l_cell_wire[765];							inform_L[766][0] = l_cell_wire[766];							inform_L[767][0] = l_cell_wire[767];							inform_L[768][0] = l_cell_wire[768];							inform_L[769][0] = l_cell_wire[769];							inform_L[770][0] = l_cell_wire[770];							inform_L[771][0] = l_cell_wire[771];							inform_L[772][0] = l_cell_wire[772];							inform_L[773][0] = l_cell_wire[773];							inform_L[774][0] = l_cell_wire[774];							inform_L[775][0] = l_cell_wire[775];							inform_L[776][0] = l_cell_wire[776];							inform_L[777][0] = l_cell_wire[777];							inform_L[778][0] = l_cell_wire[778];							inform_L[779][0] = l_cell_wire[779];							inform_L[780][0] = l_cell_wire[780];							inform_L[781][0] = l_cell_wire[781];							inform_L[782][0] = l_cell_wire[782];							inform_L[783][0] = l_cell_wire[783];							inform_L[784][0] = l_cell_wire[784];							inform_L[785][0] = l_cell_wire[785];							inform_L[786][0] = l_cell_wire[786];							inform_L[787][0] = l_cell_wire[787];							inform_L[788][0] = l_cell_wire[788];							inform_L[789][0] = l_cell_wire[789];							inform_L[790][0] = l_cell_wire[790];							inform_L[791][0] = l_cell_wire[791];							inform_L[792][0] = l_cell_wire[792];							inform_L[793][0] = l_cell_wire[793];							inform_L[794][0] = l_cell_wire[794];							inform_L[795][0] = l_cell_wire[795];							inform_L[796][0] = l_cell_wire[796];							inform_L[797][0] = l_cell_wire[797];							inform_L[798][0] = l_cell_wire[798];							inform_L[799][0] = l_cell_wire[799];							inform_L[800][0] = l_cell_wire[800];							inform_L[801][0] = l_cell_wire[801];							inform_L[802][0] = l_cell_wire[802];							inform_L[803][0] = l_cell_wire[803];							inform_L[804][0] = l_cell_wire[804];							inform_L[805][0] = l_cell_wire[805];							inform_L[806][0] = l_cell_wire[806];							inform_L[807][0] = l_cell_wire[807];							inform_L[808][0] = l_cell_wire[808];							inform_L[809][0] = l_cell_wire[809];							inform_L[810][0] = l_cell_wire[810];							inform_L[811][0] = l_cell_wire[811];							inform_L[812][0] = l_cell_wire[812];							inform_L[813][0] = l_cell_wire[813];							inform_L[814][0] = l_cell_wire[814];							inform_L[815][0] = l_cell_wire[815];							inform_L[816][0] = l_cell_wire[816];							inform_L[817][0] = l_cell_wire[817];							inform_L[818][0] = l_cell_wire[818];							inform_L[819][0] = l_cell_wire[819];							inform_L[820][0] = l_cell_wire[820];							inform_L[821][0] = l_cell_wire[821];							inform_L[822][0] = l_cell_wire[822];							inform_L[823][0] = l_cell_wire[823];							inform_L[824][0] = l_cell_wire[824];							inform_L[825][0] = l_cell_wire[825];							inform_L[826][0] = l_cell_wire[826];							inform_L[827][0] = l_cell_wire[827];							inform_L[828][0] = l_cell_wire[828];							inform_L[829][0] = l_cell_wire[829];							inform_L[830][0] = l_cell_wire[830];							inform_L[831][0] = l_cell_wire[831];							inform_L[832][0] = l_cell_wire[832];							inform_L[833][0] = l_cell_wire[833];							inform_L[834][0] = l_cell_wire[834];							inform_L[835][0] = l_cell_wire[835];							inform_L[836][0] = l_cell_wire[836];							inform_L[837][0] = l_cell_wire[837];							inform_L[838][0] = l_cell_wire[838];							inform_L[839][0] = l_cell_wire[839];							inform_L[840][0] = l_cell_wire[840];							inform_L[841][0] = l_cell_wire[841];							inform_L[842][0] = l_cell_wire[842];							inform_L[843][0] = l_cell_wire[843];							inform_L[844][0] = l_cell_wire[844];							inform_L[845][0] = l_cell_wire[845];							inform_L[846][0] = l_cell_wire[846];							inform_L[847][0] = l_cell_wire[847];							inform_L[848][0] = l_cell_wire[848];							inform_L[849][0] = l_cell_wire[849];							inform_L[850][0] = l_cell_wire[850];							inform_L[851][0] = l_cell_wire[851];							inform_L[852][0] = l_cell_wire[852];							inform_L[853][0] = l_cell_wire[853];							inform_L[854][0] = l_cell_wire[854];							inform_L[855][0] = l_cell_wire[855];							inform_L[856][0] = l_cell_wire[856];							inform_L[857][0] = l_cell_wire[857];							inform_L[858][0] = l_cell_wire[858];							inform_L[859][0] = l_cell_wire[859];							inform_L[860][0] = l_cell_wire[860];							inform_L[861][0] = l_cell_wire[861];							inform_L[862][0] = l_cell_wire[862];							inform_L[863][0] = l_cell_wire[863];							inform_L[864][0] = l_cell_wire[864];							inform_L[865][0] = l_cell_wire[865];							inform_L[866][0] = l_cell_wire[866];							inform_L[867][0] = l_cell_wire[867];							inform_L[868][0] = l_cell_wire[868];							inform_L[869][0] = l_cell_wire[869];							inform_L[870][0] = l_cell_wire[870];							inform_L[871][0] = l_cell_wire[871];							inform_L[872][0] = l_cell_wire[872];							inform_L[873][0] = l_cell_wire[873];							inform_L[874][0] = l_cell_wire[874];							inform_L[875][0] = l_cell_wire[875];							inform_L[876][0] = l_cell_wire[876];							inform_L[877][0] = l_cell_wire[877];							inform_L[878][0] = l_cell_wire[878];							inform_L[879][0] = l_cell_wire[879];							inform_L[880][0] = l_cell_wire[880];							inform_L[881][0] = l_cell_wire[881];							inform_L[882][0] = l_cell_wire[882];							inform_L[883][0] = l_cell_wire[883];							inform_L[884][0] = l_cell_wire[884];							inform_L[885][0] = l_cell_wire[885];							inform_L[886][0] = l_cell_wire[886];							inform_L[887][0] = l_cell_wire[887];							inform_L[888][0] = l_cell_wire[888];							inform_L[889][0] = l_cell_wire[889];							inform_L[890][0] = l_cell_wire[890];							inform_L[891][0] = l_cell_wire[891];							inform_L[892][0] = l_cell_wire[892];							inform_L[893][0] = l_cell_wire[893];							inform_L[894][0] = l_cell_wire[894];							inform_L[895][0] = l_cell_wire[895];							inform_L[896][0] = l_cell_wire[896];							inform_L[897][0] = l_cell_wire[897];							inform_L[898][0] = l_cell_wire[898];							inform_L[899][0] = l_cell_wire[899];							inform_L[900][0] = l_cell_wire[900];							inform_L[901][0] = l_cell_wire[901];							inform_L[902][0] = l_cell_wire[902];							inform_L[903][0] = l_cell_wire[903];							inform_L[904][0] = l_cell_wire[904];							inform_L[905][0] = l_cell_wire[905];							inform_L[906][0] = l_cell_wire[906];							inform_L[907][0] = l_cell_wire[907];							inform_L[908][0] = l_cell_wire[908];							inform_L[909][0] = l_cell_wire[909];							inform_L[910][0] = l_cell_wire[910];							inform_L[911][0] = l_cell_wire[911];							inform_L[912][0] = l_cell_wire[912];							inform_L[913][0] = l_cell_wire[913];							inform_L[914][0] = l_cell_wire[914];							inform_L[915][0] = l_cell_wire[915];							inform_L[916][0] = l_cell_wire[916];							inform_L[917][0] = l_cell_wire[917];							inform_L[918][0] = l_cell_wire[918];							inform_L[919][0] = l_cell_wire[919];							inform_L[920][0] = l_cell_wire[920];							inform_L[921][0] = l_cell_wire[921];							inform_L[922][0] = l_cell_wire[922];							inform_L[923][0] = l_cell_wire[923];							inform_L[924][0] = l_cell_wire[924];							inform_L[925][0] = l_cell_wire[925];							inform_L[926][0] = l_cell_wire[926];							inform_L[927][0] = l_cell_wire[927];							inform_L[928][0] = l_cell_wire[928];							inform_L[929][0] = l_cell_wire[929];							inform_L[930][0] = l_cell_wire[930];							inform_L[931][0] = l_cell_wire[931];							inform_L[932][0] = l_cell_wire[932];							inform_L[933][0] = l_cell_wire[933];							inform_L[934][0] = l_cell_wire[934];							inform_L[935][0] = l_cell_wire[935];							inform_L[936][0] = l_cell_wire[936];							inform_L[937][0] = l_cell_wire[937];							inform_L[938][0] = l_cell_wire[938];							inform_L[939][0] = l_cell_wire[939];							inform_L[940][0] = l_cell_wire[940];							inform_L[941][0] = l_cell_wire[941];							inform_L[942][0] = l_cell_wire[942];							inform_L[943][0] = l_cell_wire[943];							inform_L[944][0] = l_cell_wire[944];							inform_L[945][0] = l_cell_wire[945];							inform_L[946][0] = l_cell_wire[946];							inform_L[947][0] = l_cell_wire[947];							inform_L[948][0] = l_cell_wire[948];							inform_L[949][0] = l_cell_wire[949];							inform_L[950][0] = l_cell_wire[950];							inform_L[951][0] = l_cell_wire[951];							inform_L[952][0] = l_cell_wire[952];							inform_L[953][0] = l_cell_wire[953];							inform_L[954][0] = l_cell_wire[954];							inform_L[955][0] = l_cell_wire[955];							inform_L[956][0] = l_cell_wire[956];							inform_L[957][0] = l_cell_wire[957];							inform_L[958][0] = l_cell_wire[958];							inform_L[959][0] = l_cell_wire[959];							inform_L[960][0] = l_cell_wire[960];							inform_L[961][0] = l_cell_wire[961];							inform_L[962][0] = l_cell_wire[962];							inform_L[963][0] = l_cell_wire[963];							inform_L[964][0] = l_cell_wire[964];							inform_L[965][0] = l_cell_wire[965];							inform_L[966][0] = l_cell_wire[966];							inform_L[967][0] = l_cell_wire[967];							inform_L[968][0] = l_cell_wire[968];							inform_L[969][0] = l_cell_wire[969];							inform_L[970][0] = l_cell_wire[970];							inform_L[971][0] = l_cell_wire[971];							inform_L[972][0] = l_cell_wire[972];							inform_L[973][0] = l_cell_wire[973];							inform_L[974][0] = l_cell_wire[974];							inform_L[975][0] = l_cell_wire[975];							inform_L[976][0] = l_cell_wire[976];							inform_L[977][0] = l_cell_wire[977];							inform_L[978][0] = l_cell_wire[978];							inform_L[979][0] = l_cell_wire[979];							inform_L[980][0] = l_cell_wire[980];							inform_L[981][0] = l_cell_wire[981];							inform_L[982][0] = l_cell_wire[982];							inform_L[983][0] = l_cell_wire[983];							inform_L[984][0] = l_cell_wire[984];							inform_L[985][0] = l_cell_wire[985];							inform_L[986][0] = l_cell_wire[986];							inform_L[987][0] = l_cell_wire[987];							inform_L[988][0] = l_cell_wire[988];							inform_L[989][0] = l_cell_wire[989];							inform_L[990][0] = l_cell_wire[990];							inform_L[991][0] = l_cell_wire[991];							inform_L[992][0] = l_cell_wire[992];							inform_L[993][0] = l_cell_wire[993];							inform_L[994][0] = l_cell_wire[994];							inform_L[995][0] = l_cell_wire[995];							inform_L[996][0] = l_cell_wire[996];							inform_L[997][0] = l_cell_wire[997];							inform_L[998][0] = l_cell_wire[998];							inform_L[999][0] = l_cell_wire[999];							inform_L[1000][0] = l_cell_wire[1000];							inform_L[1001][0] = l_cell_wire[1001];							inform_L[1002][0] = l_cell_wire[1002];							inform_L[1003][0] = l_cell_wire[1003];							inform_L[1004][0] = l_cell_wire[1004];							inform_L[1005][0] = l_cell_wire[1005];							inform_L[1006][0] = l_cell_wire[1006];							inform_L[1007][0] = l_cell_wire[1007];							inform_L[1008][0] = l_cell_wire[1008];							inform_L[1009][0] = l_cell_wire[1009];							inform_L[1010][0] = l_cell_wire[1010];							inform_L[1011][0] = l_cell_wire[1011];							inform_L[1012][0] = l_cell_wire[1012];							inform_L[1013][0] = l_cell_wire[1013];							inform_L[1014][0] = l_cell_wire[1014];							inform_L[1015][0] = l_cell_wire[1015];							inform_L[1016][0] = l_cell_wire[1016];							inform_L[1017][0] = l_cell_wire[1017];							inform_L[1018][0] = l_cell_wire[1018];							inform_L[1019][0] = l_cell_wire[1019];							inform_L[1020][0] = l_cell_wire[1020];							inform_L[1021][0] = l_cell_wire[1021];							inform_L[1022][0] = l_cell_wire[1022];							inform_L[1023][0] = l_cell_wire[1023];						end
						2:						begin							inform_R[0][2] = r_cell_wire[0];							inform_R[2][2] = r_cell_wire[1];							inform_R[1][2] = r_cell_wire[2];							inform_R[3][2] = r_cell_wire[3];							inform_R[4][2] = r_cell_wire[4];							inform_R[6][2] = r_cell_wire[5];							inform_R[5][2] = r_cell_wire[6];							inform_R[7][2] = r_cell_wire[7];							inform_R[8][2] = r_cell_wire[8];							inform_R[10][2] = r_cell_wire[9];							inform_R[9][2] = r_cell_wire[10];							inform_R[11][2] = r_cell_wire[11];							inform_R[12][2] = r_cell_wire[12];							inform_R[14][2] = r_cell_wire[13];							inform_R[13][2] = r_cell_wire[14];							inform_R[15][2] = r_cell_wire[15];							inform_R[16][2] = r_cell_wire[16];							inform_R[18][2] = r_cell_wire[17];							inform_R[17][2] = r_cell_wire[18];							inform_R[19][2] = r_cell_wire[19];							inform_R[20][2] = r_cell_wire[20];							inform_R[22][2] = r_cell_wire[21];							inform_R[21][2] = r_cell_wire[22];							inform_R[23][2] = r_cell_wire[23];							inform_R[24][2] = r_cell_wire[24];							inform_R[26][2] = r_cell_wire[25];							inform_R[25][2] = r_cell_wire[26];							inform_R[27][2] = r_cell_wire[27];							inform_R[28][2] = r_cell_wire[28];							inform_R[30][2] = r_cell_wire[29];							inform_R[29][2] = r_cell_wire[30];							inform_R[31][2] = r_cell_wire[31];							inform_R[32][2] = r_cell_wire[32];							inform_R[34][2] = r_cell_wire[33];							inform_R[33][2] = r_cell_wire[34];							inform_R[35][2] = r_cell_wire[35];							inform_R[36][2] = r_cell_wire[36];							inform_R[38][2] = r_cell_wire[37];							inform_R[37][2] = r_cell_wire[38];							inform_R[39][2] = r_cell_wire[39];							inform_R[40][2] = r_cell_wire[40];							inform_R[42][2] = r_cell_wire[41];							inform_R[41][2] = r_cell_wire[42];							inform_R[43][2] = r_cell_wire[43];							inform_R[44][2] = r_cell_wire[44];							inform_R[46][2] = r_cell_wire[45];							inform_R[45][2] = r_cell_wire[46];							inform_R[47][2] = r_cell_wire[47];							inform_R[48][2] = r_cell_wire[48];							inform_R[50][2] = r_cell_wire[49];							inform_R[49][2] = r_cell_wire[50];							inform_R[51][2] = r_cell_wire[51];							inform_R[52][2] = r_cell_wire[52];							inform_R[54][2] = r_cell_wire[53];							inform_R[53][2] = r_cell_wire[54];							inform_R[55][2] = r_cell_wire[55];							inform_R[56][2] = r_cell_wire[56];							inform_R[58][2] = r_cell_wire[57];							inform_R[57][2] = r_cell_wire[58];							inform_R[59][2] = r_cell_wire[59];							inform_R[60][2] = r_cell_wire[60];							inform_R[62][2] = r_cell_wire[61];							inform_R[61][2] = r_cell_wire[62];							inform_R[63][2] = r_cell_wire[63];							inform_R[64][2] = r_cell_wire[64];							inform_R[66][2] = r_cell_wire[65];							inform_R[65][2] = r_cell_wire[66];							inform_R[67][2] = r_cell_wire[67];							inform_R[68][2] = r_cell_wire[68];							inform_R[70][2] = r_cell_wire[69];							inform_R[69][2] = r_cell_wire[70];							inform_R[71][2] = r_cell_wire[71];							inform_R[72][2] = r_cell_wire[72];							inform_R[74][2] = r_cell_wire[73];							inform_R[73][2] = r_cell_wire[74];							inform_R[75][2] = r_cell_wire[75];							inform_R[76][2] = r_cell_wire[76];							inform_R[78][2] = r_cell_wire[77];							inform_R[77][2] = r_cell_wire[78];							inform_R[79][2] = r_cell_wire[79];							inform_R[80][2] = r_cell_wire[80];							inform_R[82][2] = r_cell_wire[81];							inform_R[81][2] = r_cell_wire[82];							inform_R[83][2] = r_cell_wire[83];							inform_R[84][2] = r_cell_wire[84];							inform_R[86][2] = r_cell_wire[85];							inform_R[85][2] = r_cell_wire[86];							inform_R[87][2] = r_cell_wire[87];							inform_R[88][2] = r_cell_wire[88];							inform_R[90][2] = r_cell_wire[89];							inform_R[89][2] = r_cell_wire[90];							inform_R[91][2] = r_cell_wire[91];							inform_R[92][2] = r_cell_wire[92];							inform_R[94][2] = r_cell_wire[93];							inform_R[93][2] = r_cell_wire[94];							inform_R[95][2] = r_cell_wire[95];							inform_R[96][2] = r_cell_wire[96];							inform_R[98][2] = r_cell_wire[97];							inform_R[97][2] = r_cell_wire[98];							inform_R[99][2] = r_cell_wire[99];							inform_R[100][2] = r_cell_wire[100];							inform_R[102][2] = r_cell_wire[101];							inform_R[101][2] = r_cell_wire[102];							inform_R[103][2] = r_cell_wire[103];							inform_R[104][2] = r_cell_wire[104];							inform_R[106][2] = r_cell_wire[105];							inform_R[105][2] = r_cell_wire[106];							inform_R[107][2] = r_cell_wire[107];							inform_R[108][2] = r_cell_wire[108];							inform_R[110][2] = r_cell_wire[109];							inform_R[109][2] = r_cell_wire[110];							inform_R[111][2] = r_cell_wire[111];							inform_R[112][2] = r_cell_wire[112];							inform_R[114][2] = r_cell_wire[113];							inform_R[113][2] = r_cell_wire[114];							inform_R[115][2] = r_cell_wire[115];							inform_R[116][2] = r_cell_wire[116];							inform_R[118][2] = r_cell_wire[117];							inform_R[117][2] = r_cell_wire[118];							inform_R[119][2] = r_cell_wire[119];							inform_R[120][2] = r_cell_wire[120];							inform_R[122][2] = r_cell_wire[121];							inform_R[121][2] = r_cell_wire[122];							inform_R[123][2] = r_cell_wire[123];							inform_R[124][2] = r_cell_wire[124];							inform_R[126][2] = r_cell_wire[125];							inform_R[125][2] = r_cell_wire[126];							inform_R[127][2] = r_cell_wire[127];							inform_R[128][2] = r_cell_wire[128];							inform_R[130][2] = r_cell_wire[129];							inform_R[129][2] = r_cell_wire[130];							inform_R[131][2] = r_cell_wire[131];							inform_R[132][2] = r_cell_wire[132];							inform_R[134][2] = r_cell_wire[133];							inform_R[133][2] = r_cell_wire[134];							inform_R[135][2] = r_cell_wire[135];							inform_R[136][2] = r_cell_wire[136];							inform_R[138][2] = r_cell_wire[137];							inform_R[137][2] = r_cell_wire[138];							inform_R[139][2] = r_cell_wire[139];							inform_R[140][2] = r_cell_wire[140];							inform_R[142][2] = r_cell_wire[141];							inform_R[141][2] = r_cell_wire[142];							inform_R[143][2] = r_cell_wire[143];							inform_R[144][2] = r_cell_wire[144];							inform_R[146][2] = r_cell_wire[145];							inform_R[145][2] = r_cell_wire[146];							inform_R[147][2] = r_cell_wire[147];							inform_R[148][2] = r_cell_wire[148];							inform_R[150][2] = r_cell_wire[149];							inform_R[149][2] = r_cell_wire[150];							inform_R[151][2] = r_cell_wire[151];							inform_R[152][2] = r_cell_wire[152];							inform_R[154][2] = r_cell_wire[153];							inform_R[153][2] = r_cell_wire[154];							inform_R[155][2] = r_cell_wire[155];							inform_R[156][2] = r_cell_wire[156];							inform_R[158][2] = r_cell_wire[157];							inform_R[157][2] = r_cell_wire[158];							inform_R[159][2] = r_cell_wire[159];							inform_R[160][2] = r_cell_wire[160];							inform_R[162][2] = r_cell_wire[161];							inform_R[161][2] = r_cell_wire[162];							inform_R[163][2] = r_cell_wire[163];							inform_R[164][2] = r_cell_wire[164];							inform_R[166][2] = r_cell_wire[165];							inform_R[165][2] = r_cell_wire[166];							inform_R[167][2] = r_cell_wire[167];							inform_R[168][2] = r_cell_wire[168];							inform_R[170][2] = r_cell_wire[169];							inform_R[169][2] = r_cell_wire[170];							inform_R[171][2] = r_cell_wire[171];							inform_R[172][2] = r_cell_wire[172];							inform_R[174][2] = r_cell_wire[173];							inform_R[173][2] = r_cell_wire[174];							inform_R[175][2] = r_cell_wire[175];							inform_R[176][2] = r_cell_wire[176];							inform_R[178][2] = r_cell_wire[177];							inform_R[177][2] = r_cell_wire[178];							inform_R[179][2] = r_cell_wire[179];							inform_R[180][2] = r_cell_wire[180];							inform_R[182][2] = r_cell_wire[181];							inform_R[181][2] = r_cell_wire[182];							inform_R[183][2] = r_cell_wire[183];							inform_R[184][2] = r_cell_wire[184];							inform_R[186][2] = r_cell_wire[185];							inform_R[185][2] = r_cell_wire[186];							inform_R[187][2] = r_cell_wire[187];							inform_R[188][2] = r_cell_wire[188];							inform_R[190][2] = r_cell_wire[189];							inform_R[189][2] = r_cell_wire[190];							inform_R[191][2] = r_cell_wire[191];							inform_R[192][2] = r_cell_wire[192];							inform_R[194][2] = r_cell_wire[193];							inform_R[193][2] = r_cell_wire[194];							inform_R[195][2] = r_cell_wire[195];							inform_R[196][2] = r_cell_wire[196];							inform_R[198][2] = r_cell_wire[197];							inform_R[197][2] = r_cell_wire[198];							inform_R[199][2] = r_cell_wire[199];							inform_R[200][2] = r_cell_wire[200];							inform_R[202][2] = r_cell_wire[201];							inform_R[201][2] = r_cell_wire[202];							inform_R[203][2] = r_cell_wire[203];							inform_R[204][2] = r_cell_wire[204];							inform_R[206][2] = r_cell_wire[205];							inform_R[205][2] = r_cell_wire[206];							inform_R[207][2] = r_cell_wire[207];							inform_R[208][2] = r_cell_wire[208];							inform_R[210][2] = r_cell_wire[209];							inform_R[209][2] = r_cell_wire[210];							inform_R[211][2] = r_cell_wire[211];							inform_R[212][2] = r_cell_wire[212];							inform_R[214][2] = r_cell_wire[213];							inform_R[213][2] = r_cell_wire[214];							inform_R[215][2] = r_cell_wire[215];							inform_R[216][2] = r_cell_wire[216];							inform_R[218][2] = r_cell_wire[217];							inform_R[217][2] = r_cell_wire[218];							inform_R[219][2] = r_cell_wire[219];							inform_R[220][2] = r_cell_wire[220];							inform_R[222][2] = r_cell_wire[221];							inform_R[221][2] = r_cell_wire[222];							inform_R[223][2] = r_cell_wire[223];							inform_R[224][2] = r_cell_wire[224];							inform_R[226][2] = r_cell_wire[225];							inform_R[225][2] = r_cell_wire[226];							inform_R[227][2] = r_cell_wire[227];							inform_R[228][2] = r_cell_wire[228];							inform_R[230][2] = r_cell_wire[229];							inform_R[229][2] = r_cell_wire[230];							inform_R[231][2] = r_cell_wire[231];							inform_R[232][2] = r_cell_wire[232];							inform_R[234][2] = r_cell_wire[233];							inform_R[233][2] = r_cell_wire[234];							inform_R[235][2] = r_cell_wire[235];							inform_R[236][2] = r_cell_wire[236];							inform_R[238][2] = r_cell_wire[237];							inform_R[237][2] = r_cell_wire[238];							inform_R[239][2] = r_cell_wire[239];							inform_R[240][2] = r_cell_wire[240];							inform_R[242][2] = r_cell_wire[241];							inform_R[241][2] = r_cell_wire[242];							inform_R[243][2] = r_cell_wire[243];							inform_R[244][2] = r_cell_wire[244];							inform_R[246][2] = r_cell_wire[245];							inform_R[245][2] = r_cell_wire[246];							inform_R[247][2] = r_cell_wire[247];							inform_R[248][2] = r_cell_wire[248];							inform_R[250][2] = r_cell_wire[249];							inform_R[249][2] = r_cell_wire[250];							inform_R[251][2] = r_cell_wire[251];							inform_R[252][2] = r_cell_wire[252];							inform_R[254][2] = r_cell_wire[253];							inform_R[253][2] = r_cell_wire[254];							inform_R[255][2] = r_cell_wire[255];							inform_R[256][2] = r_cell_wire[256];							inform_R[258][2] = r_cell_wire[257];							inform_R[257][2] = r_cell_wire[258];							inform_R[259][2] = r_cell_wire[259];							inform_R[260][2] = r_cell_wire[260];							inform_R[262][2] = r_cell_wire[261];							inform_R[261][2] = r_cell_wire[262];							inform_R[263][2] = r_cell_wire[263];							inform_R[264][2] = r_cell_wire[264];							inform_R[266][2] = r_cell_wire[265];							inform_R[265][2] = r_cell_wire[266];							inform_R[267][2] = r_cell_wire[267];							inform_R[268][2] = r_cell_wire[268];							inform_R[270][2] = r_cell_wire[269];							inform_R[269][2] = r_cell_wire[270];							inform_R[271][2] = r_cell_wire[271];							inform_R[272][2] = r_cell_wire[272];							inform_R[274][2] = r_cell_wire[273];							inform_R[273][2] = r_cell_wire[274];							inform_R[275][2] = r_cell_wire[275];							inform_R[276][2] = r_cell_wire[276];							inform_R[278][2] = r_cell_wire[277];							inform_R[277][2] = r_cell_wire[278];							inform_R[279][2] = r_cell_wire[279];							inform_R[280][2] = r_cell_wire[280];							inform_R[282][2] = r_cell_wire[281];							inform_R[281][2] = r_cell_wire[282];							inform_R[283][2] = r_cell_wire[283];							inform_R[284][2] = r_cell_wire[284];							inform_R[286][2] = r_cell_wire[285];							inform_R[285][2] = r_cell_wire[286];							inform_R[287][2] = r_cell_wire[287];							inform_R[288][2] = r_cell_wire[288];							inform_R[290][2] = r_cell_wire[289];							inform_R[289][2] = r_cell_wire[290];							inform_R[291][2] = r_cell_wire[291];							inform_R[292][2] = r_cell_wire[292];							inform_R[294][2] = r_cell_wire[293];							inform_R[293][2] = r_cell_wire[294];							inform_R[295][2] = r_cell_wire[295];							inform_R[296][2] = r_cell_wire[296];							inform_R[298][2] = r_cell_wire[297];							inform_R[297][2] = r_cell_wire[298];							inform_R[299][2] = r_cell_wire[299];							inform_R[300][2] = r_cell_wire[300];							inform_R[302][2] = r_cell_wire[301];							inform_R[301][2] = r_cell_wire[302];							inform_R[303][2] = r_cell_wire[303];							inform_R[304][2] = r_cell_wire[304];							inform_R[306][2] = r_cell_wire[305];							inform_R[305][2] = r_cell_wire[306];							inform_R[307][2] = r_cell_wire[307];							inform_R[308][2] = r_cell_wire[308];							inform_R[310][2] = r_cell_wire[309];							inform_R[309][2] = r_cell_wire[310];							inform_R[311][2] = r_cell_wire[311];							inform_R[312][2] = r_cell_wire[312];							inform_R[314][2] = r_cell_wire[313];							inform_R[313][2] = r_cell_wire[314];							inform_R[315][2] = r_cell_wire[315];							inform_R[316][2] = r_cell_wire[316];							inform_R[318][2] = r_cell_wire[317];							inform_R[317][2] = r_cell_wire[318];							inform_R[319][2] = r_cell_wire[319];							inform_R[320][2] = r_cell_wire[320];							inform_R[322][2] = r_cell_wire[321];							inform_R[321][2] = r_cell_wire[322];							inform_R[323][2] = r_cell_wire[323];							inform_R[324][2] = r_cell_wire[324];							inform_R[326][2] = r_cell_wire[325];							inform_R[325][2] = r_cell_wire[326];							inform_R[327][2] = r_cell_wire[327];							inform_R[328][2] = r_cell_wire[328];							inform_R[330][2] = r_cell_wire[329];							inform_R[329][2] = r_cell_wire[330];							inform_R[331][2] = r_cell_wire[331];							inform_R[332][2] = r_cell_wire[332];							inform_R[334][2] = r_cell_wire[333];							inform_R[333][2] = r_cell_wire[334];							inform_R[335][2] = r_cell_wire[335];							inform_R[336][2] = r_cell_wire[336];							inform_R[338][2] = r_cell_wire[337];							inform_R[337][2] = r_cell_wire[338];							inform_R[339][2] = r_cell_wire[339];							inform_R[340][2] = r_cell_wire[340];							inform_R[342][2] = r_cell_wire[341];							inform_R[341][2] = r_cell_wire[342];							inform_R[343][2] = r_cell_wire[343];							inform_R[344][2] = r_cell_wire[344];							inform_R[346][2] = r_cell_wire[345];							inform_R[345][2] = r_cell_wire[346];							inform_R[347][2] = r_cell_wire[347];							inform_R[348][2] = r_cell_wire[348];							inform_R[350][2] = r_cell_wire[349];							inform_R[349][2] = r_cell_wire[350];							inform_R[351][2] = r_cell_wire[351];							inform_R[352][2] = r_cell_wire[352];							inform_R[354][2] = r_cell_wire[353];							inform_R[353][2] = r_cell_wire[354];							inform_R[355][2] = r_cell_wire[355];							inform_R[356][2] = r_cell_wire[356];							inform_R[358][2] = r_cell_wire[357];							inform_R[357][2] = r_cell_wire[358];							inform_R[359][2] = r_cell_wire[359];							inform_R[360][2] = r_cell_wire[360];							inform_R[362][2] = r_cell_wire[361];							inform_R[361][2] = r_cell_wire[362];							inform_R[363][2] = r_cell_wire[363];							inform_R[364][2] = r_cell_wire[364];							inform_R[366][2] = r_cell_wire[365];							inform_R[365][2] = r_cell_wire[366];							inform_R[367][2] = r_cell_wire[367];							inform_R[368][2] = r_cell_wire[368];							inform_R[370][2] = r_cell_wire[369];							inform_R[369][2] = r_cell_wire[370];							inform_R[371][2] = r_cell_wire[371];							inform_R[372][2] = r_cell_wire[372];							inform_R[374][2] = r_cell_wire[373];							inform_R[373][2] = r_cell_wire[374];							inform_R[375][2] = r_cell_wire[375];							inform_R[376][2] = r_cell_wire[376];							inform_R[378][2] = r_cell_wire[377];							inform_R[377][2] = r_cell_wire[378];							inform_R[379][2] = r_cell_wire[379];							inform_R[380][2] = r_cell_wire[380];							inform_R[382][2] = r_cell_wire[381];							inform_R[381][2] = r_cell_wire[382];							inform_R[383][2] = r_cell_wire[383];							inform_R[384][2] = r_cell_wire[384];							inform_R[386][2] = r_cell_wire[385];							inform_R[385][2] = r_cell_wire[386];							inform_R[387][2] = r_cell_wire[387];							inform_R[388][2] = r_cell_wire[388];							inform_R[390][2] = r_cell_wire[389];							inform_R[389][2] = r_cell_wire[390];							inform_R[391][2] = r_cell_wire[391];							inform_R[392][2] = r_cell_wire[392];							inform_R[394][2] = r_cell_wire[393];							inform_R[393][2] = r_cell_wire[394];							inform_R[395][2] = r_cell_wire[395];							inform_R[396][2] = r_cell_wire[396];							inform_R[398][2] = r_cell_wire[397];							inform_R[397][2] = r_cell_wire[398];							inform_R[399][2] = r_cell_wire[399];							inform_R[400][2] = r_cell_wire[400];							inform_R[402][2] = r_cell_wire[401];							inform_R[401][2] = r_cell_wire[402];							inform_R[403][2] = r_cell_wire[403];							inform_R[404][2] = r_cell_wire[404];							inform_R[406][2] = r_cell_wire[405];							inform_R[405][2] = r_cell_wire[406];							inform_R[407][2] = r_cell_wire[407];							inform_R[408][2] = r_cell_wire[408];							inform_R[410][2] = r_cell_wire[409];							inform_R[409][2] = r_cell_wire[410];							inform_R[411][2] = r_cell_wire[411];							inform_R[412][2] = r_cell_wire[412];							inform_R[414][2] = r_cell_wire[413];							inform_R[413][2] = r_cell_wire[414];							inform_R[415][2] = r_cell_wire[415];							inform_R[416][2] = r_cell_wire[416];							inform_R[418][2] = r_cell_wire[417];							inform_R[417][2] = r_cell_wire[418];							inform_R[419][2] = r_cell_wire[419];							inform_R[420][2] = r_cell_wire[420];							inform_R[422][2] = r_cell_wire[421];							inform_R[421][2] = r_cell_wire[422];							inform_R[423][2] = r_cell_wire[423];							inform_R[424][2] = r_cell_wire[424];							inform_R[426][2] = r_cell_wire[425];							inform_R[425][2] = r_cell_wire[426];							inform_R[427][2] = r_cell_wire[427];							inform_R[428][2] = r_cell_wire[428];							inform_R[430][2] = r_cell_wire[429];							inform_R[429][2] = r_cell_wire[430];							inform_R[431][2] = r_cell_wire[431];							inform_R[432][2] = r_cell_wire[432];							inform_R[434][2] = r_cell_wire[433];							inform_R[433][2] = r_cell_wire[434];							inform_R[435][2] = r_cell_wire[435];							inform_R[436][2] = r_cell_wire[436];							inform_R[438][2] = r_cell_wire[437];							inform_R[437][2] = r_cell_wire[438];							inform_R[439][2] = r_cell_wire[439];							inform_R[440][2] = r_cell_wire[440];							inform_R[442][2] = r_cell_wire[441];							inform_R[441][2] = r_cell_wire[442];							inform_R[443][2] = r_cell_wire[443];							inform_R[444][2] = r_cell_wire[444];							inform_R[446][2] = r_cell_wire[445];							inform_R[445][2] = r_cell_wire[446];							inform_R[447][2] = r_cell_wire[447];							inform_R[448][2] = r_cell_wire[448];							inform_R[450][2] = r_cell_wire[449];							inform_R[449][2] = r_cell_wire[450];							inform_R[451][2] = r_cell_wire[451];							inform_R[452][2] = r_cell_wire[452];							inform_R[454][2] = r_cell_wire[453];							inform_R[453][2] = r_cell_wire[454];							inform_R[455][2] = r_cell_wire[455];							inform_R[456][2] = r_cell_wire[456];							inform_R[458][2] = r_cell_wire[457];							inform_R[457][2] = r_cell_wire[458];							inform_R[459][2] = r_cell_wire[459];							inform_R[460][2] = r_cell_wire[460];							inform_R[462][2] = r_cell_wire[461];							inform_R[461][2] = r_cell_wire[462];							inform_R[463][2] = r_cell_wire[463];							inform_R[464][2] = r_cell_wire[464];							inform_R[466][2] = r_cell_wire[465];							inform_R[465][2] = r_cell_wire[466];							inform_R[467][2] = r_cell_wire[467];							inform_R[468][2] = r_cell_wire[468];							inform_R[470][2] = r_cell_wire[469];							inform_R[469][2] = r_cell_wire[470];							inform_R[471][2] = r_cell_wire[471];							inform_R[472][2] = r_cell_wire[472];							inform_R[474][2] = r_cell_wire[473];							inform_R[473][2] = r_cell_wire[474];							inform_R[475][2] = r_cell_wire[475];							inform_R[476][2] = r_cell_wire[476];							inform_R[478][2] = r_cell_wire[477];							inform_R[477][2] = r_cell_wire[478];							inform_R[479][2] = r_cell_wire[479];							inform_R[480][2] = r_cell_wire[480];							inform_R[482][2] = r_cell_wire[481];							inform_R[481][2] = r_cell_wire[482];							inform_R[483][2] = r_cell_wire[483];							inform_R[484][2] = r_cell_wire[484];							inform_R[486][2] = r_cell_wire[485];							inform_R[485][2] = r_cell_wire[486];							inform_R[487][2] = r_cell_wire[487];							inform_R[488][2] = r_cell_wire[488];							inform_R[490][2] = r_cell_wire[489];							inform_R[489][2] = r_cell_wire[490];							inform_R[491][2] = r_cell_wire[491];							inform_R[492][2] = r_cell_wire[492];							inform_R[494][2] = r_cell_wire[493];							inform_R[493][2] = r_cell_wire[494];							inform_R[495][2] = r_cell_wire[495];							inform_R[496][2] = r_cell_wire[496];							inform_R[498][2] = r_cell_wire[497];							inform_R[497][2] = r_cell_wire[498];							inform_R[499][2] = r_cell_wire[499];							inform_R[500][2] = r_cell_wire[500];							inform_R[502][2] = r_cell_wire[501];							inform_R[501][2] = r_cell_wire[502];							inform_R[503][2] = r_cell_wire[503];							inform_R[504][2] = r_cell_wire[504];							inform_R[506][2] = r_cell_wire[505];							inform_R[505][2] = r_cell_wire[506];							inform_R[507][2] = r_cell_wire[507];							inform_R[508][2] = r_cell_wire[508];							inform_R[510][2] = r_cell_wire[509];							inform_R[509][2] = r_cell_wire[510];							inform_R[511][2] = r_cell_wire[511];							inform_R[512][2] = r_cell_wire[512];							inform_R[514][2] = r_cell_wire[513];							inform_R[513][2] = r_cell_wire[514];							inform_R[515][2] = r_cell_wire[515];							inform_R[516][2] = r_cell_wire[516];							inform_R[518][2] = r_cell_wire[517];							inform_R[517][2] = r_cell_wire[518];							inform_R[519][2] = r_cell_wire[519];							inform_R[520][2] = r_cell_wire[520];							inform_R[522][2] = r_cell_wire[521];							inform_R[521][2] = r_cell_wire[522];							inform_R[523][2] = r_cell_wire[523];							inform_R[524][2] = r_cell_wire[524];							inform_R[526][2] = r_cell_wire[525];							inform_R[525][2] = r_cell_wire[526];							inform_R[527][2] = r_cell_wire[527];							inform_R[528][2] = r_cell_wire[528];							inform_R[530][2] = r_cell_wire[529];							inform_R[529][2] = r_cell_wire[530];							inform_R[531][2] = r_cell_wire[531];							inform_R[532][2] = r_cell_wire[532];							inform_R[534][2] = r_cell_wire[533];							inform_R[533][2] = r_cell_wire[534];							inform_R[535][2] = r_cell_wire[535];							inform_R[536][2] = r_cell_wire[536];							inform_R[538][2] = r_cell_wire[537];							inform_R[537][2] = r_cell_wire[538];							inform_R[539][2] = r_cell_wire[539];							inform_R[540][2] = r_cell_wire[540];							inform_R[542][2] = r_cell_wire[541];							inform_R[541][2] = r_cell_wire[542];							inform_R[543][2] = r_cell_wire[543];							inform_R[544][2] = r_cell_wire[544];							inform_R[546][2] = r_cell_wire[545];							inform_R[545][2] = r_cell_wire[546];							inform_R[547][2] = r_cell_wire[547];							inform_R[548][2] = r_cell_wire[548];							inform_R[550][2] = r_cell_wire[549];							inform_R[549][2] = r_cell_wire[550];							inform_R[551][2] = r_cell_wire[551];							inform_R[552][2] = r_cell_wire[552];							inform_R[554][2] = r_cell_wire[553];							inform_R[553][2] = r_cell_wire[554];							inform_R[555][2] = r_cell_wire[555];							inform_R[556][2] = r_cell_wire[556];							inform_R[558][2] = r_cell_wire[557];							inform_R[557][2] = r_cell_wire[558];							inform_R[559][2] = r_cell_wire[559];							inform_R[560][2] = r_cell_wire[560];							inform_R[562][2] = r_cell_wire[561];							inform_R[561][2] = r_cell_wire[562];							inform_R[563][2] = r_cell_wire[563];							inform_R[564][2] = r_cell_wire[564];							inform_R[566][2] = r_cell_wire[565];							inform_R[565][2] = r_cell_wire[566];							inform_R[567][2] = r_cell_wire[567];							inform_R[568][2] = r_cell_wire[568];							inform_R[570][2] = r_cell_wire[569];							inform_R[569][2] = r_cell_wire[570];							inform_R[571][2] = r_cell_wire[571];							inform_R[572][2] = r_cell_wire[572];							inform_R[574][2] = r_cell_wire[573];							inform_R[573][2] = r_cell_wire[574];							inform_R[575][2] = r_cell_wire[575];							inform_R[576][2] = r_cell_wire[576];							inform_R[578][2] = r_cell_wire[577];							inform_R[577][2] = r_cell_wire[578];							inform_R[579][2] = r_cell_wire[579];							inform_R[580][2] = r_cell_wire[580];							inform_R[582][2] = r_cell_wire[581];							inform_R[581][2] = r_cell_wire[582];							inform_R[583][2] = r_cell_wire[583];							inform_R[584][2] = r_cell_wire[584];							inform_R[586][2] = r_cell_wire[585];							inform_R[585][2] = r_cell_wire[586];							inform_R[587][2] = r_cell_wire[587];							inform_R[588][2] = r_cell_wire[588];							inform_R[590][2] = r_cell_wire[589];							inform_R[589][2] = r_cell_wire[590];							inform_R[591][2] = r_cell_wire[591];							inform_R[592][2] = r_cell_wire[592];							inform_R[594][2] = r_cell_wire[593];							inform_R[593][2] = r_cell_wire[594];							inform_R[595][2] = r_cell_wire[595];							inform_R[596][2] = r_cell_wire[596];							inform_R[598][2] = r_cell_wire[597];							inform_R[597][2] = r_cell_wire[598];							inform_R[599][2] = r_cell_wire[599];							inform_R[600][2] = r_cell_wire[600];							inform_R[602][2] = r_cell_wire[601];							inform_R[601][2] = r_cell_wire[602];							inform_R[603][2] = r_cell_wire[603];							inform_R[604][2] = r_cell_wire[604];							inform_R[606][2] = r_cell_wire[605];							inform_R[605][2] = r_cell_wire[606];							inform_R[607][2] = r_cell_wire[607];							inform_R[608][2] = r_cell_wire[608];							inform_R[610][2] = r_cell_wire[609];							inform_R[609][2] = r_cell_wire[610];							inform_R[611][2] = r_cell_wire[611];							inform_R[612][2] = r_cell_wire[612];							inform_R[614][2] = r_cell_wire[613];							inform_R[613][2] = r_cell_wire[614];							inform_R[615][2] = r_cell_wire[615];							inform_R[616][2] = r_cell_wire[616];							inform_R[618][2] = r_cell_wire[617];							inform_R[617][2] = r_cell_wire[618];							inform_R[619][2] = r_cell_wire[619];							inform_R[620][2] = r_cell_wire[620];							inform_R[622][2] = r_cell_wire[621];							inform_R[621][2] = r_cell_wire[622];							inform_R[623][2] = r_cell_wire[623];							inform_R[624][2] = r_cell_wire[624];							inform_R[626][2] = r_cell_wire[625];							inform_R[625][2] = r_cell_wire[626];							inform_R[627][2] = r_cell_wire[627];							inform_R[628][2] = r_cell_wire[628];							inform_R[630][2] = r_cell_wire[629];							inform_R[629][2] = r_cell_wire[630];							inform_R[631][2] = r_cell_wire[631];							inform_R[632][2] = r_cell_wire[632];							inform_R[634][2] = r_cell_wire[633];							inform_R[633][2] = r_cell_wire[634];							inform_R[635][2] = r_cell_wire[635];							inform_R[636][2] = r_cell_wire[636];							inform_R[638][2] = r_cell_wire[637];							inform_R[637][2] = r_cell_wire[638];							inform_R[639][2] = r_cell_wire[639];							inform_R[640][2] = r_cell_wire[640];							inform_R[642][2] = r_cell_wire[641];							inform_R[641][2] = r_cell_wire[642];							inform_R[643][2] = r_cell_wire[643];							inform_R[644][2] = r_cell_wire[644];							inform_R[646][2] = r_cell_wire[645];							inform_R[645][2] = r_cell_wire[646];							inform_R[647][2] = r_cell_wire[647];							inform_R[648][2] = r_cell_wire[648];							inform_R[650][2] = r_cell_wire[649];							inform_R[649][2] = r_cell_wire[650];							inform_R[651][2] = r_cell_wire[651];							inform_R[652][2] = r_cell_wire[652];							inform_R[654][2] = r_cell_wire[653];							inform_R[653][2] = r_cell_wire[654];							inform_R[655][2] = r_cell_wire[655];							inform_R[656][2] = r_cell_wire[656];							inform_R[658][2] = r_cell_wire[657];							inform_R[657][2] = r_cell_wire[658];							inform_R[659][2] = r_cell_wire[659];							inform_R[660][2] = r_cell_wire[660];							inform_R[662][2] = r_cell_wire[661];							inform_R[661][2] = r_cell_wire[662];							inform_R[663][2] = r_cell_wire[663];							inform_R[664][2] = r_cell_wire[664];							inform_R[666][2] = r_cell_wire[665];							inform_R[665][2] = r_cell_wire[666];							inform_R[667][2] = r_cell_wire[667];							inform_R[668][2] = r_cell_wire[668];							inform_R[670][2] = r_cell_wire[669];							inform_R[669][2] = r_cell_wire[670];							inform_R[671][2] = r_cell_wire[671];							inform_R[672][2] = r_cell_wire[672];							inform_R[674][2] = r_cell_wire[673];							inform_R[673][2] = r_cell_wire[674];							inform_R[675][2] = r_cell_wire[675];							inform_R[676][2] = r_cell_wire[676];							inform_R[678][2] = r_cell_wire[677];							inform_R[677][2] = r_cell_wire[678];							inform_R[679][2] = r_cell_wire[679];							inform_R[680][2] = r_cell_wire[680];							inform_R[682][2] = r_cell_wire[681];							inform_R[681][2] = r_cell_wire[682];							inform_R[683][2] = r_cell_wire[683];							inform_R[684][2] = r_cell_wire[684];							inform_R[686][2] = r_cell_wire[685];							inform_R[685][2] = r_cell_wire[686];							inform_R[687][2] = r_cell_wire[687];							inform_R[688][2] = r_cell_wire[688];							inform_R[690][2] = r_cell_wire[689];							inform_R[689][2] = r_cell_wire[690];							inform_R[691][2] = r_cell_wire[691];							inform_R[692][2] = r_cell_wire[692];							inform_R[694][2] = r_cell_wire[693];							inform_R[693][2] = r_cell_wire[694];							inform_R[695][2] = r_cell_wire[695];							inform_R[696][2] = r_cell_wire[696];							inform_R[698][2] = r_cell_wire[697];							inform_R[697][2] = r_cell_wire[698];							inform_R[699][2] = r_cell_wire[699];							inform_R[700][2] = r_cell_wire[700];							inform_R[702][2] = r_cell_wire[701];							inform_R[701][2] = r_cell_wire[702];							inform_R[703][2] = r_cell_wire[703];							inform_R[704][2] = r_cell_wire[704];							inform_R[706][2] = r_cell_wire[705];							inform_R[705][2] = r_cell_wire[706];							inform_R[707][2] = r_cell_wire[707];							inform_R[708][2] = r_cell_wire[708];							inform_R[710][2] = r_cell_wire[709];							inform_R[709][2] = r_cell_wire[710];							inform_R[711][2] = r_cell_wire[711];							inform_R[712][2] = r_cell_wire[712];							inform_R[714][2] = r_cell_wire[713];							inform_R[713][2] = r_cell_wire[714];							inform_R[715][2] = r_cell_wire[715];							inform_R[716][2] = r_cell_wire[716];							inform_R[718][2] = r_cell_wire[717];							inform_R[717][2] = r_cell_wire[718];							inform_R[719][2] = r_cell_wire[719];							inform_R[720][2] = r_cell_wire[720];							inform_R[722][2] = r_cell_wire[721];							inform_R[721][2] = r_cell_wire[722];							inform_R[723][2] = r_cell_wire[723];							inform_R[724][2] = r_cell_wire[724];							inform_R[726][2] = r_cell_wire[725];							inform_R[725][2] = r_cell_wire[726];							inform_R[727][2] = r_cell_wire[727];							inform_R[728][2] = r_cell_wire[728];							inform_R[730][2] = r_cell_wire[729];							inform_R[729][2] = r_cell_wire[730];							inform_R[731][2] = r_cell_wire[731];							inform_R[732][2] = r_cell_wire[732];							inform_R[734][2] = r_cell_wire[733];							inform_R[733][2] = r_cell_wire[734];							inform_R[735][2] = r_cell_wire[735];							inform_R[736][2] = r_cell_wire[736];							inform_R[738][2] = r_cell_wire[737];							inform_R[737][2] = r_cell_wire[738];							inform_R[739][2] = r_cell_wire[739];							inform_R[740][2] = r_cell_wire[740];							inform_R[742][2] = r_cell_wire[741];							inform_R[741][2] = r_cell_wire[742];							inform_R[743][2] = r_cell_wire[743];							inform_R[744][2] = r_cell_wire[744];							inform_R[746][2] = r_cell_wire[745];							inform_R[745][2] = r_cell_wire[746];							inform_R[747][2] = r_cell_wire[747];							inform_R[748][2] = r_cell_wire[748];							inform_R[750][2] = r_cell_wire[749];							inform_R[749][2] = r_cell_wire[750];							inform_R[751][2] = r_cell_wire[751];							inform_R[752][2] = r_cell_wire[752];							inform_R[754][2] = r_cell_wire[753];							inform_R[753][2] = r_cell_wire[754];							inform_R[755][2] = r_cell_wire[755];							inform_R[756][2] = r_cell_wire[756];							inform_R[758][2] = r_cell_wire[757];							inform_R[757][2] = r_cell_wire[758];							inform_R[759][2] = r_cell_wire[759];							inform_R[760][2] = r_cell_wire[760];							inform_R[762][2] = r_cell_wire[761];							inform_R[761][2] = r_cell_wire[762];							inform_R[763][2] = r_cell_wire[763];							inform_R[764][2] = r_cell_wire[764];							inform_R[766][2] = r_cell_wire[765];							inform_R[765][2] = r_cell_wire[766];							inform_R[767][2] = r_cell_wire[767];							inform_R[768][2] = r_cell_wire[768];							inform_R[770][2] = r_cell_wire[769];							inform_R[769][2] = r_cell_wire[770];							inform_R[771][2] = r_cell_wire[771];							inform_R[772][2] = r_cell_wire[772];							inform_R[774][2] = r_cell_wire[773];							inform_R[773][2] = r_cell_wire[774];							inform_R[775][2] = r_cell_wire[775];							inform_R[776][2] = r_cell_wire[776];							inform_R[778][2] = r_cell_wire[777];							inform_R[777][2] = r_cell_wire[778];							inform_R[779][2] = r_cell_wire[779];							inform_R[780][2] = r_cell_wire[780];							inform_R[782][2] = r_cell_wire[781];							inform_R[781][2] = r_cell_wire[782];							inform_R[783][2] = r_cell_wire[783];							inform_R[784][2] = r_cell_wire[784];							inform_R[786][2] = r_cell_wire[785];							inform_R[785][2] = r_cell_wire[786];							inform_R[787][2] = r_cell_wire[787];							inform_R[788][2] = r_cell_wire[788];							inform_R[790][2] = r_cell_wire[789];							inform_R[789][2] = r_cell_wire[790];							inform_R[791][2] = r_cell_wire[791];							inform_R[792][2] = r_cell_wire[792];							inform_R[794][2] = r_cell_wire[793];							inform_R[793][2] = r_cell_wire[794];							inform_R[795][2] = r_cell_wire[795];							inform_R[796][2] = r_cell_wire[796];							inform_R[798][2] = r_cell_wire[797];							inform_R[797][2] = r_cell_wire[798];							inform_R[799][2] = r_cell_wire[799];							inform_R[800][2] = r_cell_wire[800];							inform_R[802][2] = r_cell_wire[801];							inform_R[801][2] = r_cell_wire[802];							inform_R[803][2] = r_cell_wire[803];							inform_R[804][2] = r_cell_wire[804];							inform_R[806][2] = r_cell_wire[805];							inform_R[805][2] = r_cell_wire[806];							inform_R[807][2] = r_cell_wire[807];							inform_R[808][2] = r_cell_wire[808];							inform_R[810][2] = r_cell_wire[809];							inform_R[809][2] = r_cell_wire[810];							inform_R[811][2] = r_cell_wire[811];							inform_R[812][2] = r_cell_wire[812];							inform_R[814][2] = r_cell_wire[813];							inform_R[813][2] = r_cell_wire[814];							inform_R[815][2] = r_cell_wire[815];							inform_R[816][2] = r_cell_wire[816];							inform_R[818][2] = r_cell_wire[817];							inform_R[817][2] = r_cell_wire[818];							inform_R[819][2] = r_cell_wire[819];							inform_R[820][2] = r_cell_wire[820];							inform_R[822][2] = r_cell_wire[821];							inform_R[821][2] = r_cell_wire[822];							inform_R[823][2] = r_cell_wire[823];							inform_R[824][2] = r_cell_wire[824];							inform_R[826][2] = r_cell_wire[825];							inform_R[825][2] = r_cell_wire[826];							inform_R[827][2] = r_cell_wire[827];							inform_R[828][2] = r_cell_wire[828];							inform_R[830][2] = r_cell_wire[829];							inform_R[829][2] = r_cell_wire[830];							inform_R[831][2] = r_cell_wire[831];							inform_R[832][2] = r_cell_wire[832];							inform_R[834][2] = r_cell_wire[833];							inform_R[833][2] = r_cell_wire[834];							inform_R[835][2] = r_cell_wire[835];							inform_R[836][2] = r_cell_wire[836];							inform_R[838][2] = r_cell_wire[837];							inform_R[837][2] = r_cell_wire[838];							inform_R[839][2] = r_cell_wire[839];							inform_R[840][2] = r_cell_wire[840];							inform_R[842][2] = r_cell_wire[841];							inform_R[841][2] = r_cell_wire[842];							inform_R[843][2] = r_cell_wire[843];							inform_R[844][2] = r_cell_wire[844];							inform_R[846][2] = r_cell_wire[845];							inform_R[845][2] = r_cell_wire[846];							inform_R[847][2] = r_cell_wire[847];							inform_R[848][2] = r_cell_wire[848];							inform_R[850][2] = r_cell_wire[849];							inform_R[849][2] = r_cell_wire[850];							inform_R[851][2] = r_cell_wire[851];							inform_R[852][2] = r_cell_wire[852];							inform_R[854][2] = r_cell_wire[853];							inform_R[853][2] = r_cell_wire[854];							inform_R[855][2] = r_cell_wire[855];							inform_R[856][2] = r_cell_wire[856];							inform_R[858][2] = r_cell_wire[857];							inform_R[857][2] = r_cell_wire[858];							inform_R[859][2] = r_cell_wire[859];							inform_R[860][2] = r_cell_wire[860];							inform_R[862][2] = r_cell_wire[861];							inform_R[861][2] = r_cell_wire[862];							inform_R[863][2] = r_cell_wire[863];							inform_R[864][2] = r_cell_wire[864];							inform_R[866][2] = r_cell_wire[865];							inform_R[865][2] = r_cell_wire[866];							inform_R[867][2] = r_cell_wire[867];							inform_R[868][2] = r_cell_wire[868];							inform_R[870][2] = r_cell_wire[869];							inform_R[869][2] = r_cell_wire[870];							inform_R[871][2] = r_cell_wire[871];							inform_R[872][2] = r_cell_wire[872];							inform_R[874][2] = r_cell_wire[873];							inform_R[873][2] = r_cell_wire[874];							inform_R[875][2] = r_cell_wire[875];							inform_R[876][2] = r_cell_wire[876];							inform_R[878][2] = r_cell_wire[877];							inform_R[877][2] = r_cell_wire[878];							inform_R[879][2] = r_cell_wire[879];							inform_R[880][2] = r_cell_wire[880];							inform_R[882][2] = r_cell_wire[881];							inform_R[881][2] = r_cell_wire[882];							inform_R[883][2] = r_cell_wire[883];							inform_R[884][2] = r_cell_wire[884];							inform_R[886][2] = r_cell_wire[885];							inform_R[885][2] = r_cell_wire[886];							inform_R[887][2] = r_cell_wire[887];							inform_R[888][2] = r_cell_wire[888];							inform_R[890][2] = r_cell_wire[889];							inform_R[889][2] = r_cell_wire[890];							inform_R[891][2] = r_cell_wire[891];							inform_R[892][2] = r_cell_wire[892];							inform_R[894][2] = r_cell_wire[893];							inform_R[893][2] = r_cell_wire[894];							inform_R[895][2] = r_cell_wire[895];							inform_R[896][2] = r_cell_wire[896];							inform_R[898][2] = r_cell_wire[897];							inform_R[897][2] = r_cell_wire[898];							inform_R[899][2] = r_cell_wire[899];							inform_R[900][2] = r_cell_wire[900];							inform_R[902][2] = r_cell_wire[901];							inform_R[901][2] = r_cell_wire[902];							inform_R[903][2] = r_cell_wire[903];							inform_R[904][2] = r_cell_wire[904];							inform_R[906][2] = r_cell_wire[905];							inform_R[905][2] = r_cell_wire[906];							inform_R[907][2] = r_cell_wire[907];							inform_R[908][2] = r_cell_wire[908];							inform_R[910][2] = r_cell_wire[909];							inform_R[909][2] = r_cell_wire[910];							inform_R[911][2] = r_cell_wire[911];							inform_R[912][2] = r_cell_wire[912];							inform_R[914][2] = r_cell_wire[913];							inform_R[913][2] = r_cell_wire[914];							inform_R[915][2] = r_cell_wire[915];							inform_R[916][2] = r_cell_wire[916];							inform_R[918][2] = r_cell_wire[917];							inform_R[917][2] = r_cell_wire[918];							inform_R[919][2] = r_cell_wire[919];							inform_R[920][2] = r_cell_wire[920];							inform_R[922][2] = r_cell_wire[921];							inform_R[921][2] = r_cell_wire[922];							inform_R[923][2] = r_cell_wire[923];							inform_R[924][2] = r_cell_wire[924];							inform_R[926][2] = r_cell_wire[925];							inform_R[925][2] = r_cell_wire[926];							inform_R[927][2] = r_cell_wire[927];							inform_R[928][2] = r_cell_wire[928];							inform_R[930][2] = r_cell_wire[929];							inform_R[929][2] = r_cell_wire[930];							inform_R[931][2] = r_cell_wire[931];							inform_R[932][2] = r_cell_wire[932];							inform_R[934][2] = r_cell_wire[933];							inform_R[933][2] = r_cell_wire[934];							inform_R[935][2] = r_cell_wire[935];							inform_R[936][2] = r_cell_wire[936];							inform_R[938][2] = r_cell_wire[937];							inform_R[937][2] = r_cell_wire[938];							inform_R[939][2] = r_cell_wire[939];							inform_R[940][2] = r_cell_wire[940];							inform_R[942][2] = r_cell_wire[941];							inform_R[941][2] = r_cell_wire[942];							inform_R[943][2] = r_cell_wire[943];							inform_R[944][2] = r_cell_wire[944];							inform_R[946][2] = r_cell_wire[945];							inform_R[945][2] = r_cell_wire[946];							inform_R[947][2] = r_cell_wire[947];							inform_R[948][2] = r_cell_wire[948];							inform_R[950][2] = r_cell_wire[949];							inform_R[949][2] = r_cell_wire[950];							inform_R[951][2] = r_cell_wire[951];							inform_R[952][2] = r_cell_wire[952];							inform_R[954][2] = r_cell_wire[953];							inform_R[953][2] = r_cell_wire[954];							inform_R[955][2] = r_cell_wire[955];							inform_R[956][2] = r_cell_wire[956];							inform_R[958][2] = r_cell_wire[957];							inform_R[957][2] = r_cell_wire[958];							inform_R[959][2] = r_cell_wire[959];							inform_R[960][2] = r_cell_wire[960];							inform_R[962][2] = r_cell_wire[961];							inform_R[961][2] = r_cell_wire[962];							inform_R[963][2] = r_cell_wire[963];							inform_R[964][2] = r_cell_wire[964];							inform_R[966][2] = r_cell_wire[965];							inform_R[965][2] = r_cell_wire[966];							inform_R[967][2] = r_cell_wire[967];							inform_R[968][2] = r_cell_wire[968];							inform_R[970][2] = r_cell_wire[969];							inform_R[969][2] = r_cell_wire[970];							inform_R[971][2] = r_cell_wire[971];							inform_R[972][2] = r_cell_wire[972];							inform_R[974][2] = r_cell_wire[973];							inform_R[973][2] = r_cell_wire[974];							inform_R[975][2] = r_cell_wire[975];							inform_R[976][2] = r_cell_wire[976];							inform_R[978][2] = r_cell_wire[977];							inform_R[977][2] = r_cell_wire[978];							inform_R[979][2] = r_cell_wire[979];							inform_R[980][2] = r_cell_wire[980];							inform_R[982][2] = r_cell_wire[981];							inform_R[981][2] = r_cell_wire[982];							inform_R[983][2] = r_cell_wire[983];							inform_R[984][2] = r_cell_wire[984];							inform_R[986][2] = r_cell_wire[985];							inform_R[985][2] = r_cell_wire[986];							inform_R[987][2] = r_cell_wire[987];							inform_R[988][2] = r_cell_wire[988];							inform_R[990][2] = r_cell_wire[989];							inform_R[989][2] = r_cell_wire[990];							inform_R[991][2] = r_cell_wire[991];							inform_R[992][2] = r_cell_wire[992];							inform_R[994][2] = r_cell_wire[993];							inform_R[993][2] = r_cell_wire[994];							inform_R[995][2] = r_cell_wire[995];							inform_R[996][2] = r_cell_wire[996];							inform_R[998][2] = r_cell_wire[997];							inform_R[997][2] = r_cell_wire[998];							inform_R[999][2] = r_cell_wire[999];							inform_R[1000][2] = r_cell_wire[1000];							inform_R[1002][2] = r_cell_wire[1001];							inform_R[1001][2] = r_cell_wire[1002];							inform_R[1003][2] = r_cell_wire[1003];							inform_R[1004][2] = r_cell_wire[1004];							inform_R[1006][2] = r_cell_wire[1005];							inform_R[1005][2] = r_cell_wire[1006];							inform_R[1007][2] = r_cell_wire[1007];							inform_R[1008][2] = r_cell_wire[1008];							inform_R[1010][2] = r_cell_wire[1009];							inform_R[1009][2] = r_cell_wire[1010];							inform_R[1011][2] = r_cell_wire[1011];							inform_R[1012][2] = r_cell_wire[1012];							inform_R[1014][2] = r_cell_wire[1013];							inform_R[1013][2] = r_cell_wire[1014];							inform_R[1015][2] = r_cell_wire[1015];							inform_R[1016][2] = r_cell_wire[1016];							inform_R[1018][2] = r_cell_wire[1017];							inform_R[1017][2] = r_cell_wire[1018];							inform_R[1019][2] = r_cell_wire[1019];							inform_R[1020][2] = r_cell_wire[1020];							inform_R[1022][2] = r_cell_wire[1021];							inform_R[1021][2] = r_cell_wire[1022];							inform_R[1023][2] = r_cell_wire[1023];							inform_L[0][1] = l_cell_wire[0];							inform_L[2][1] = l_cell_wire[1];							inform_L[1][1] = l_cell_wire[2];							inform_L[3][1] = l_cell_wire[3];							inform_L[4][1] = l_cell_wire[4];							inform_L[6][1] = l_cell_wire[5];							inform_L[5][1] = l_cell_wire[6];							inform_L[7][1] = l_cell_wire[7];							inform_L[8][1] = l_cell_wire[8];							inform_L[10][1] = l_cell_wire[9];							inform_L[9][1] = l_cell_wire[10];							inform_L[11][1] = l_cell_wire[11];							inform_L[12][1] = l_cell_wire[12];							inform_L[14][1] = l_cell_wire[13];							inform_L[13][1] = l_cell_wire[14];							inform_L[15][1] = l_cell_wire[15];							inform_L[16][1] = l_cell_wire[16];							inform_L[18][1] = l_cell_wire[17];							inform_L[17][1] = l_cell_wire[18];							inform_L[19][1] = l_cell_wire[19];							inform_L[20][1] = l_cell_wire[20];							inform_L[22][1] = l_cell_wire[21];							inform_L[21][1] = l_cell_wire[22];							inform_L[23][1] = l_cell_wire[23];							inform_L[24][1] = l_cell_wire[24];							inform_L[26][1] = l_cell_wire[25];							inform_L[25][1] = l_cell_wire[26];							inform_L[27][1] = l_cell_wire[27];							inform_L[28][1] = l_cell_wire[28];							inform_L[30][1] = l_cell_wire[29];							inform_L[29][1] = l_cell_wire[30];							inform_L[31][1] = l_cell_wire[31];							inform_L[32][1] = l_cell_wire[32];							inform_L[34][1] = l_cell_wire[33];							inform_L[33][1] = l_cell_wire[34];							inform_L[35][1] = l_cell_wire[35];							inform_L[36][1] = l_cell_wire[36];							inform_L[38][1] = l_cell_wire[37];							inform_L[37][1] = l_cell_wire[38];							inform_L[39][1] = l_cell_wire[39];							inform_L[40][1] = l_cell_wire[40];							inform_L[42][1] = l_cell_wire[41];							inform_L[41][1] = l_cell_wire[42];							inform_L[43][1] = l_cell_wire[43];							inform_L[44][1] = l_cell_wire[44];							inform_L[46][1] = l_cell_wire[45];							inform_L[45][1] = l_cell_wire[46];							inform_L[47][1] = l_cell_wire[47];							inform_L[48][1] = l_cell_wire[48];							inform_L[50][1] = l_cell_wire[49];							inform_L[49][1] = l_cell_wire[50];							inform_L[51][1] = l_cell_wire[51];							inform_L[52][1] = l_cell_wire[52];							inform_L[54][1] = l_cell_wire[53];							inform_L[53][1] = l_cell_wire[54];							inform_L[55][1] = l_cell_wire[55];							inform_L[56][1] = l_cell_wire[56];							inform_L[58][1] = l_cell_wire[57];							inform_L[57][1] = l_cell_wire[58];							inform_L[59][1] = l_cell_wire[59];							inform_L[60][1] = l_cell_wire[60];							inform_L[62][1] = l_cell_wire[61];							inform_L[61][1] = l_cell_wire[62];							inform_L[63][1] = l_cell_wire[63];							inform_L[64][1] = l_cell_wire[64];							inform_L[66][1] = l_cell_wire[65];							inform_L[65][1] = l_cell_wire[66];							inform_L[67][1] = l_cell_wire[67];							inform_L[68][1] = l_cell_wire[68];							inform_L[70][1] = l_cell_wire[69];							inform_L[69][1] = l_cell_wire[70];							inform_L[71][1] = l_cell_wire[71];							inform_L[72][1] = l_cell_wire[72];							inform_L[74][1] = l_cell_wire[73];							inform_L[73][1] = l_cell_wire[74];							inform_L[75][1] = l_cell_wire[75];							inform_L[76][1] = l_cell_wire[76];							inform_L[78][1] = l_cell_wire[77];							inform_L[77][1] = l_cell_wire[78];							inform_L[79][1] = l_cell_wire[79];							inform_L[80][1] = l_cell_wire[80];							inform_L[82][1] = l_cell_wire[81];							inform_L[81][1] = l_cell_wire[82];							inform_L[83][1] = l_cell_wire[83];							inform_L[84][1] = l_cell_wire[84];							inform_L[86][1] = l_cell_wire[85];							inform_L[85][1] = l_cell_wire[86];							inform_L[87][1] = l_cell_wire[87];							inform_L[88][1] = l_cell_wire[88];							inform_L[90][1] = l_cell_wire[89];							inform_L[89][1] = l_cell_wire[90];							inform_L[91][1] = l_cell_wire[91];							inform_L[92][1] = l_cell_wire[92];							inform_L[94][1] = l_cell_wire[93];							inform_L[93][1] = l_cell_wire[94];							inform_L[95][1] = l_cell_wire[95];							inform_L[96][1] = l_cell_wire[96];							inform_L[98][1] = l_cell_wire[97];							inform_L[97][1] = l_cell_wire[98];							inform_L[99][1] = l_cell_wire[99];							inform_L[100][1] = l_cell_wire[100];							inform_L[102][1] = l_cell_wire[101];							inform_L[101][1] = l_cell_wire[102];							inform_L[103][1] = l_cell_wire[103];							inform_L[104][1] = l_cell_wire[104];							inform_L[106][1] = l_cell_wire[105];							inform_L[105][1] = l_cell_wire[106];							inform_L[107][1] = l_cell_wire[107];							inform_L[108][1] = l_cell_wire[108];							inform_L[110][1] = l_cell_wire[109];							inform_L[109][1] = l_cell_wire[110];							inform_L[111][1] = l_cell_wire[111];							inform_L[112][1] = l_cell_wire[112];							inform_L[114][1] = l_cell_wire[113];							inform_L[113][1] = l_cell_wire[114];							inform_L[115][1] = l_cell_wire[115];							inform_L[116][1] = l_cell_wire[116];							inform_L[118][1] = l_cell_wire[117];							inform_L[117][1] = l_cell_wire[118];							inform_L[119][1] = l_cell_wire[119];							inform_L[120][1] = l_cell_wire[120];							inform_L[122][1] = l_cell_wire[121];							inform_L[121][1] = l_cell_wire[122];							inform_L[123][1] = l_cell_wire[123];							inform_L[124][1] = l_cell_wire[124];							inform_L[126][1] = l_cell_wire[125];							inform_L[125][1] = l_cell_wire[126];							inform_L[127][1] = l_cell_wire[127];							inform_L[128][1] = l_cell_wire[128];							inform_L[130][1] = l_cell_wire[129];							inform_L[129][1] = l_cell_wire[130];							inform_L[131][1] = l_cell_wire[131];							inform_L[132][1] = l_cell_wire[132];							inform_L[134][1] = l_cell_wire[133];							inform_L[133][1] = l_cell_wire[134];							inform_L[135][1] = l_cell_wire[135];							inform_L[136][1] = l_cell_wire[136];							inform_L[138][1] = l_cell_wire[137];							inform_L[137][1] = l_cell_wire[138];							inform_L[139][1] = l_cell_wire[139];							inform_L[140][1] = l_cell_wire[140];							inform_L[142][1] = l_cell_wire[141];							inform_L[141][1] = l_cell_wire[142];							inform_L[143][1] = l_cell_wire[143];							inform_L[144][1] = l_cell_wire[144];							inform_L[146][1] = l_cell_wire[145];							inform_L[145][1] = l_cell_wire[146];							inform_L[147][1] = l_cell_wire[147];							inform_L[148][1] = l_cell_wire[148];							inform_L[150][1] = l_cell_wire[149];							inform_L[149][1] = l_cell_wire[150];							inform_L[151][1] = l_cell_wire[151];							inform_L[152][1] = l_cell_wire[152];							inform_L[154][1] = l_cell_wire[153];							inform_L[153][1] = l_cell_wire[154];							inform_L[155][1] = l_cell_wire[155];							inform_L[156][1] = l_cell_wire[156];							inform_L[158][1] = l_cell_wire[157];							inform_L[157][1] = l_cell_wire[158];							inform_L[159][1] = l_cell_wire[159];							inform_L[160][1] = l_cell_wire[160];							inform_L[162][1] = l_cell_wire[161];							inform_L[161][1] = l_cell_wire[162];							inform_L[163][1] = l_cell_wire[163];							inform_L[164][1] = l_cell_wire[164];							inform_L[166][1] = l_cell_wire[165];							inform_L[165][1] = l_cell_wire[166];							inform_L[167][1] = l_cell_wire[167];							inform_L[168][1] = l_cell_wire[168];							inform_L[170][1] = l_cell_wire[169];							inform_L[169][1] = l_cell_wire[170];							inform_L[171][1] = l_cell_wire[171];							inform_L[172][1] = l_cell_wire[172];							inform_L[174][1] = l_cell_wire[173];							inform_L[173][1] = l_cell_wire[174];							inform_L[175][1] = l_cell_wire[175];							inform_L[176][1] = l_cell_wire[176];							inform_L[178][1] = l_cell_wire[177];							inform_L[177][1] = l_cell_wire[178];							inform_L[179][1] = l_cell_wire[179];							inform_L[180][1] = l_cell_wire[180];							inform_L[182][1] = l_cell_wire[181];							inform_L[181][1] = l_cell_wire[182];							inform_L[183][1] = l_cell_wire[183];							inform_L[184][1] = l_cell_wire[184];							inform_L[186][1] = l_cell_wire[185];							inform_L[185][1] = l_cell_wire[186];							inform_L[187][1] = l_cell_wire[187];							inform_L[188][1] = l_cell_wire[188];							inform_L[190][1] = l_cell_wire[189];							inform_L[189][1] = l_cell_wire[190];							inform_L[191][1] = l_cell_wire[191];							inform_L[192][1] = l_cell_wire[192];							inform_L[194][1] = l_cell_wire[193];							inform_L[193][1] = l_cell_wire[194];							inform_L[195][1] = l_cell_wire[195];							inform_L[196][1] = l_cell_wire[196];							inform_L[198][1] = l_cell_wire[197];							inform_L[197][1] = l_cell_wire[198];							inform_L[199][1] = l_cell_wire[199];							inform_L[200][1] = l_cell_wire[200];							inform_L[202][1] = l_cell_wire[201];							inform_L[201][1] = l_cell_wire[202];							inform_L[203][1] = l_cell_wire[203];							inform_L[204][1] = l_cell_wire[204];							inform_L[206][1] = l_cell_wire[205];							inform_L[205][1] = l_cell_wire[206];							inform_L[207][1] = l_cell_wire[207];							inform_L[208][1] = l_cell_wire[208];							inform_L[210][1] = l_cell_wire[209];							inform_L[209][1] = l_cell_wire[210];							inform_L[211][1] = l_cell_wire[211];							inform_L[212][1] = l_cell_wire[212];							inform_L[214][1] = l_cell_wire[213];							inform_L[213][1] = l_cell_wire[214];							inform_L[215][1] = l_cell_wire[215];							inform_L[216][1] = l_cell_wire[216];							inform_L[218][1] = l_cell_wire[217];							inform_L[217][1] = l_cell_wire[218];							inform_L[219][1] = l_cell_wire[219];							inform_L[220][1] = l_cell_wire[220];							inform_L[222][1] = l_cell_wire[221];							inform_L[221][1] = l_cell_wire[222];							inform_L[223][1] = l_cell_wire[223];							inform_L[224][1] = l_cell_wire[224];							inform_L[226][1] = l_cell_wire[225];							inform_L[225][1] = l_cell_wire[226];							inform_L[227][1] = l_cell_wire[227];							inform_L[228][1] = l_cell_wire[228];							inform_L[230][1] = l_cell_wire[229];							inform_L[229][1] = l_cell_wire[230];							inform_L[231][1] = l_cell_wire[231];							inform_L[232][1] = l_cell_wire[232];							inform_L[234][1] = l_cell_wire[233];							inform_L[233][1] = l_cell_wire[234];							inform_L[235][1] = l_cell_wire[235];							inform_L[236][1] = l_cell_wire[236];							inform_L[238][1] = l_cell_wire[237];							inform_L[237][1] = l_cell_wire[238];							inform_L[239][1] = l_cell_wire[239];							inform_L[240][1] = l_cell_wire[240];							inform_L[242][1] = l_cell_wire[241];							inform_L[241][1] = l_cell_wire[242];							inform_L[243][1] = l_cell_wire[243];							inform_L[244][1] = l_cell_wire[244];							inform_L[246][1] = l_cell_wire[245];							inform_L[245][1] = l_cell_wire[246];							inform_L[247][1] = l_cell_wire[247];							inform_L[248][1] = l_cell_wire[248];							inform_L[250][1] = l_cell_wire[249];							inform_L[249][1] = l_cell_wire[250];							inform_L[251][1] = l_cell_wire[251];							inform_L[252][1] = l_cell_wire[252];							inform_L[254][1] = l_cell_wire[253];							inform_L[253][1] = l_cell_wire[254];							inform_L[255][1] = l_cell_wire[255];							inform_L[256][1] = l_cell_wire[256];							inform_L[258][1] = l_cell_wire[257];							inform_L[257][1] = l_cell_wire[258];							inform_L[259][1] = l_cell_wire[259];							inform_L[260][1] = l_cell_wire[260];							inform_L[262][1] = l_cell_wire[261];							inform_L[261][1] = l_cell_wire[262];							inform_L[263][1] = l_cell_wire[263];							inform_L[264][1] = l_cell_wire[264];							inform_L[266][1] = l_cell_wire[265];							inform_L[265][1] = l_cell_wire[266];							inform_L[267][1] = l_cell_wire[267];							inform_L[268][1] = l_cell_wire[268];							inform_L[270][1] = l_cell_wire[269];							inform_L[269][1] = l_cell_wire[270];							inform_L[271][1] = l_cell_wire[271];							inform_L[272][1] = l_cell_wire[272];							inform_L[274][1] = l_cell_wire[273];							inform_L[273][1] = l_cell_wire[274];							inform_L[275][1] = l_cell_wire[275];							inform_L[276][1] = l_cell_wire[276];							inform_L[278][1] = l_cell_wire[277];							inform_L[277][1] = l_cell_wire[278];							inform_L[279][1] = l_cell_wire[279];							inform_L[280][1] = l_cell_wire[280];							inform_L[282][1] = l_cell_wire[281];							inform_L[281][1] = l_cell_wire[282];							inform_L[283][1] = l_cell_wire[283];							inform_L[284][1] = l_cell_wire[284];							inform_L[286][1] = l_cell_wire[285];							inform_L[285][1] = l_cell_wire[286];							inform_L[287][1] = l_cell_wire[287];							inform_L[288][1] = l_cell_wire[288];							inform_L[290][1] = l_cell_wire[289];							inform_L[289][1] = l_cell_wire[290];							inform_L[291][1] = l_cell_wire[291];							inform_L[292][1] = l_cell_wire[292];							inform_L[294][1] = l_cell_wire[293];							inform_L[293][1] = l_cell_wire[294];							inform_L[295][1] = l_cell_wire[295];							inform_L[296][1] = l_cell_wire[296];							inform_L[298][1] = l_cell_wire[297];							inform_L[297][1] = l_cell_wire[298];							inform_L[299][1] = l_cell_wire[299];							inform_L[300][1] = l_cell_wire[300];							inform_L[302][1] = l_cell_wire[301];							inform_L[301][1] = l_cell_wire[302];							inform_L[303][1] = l_cell_wire[303];							inform_L[304][1] = l_cell_wire[304];							inform_L[306][1] = l_cell_wire[305];							inform_L[305][1] = l_cell_wire[306];							inform_L[307][1] = l_cell_wire[307];							inform_L[308][1] = l_cell_wire[308];							inform_L[310][1] = l_cell_wire[309];							inform_L[309][1] = l_cell_wire[310];							inform_L[311][1] = l_cell_wire[311];							inform_L[312][1] = l_cell_wire[312];							inform_L[314][1] = l_cell_wire[313];							inform_L[313][1] = l_cell_wire[314];							inform_L[315][1] = l_cell_wire[315];							inform_L[316][1] = l_cell_wire[316];							inform_L[318][1] = l_cell_wire[317];							inform_L[317][1] = l_cell_wire[318];							inform_L[319][1] = l_cell_wire[319];							inform_L[320][1] = l_cell_wire[320];							inform_L[322][1] = l_cell_wire[321];							inform_L[321][1] = l_cell_wire[322];							inform_L[323][1] = l_cell_wire[323];							inform_L[324][1] = l_cell_wire[324];							inform_L[326][1] = l_cell_wire[325];							inform_L[325][1] = l_cell_wire[326];							inform_L[327][1] = l_cell_wire[327];							inform_L[328][1] = l_cell_wire[328];							inform_L[330][1] = l_cell_wire[329];							inform_L[329][1] = l_cell_wire[330];							inform_L[331][1] = l_cell_wire[331];							inform_L[332][1] = l_cell_wire[332];							inform_L[334][1] = l_cell_wire[333];							inform_L[333][1] = l_cell_wire[334];							inform_L[335][1] = l_cell_wire[335];							inform_L[336][1] = l_cell_wire[336];							inform_L[338][1] = l_cell_wire[337];							inform_L[337][1] = l_cell_wire[338];							inform_L[339][1] = l_cell_wire[339];							inform_L[340][1] = l_cell_wire[340];							inform_L[342][1] = l_cell_wire[341];							inform_L[341][1] = l_cell_wire[342];							inform_L[343][1] = l_cell_wire[343];							inform_L[344][1] = l_cell_wire[344];							inform_L[346][1] = l_cell_wire[345];							inform_L[345][1] = l_cell_wire[346];							inform_L[347][1] = l_cell_wire[347];							inform_L[348][1] = l_cell_wire[348];							inform_L[350][1] = l_cell_wire[349];							inform_L[349][1] = l_cell_wire[350];							inform_L[351][1] = l_cell_wire[351];							inform_L[352][1] = l_cell_wire[352];							inform_L[354][1] = l_cell_wire[353];							inform_L[353][1] = l_cell_wire[354];							inform_L[355][1] = l_cell_wire[355];							inform_L[356][1] = l_cell_wire[356];							inform_L[358][1] = l_cell_wire[357];							inform_L[357][1] = l_cell_wire[358];							inform_L[359][1] = l_cell_wire[359];							inform_L[360][1] = l_cell_wire[360];							inform_L[362][1] = l_cell_wire[361];							inform_L[361][1] = l_cell_wire[362];							inform_L[363][1] = l_cell_wire[363];							inform_L[364][1] = l_cell_wire[364];							inform_L[366][1] = l_cell_wire[365];							inform_L[365][1] = l_cell_wire[366];							inform_L[367][1] = l_cell_wire[367];							inform_L[368][1] = l_cell_wire[368];							inform_L[370][1] = l_cell_wire[369];							inform_L[369][1] = l_cell_wire[370];							inform_L[371][1] = l_cell_wire[371];							inform_L[372][1] = l_cell_wire[372];							inform_L[374][1] = l_cell_wire[373];							inform_L[373][1] = l_cell_wire[374];							inform_L[375][1] = l_cell_wire[375];							inform_L[376][1] = l_cell_wire[376];							inform_L[378][1] = l_cell_wire[377];							inform_L[377][1] = l_cell_wire[378];							inform_L[379][1] = l_cell_wire[379];							inform_L[380][1] = l_cell_wire[380];							inform_L[382][1] = l_cell_wire[381];							inform_L[381][1] = l_cell_wire[382];							inform_L[383][1] = l_cell_wire[383];							inform_L[384][1] = l_cell_wire[384];							inform_L[386][1] = l_cell_wire[385];							inform_L[385][1] = l_cell_wire[386];							inform_L[387][1] = l_cell_wire[387];							inform_L[388][1] = l_cell_wire[388];							inform_L[390][1] = l_cell_wire[389];							inform_L[389][1] = l_cell_wire[390];							inform_L[391][1] = l_cell_wire[391];							inform_L[392][1] = l_cell_wire[392];							inform_L[394][1] = l_cell_wire[393];							inform_L[393][1] = l_cell_wire[394];							inform_L[395][1] = l_cell_wire[395];							inform_L[396][1] = l_cell_wire[396];							inform_L[398][1] = l_cell_wire[397];							inform_L[397][1] = l_cell_wire[398];							inform_L[399][1] = l_cell_wire[399];							inform_L[400][1] = l_cell_wire[400];							inform_L[402][1] = l_cell_wire[401];							inform_L[401][1] = l_cell_wire[402];							inform_L[403][1] = l_cell_wire[403];							inform_L[404][1] = l_cell_wire[404];							inform_L[406][1] = l_cell_wire[405];							inform_L[405][1] = l_cell_wire[406];							inform_L[407][1] = l_cell_wire[407];							inform_L[408][1] = l_cell_wire[408];							inform_L[410][1] = l_cell_wire[409];							inform_L[409][1] = l_cell_wire[410];							inform_L[411][1] = l_cell_wire[411];							inform_L[412][1] = l_cell_wire[412];							inform_L[414][1] = l_cell_wire[413];							inform_L[413][1] = l_cell_wire[414];							inform_L[415][1] = l_cell_wire[415];							inform_L[416][1] = l_cell_wire[416];							inform_L[418][1] = l_cell_wire[417];							inform_L[417][1] = l_cell_wire[418];							inform_L[419][1] = l_cell_wire[419];							inform_L[420][1] = l_cell_wire[420];							inform_L[422][1] = l_cell_wire[421];							inform_L[421][1] = l_cell_wire[422];							inform_L[423][1] = l_cell_wire[423];							inform_L[424][1] = l_cell_wire[424];							inform_L[426][1] = l_cell_wire[425];							inform_L[425][1] = l_cell_wire[426];							inform_L[427][1] = l_cell_wire[427];							inform_L[428][1] = l_cell_wire[428];							inform_L[430][1] = l_cell_wire[429];							inform_L[429][1] = l_cell_wire[430];							inform_L[431][1] = l_cell_wire[431];							inform_L[432][1] = l_cell_wire[432];							inform_L[434][1] = l_cell_wire[433];							inform_L[433][1] = l_cell_wire[434];							inform_L[435][1] = l_cell_wire[435];							inform_L[436][1] = l_cell_wire[436];							inform_L[438][1] = l_cell_wire[437];							inform_L[437][1] = l_cell_wire[438];							inform_L[439][1] = l_cell_wire[439];							inform_L[440][1] = l_cell_wire[440];							inform_L[442][1] = l_cell_wire[441];							inform_L[441][1] = l_cell_wire[442];							inform_L[443][1] = l_cell_wire[443];							inform_L[444][1] = l_cell_wire[444];							inform_L[446][1] = l_cell_wire[445];							inform_L[445][1] = l_cell_wire[446];							inform_L[447][1] = l_cell_wire[447];							inform_L[448][1] = l_cell_wire[448];							inform_L[450][1] = l_cell_wire[449];							inform_L[449][1] = l_cell_wire[450];							inform_L[451][1] = l_cell_wire[451];							inform_L[452][1] = l_cell_wire[452];							inform_L[454][1] = l_cell_wire[453];							inform_L[453][1] = l_cell_wire[454];							inform_L[455][1] = l_cell_wire[455];							inform_L[456][1] = l_cell_wire[456];							inform_L[458][1] = l_cell_wire[457];							inform_L[457][1] = l_cell_wire[458];							inform_L[459][1] = l_cell_wire[459];							inform_L[460][1] = l_cell_wire[460];							inform_L[462][1] = l_cell_wire[461];							inform_L[461][1] = l_cell_wire[462];							inform_L[463][1] = l_cell_wire[463];							inform_L[464][1] = l_cell_wire[464];							inform_L[466][1] = l_cell_wire[465];							inform_L[465][1] = l_cell_wire[466];							inform_L[467][1] = l_cell_wire[467];							inform_L[468][1] = l_cell_wire[468];							inform_L[470][1] = l_cell_wire[469];							inform_L[469][1] = l_cell_wire[470];							inform_L[471][1] = l_cell_wire[471];							inform_L[472][1] = l_cell_wire[472];							inform_L[474][1] = l_cell_wire[473];							inform_L[473][1] = l_cell_wire[474];							inform_L[475][1] = l_cell_wire[475];							inform_L[476][1] = l_cell_wire[476];							inform_L[478][1] = l_cell_wire[477];							inform_L[477][1] = l_cell_wire[478];							inform_L[479][1] = l_cell_wire[479];							inform_L[480][1] = l_cell_wire[480];							inform_L[482][1] = l_cell_wire[481];							inform_L[481][1] = l_cell_wire[482];							inform_L[483][1] = l_cell_wire[483];							inform_L[484][1] = l_cell_wire[484];							inform_L[486][1] = l_cell_wire[485];							inform_L[485][1] = l_cell_wire[486];							inform_L[487][1] = l_cell_wire[487];							inform_L[488][1] = l_cell_wire[488];							inform_L[490][1] = l_cell_wire[489];							inform_L[489][1] = l_cell_wire[490];							inform_L[491][1] = l_cell_wire[491];							inform_L[492][1] = l_cell_wire[492];							inform_L[494][1] = l_cell_wire[493];							inform_L[493][1] = l_cell_wire[494];							inform_L[495][1] = l_cell_wire[495];							inform_L[496][1] = l_cell_wire[496];							inform_L[498][1] = l_cell_wire[497];							inform_L[497][1] = l_cell_wire[498];							inform_L[499][1] = l_cell_wire[499];							inform_L[500][1] = l_cell_wire[500];							inform_L[502][1] = l_cell_wire[501];							inform_L[501][1] = l_cell_wire[502];							inform_L[503][1] = l_cell_wire[503];							inform_L[504][1] = l_cell_wire[504];							inform_L[506][1] = l_cell_wire[505];							inform_L[505][1] = l_cell_wire[506];							inform_L[507][1] = l_cell_wire[507];							inform_L[508][1] = l_cell_wire[508];							inform_L[510][1] = l_cell_wire[509];							inform_L[509][1] = l_cell_wire[510];							inform_L[511][1] = l_cell_wire[511];							inform_L[512][1] = l_cell_wire[512];							inform_L[514][1] = l_cell_wire[513];							inform_L[513][1] = l_cell_wire[514];							inform_L[515][1] = l_cell_wire[515];							inform_L[516][1] = l_cell_wire[516];							inform_L[518][1] = l_cell_wire[517];							inform_L[517][1] = l_cell_wire[518];							inform_L[519][1] = l_cell_wire[519];							inform_L[520][1] = l_cell_wire[520];							inform_L[522][1] = l_cell_wire[521];							inform_L[521][1] = l_cell_wire[522];							inform_L[523][1] = l_cell_wire[523];							inform_L[524][1] = l_cell_wire[524];							inform_L[526][1] = l_cell_wire[525];							inform_L[525][1] = l_cell_wire[526];							inform_L[527][1] = l_cell_wire[527];							inform_L[528][1] = l_cell_wire[528];							inform_L[530][1] = l_cell_wire[529];							inform_L[529][1] = l_cell_wire[530];							inform_L[531][1] = l_cell_wire[531];							inform_L[532][1] = l_cell_wire[532];							inform_L[534][1] = l_cell_wire[533];							inform_L[533][1] = l_cell_wire[534];							inform_L[535][1] = l_cell_wire[535];							inform_L[536][1] = l_cell_wire[536];							inform_L[538][1] = l_cell_wire[537];							inform_L[537][1] = l_cell_wire[538];							inform_L[539][1] = l_cell_wire[539];							inform_L[540][1] = l_cell_wire[540];							inform_L[542][1] = l_cell_wire[541];							inform_L[541][1] = l_cell_wire[542];							inform_L[543][1] = l_cell_wire[543];							inform_L[544][1] = l_cell_wire[544];							inform_L[546][1] = l_cell_wire[545];							inform_L[545][1] = l_cell_wire[546];							inform_L[547][1] = l_cell_wire[547];							inform_L[548][1] = l_cell_wire[548];							inform_L[550][1] = l_cell_wire[549];							inform_L[549][1] = l_cell_wire[550];							inform_L[551][1] = l_cell_wire[551];							inform_L[552][1] = l_cell_wire[552];							inform_L[554][1] = l_cell_wire[553];							inform_L[553][1] = l_cell_wire[554];							inform_L[555][1] = l_cell_wire[555];							inform_L[556][1] = l_cell_wire[556];							inform_L[558][1] = l_cell_wire[557];							inform_L[557][1] = l_cell_wire[558];							inform_L[559][1] = l_cell_wire[559];							inform_L[560][1] = l_cell_wire[560];							inform_L[562][1] = l_cell_wire[561];							inform_L[561][1] = l_cell_wire[562];							inform_L[563][1] = l_cell_wire[563];							inform_L[564][1] = l_cell_wire[564];							inform_L[566][1] = l_cell_wire[565];							inform_L[565][1] = l_cell_wire[566];							inform_L[567][1] = l_cell_wire[567];							inform_L[568][1] = l_cell_wire[568];							inform_L[570][1] = l_cell_wire[569];							inform_L[569][1] = l_cell_wire[570];							inform_L[571][1] = l_cell_wire[571];							inform_L[572][1] = l_cell_wire[572];							inform_L[574][1] = l_cell_wire[573];							inform_L[573][1] = l_cell_wire[574];							inform_L[575][1] = l_cell_wire[575];							inform_L[576][1] = l_cell_wire[576];							inform_L[578][1] = l_cell_wire[577];							inform_L[577][1] = l_cell_wire[578];							inform_L[579][1] = l_cell_wire[579];							inform_L[580][1] = l_cell_wire[580];							inform_L[582][1] = l_cell_wire[581];							inform_L[581][1] = l_cell_wire[582];							inform_L[583][1] = l_cell_wire[583];							inform_L[584][1] = l_cell_wire[584];							inform_L[586][1] = l_cell_wire[585];							inform_L[585][1] = l_cell_wire[586];							inform_L[587][1] = l_cell_wire[587];							inform_L[588][1] = l_cell_wire[588];							inform_L[590][1] = l_cell_wire[589];							inform_L[589][1] = l_cell_wire[590];							inform_L[591][1] = l_cell_wire[591];							inform_L[592][1] = l_cell_wire[592];							inform_L[594][1] = l_cell_wire[593];							inform_L[593][1] = l_cell_wire[594];							inform_L[595][1] = l_cell_wire[595];							inform_L[596][1] = l_cell_wire[596];							inform_L[598][1] = l_cell_wire[597];							inform_L[597][1] = l_cell_wire[598];							inform_L[599][1] = l_cell_wire[599];							inform_L[600][1] = l_cell_wire[600];							inform_L[602][1] = l_cell_wire[601];							inform_L[601][1] = l_cell_wire[602];							inform_L[603][1] = l_cell_wire[603];							inform_L[604][1] = l_cell_wire[604];							inform_L[606][1] = l_cell_wire[605];							inform_L[605][1] = l_cell_wire[606];							inform_L[607][1] = l_cell_wire[607];							inform_L[608][1] = l_cell_wire[608];							inform_L[610][1] = l_cell_wire[609];							inform_L[609][1] = l_cell_wire[610];							inform_L[611][1] = l_cell_wire[611];							inform_L[612][1] = l_cell_wire[612];							inform_L[614][1] = l_cell_wire[613];							inform_L[613][1] = l_cell_wire[614];							inform_L[615][1] = l_cell_wire[615];							inform_L[616][1] = l_cell_wire[616];							inform_L[618][1] = l_cell_wire[617];							inform_L[617][1] = l_cell_wire[618];							inform_L[619][1] = l_cell_wire[619];							inform_L[620][1] = l_cell_wire[620];							inform_L[622][1] = l_cell_wire[621];							inform_L[621][1] = l_cell_wire[622];							inform_L[623][1] = l_cell_wire[623];							inform_L[624][1] = l_cell_wire[624];							inform_L[626][1] = l_cell_wire[625];							inform_L[625][1] = l_cell_wire[626];							inform_L[627][1] = l_cell_wire[627];							inform_L[628][1] = l_cell_wire[628];							inform_L[630][1] = l_cell_wire[629];							inform_L[629][1] = l_cell_wire[630];							inform_L[631][1] = l_cell_wire[631];							inform_L[632][1] = l_cell_wire[632];							inform_L[634][1] = l_cell_wire[633];							inform_L[633][1] = l_cell_wire[634];							inform_L[635][1] = l_cell_wire[635];							inform_L[636][1] = l_cell_wire[636];							inform_L[638][1] = l_cell_wire[637];							inform_L[637][1] = l_cell_wire[638];							inform_L[639][1] = l_cell_wire[639];							inform_L[640][1] = l_cell_wire[640];							inform_L[642][1] = l_cell_wire[641];							inform_L[641][1] = l_cell_wire[642];							inform_L[643][1] = l_cell_wire[643];							inform_L[644][1] = l_cell_wire[644];							inform_L[646][1] = l_cell_wire[645];							inform_L[645][1] = l_cell_wire[646];							inform_L[647][1] = l_cell_wire[647];							inform_L[648][1] = l_cell_wire[648];							inform_L[650][1] = l_cell_wire[649];							inform_L[649][1] = l_cell_wire[650];							inform_L[651][1] = l_cell_wire[651];							inform_L[652][1] = l_cell_wire[652];							inform_L[654][1] = l_cell_wire[653];							inform_L[653][1] = l_cell_wire[654];							inform_L[655][1] = l_cell_wire[655];							inform_L[656][1] = l_cell_wire[656];							inform_L[658][1] = l_cell_wire[657];							inform_L[657][1] = l_cell_wire[658];							inform_L[659][1] = l_cell_wire[659];							inform_L[660][1] = l_cell_wire[660];							inform_L[662][1] = l_cell_wire[661];							inform_L[661][1] = l_cell_wire[662];							inform_L[663][1] = l_cell_wire[663];							inform_L[664][1] = l_cell_wire[664];							inform_L[666][1] = l_cell_wire[665];							inform_L[665][1] = l_cell_wire[666];							inform_L[667][1] = l_cell_wire[667];							inform_L[668][1] = l_cell_wire[668];							inform_L[670][1] = l_cell_wire[669];							inform_L[669][1] = l_cell_wire[670];							inform_L[671][1] = l_cell_wire[671];							inform_L[672][1] = l_cell_wire[672];							inform_L[674][1] = l_cell_wire[673];							inform_L[673][1] = l_cell_wire[674];							inform_L[675][1] = l_cell_wire[675];							inform_L[676][1] = l_cell_wire[676];							inform_L[678][1] = l_cell_wire[677];							inform_L[677][1] = l_cell_wire[678];							inform_L[679][1] = l_cell_wire[679];							inform_L[680][1] = l_cell_wire[680];							inform_L[682][1] = l_cell_wire[681];							inform_L[681][1] = l_cell_wire[682];							inform_L[683][1] = l_cell_wire[683];							inform_L[684][1] = l_cell_wire[684];							inform_L[686][1] = l_cell_wire[685];							inform_L[685][1] = l_cell_wire[686];							inform_L[687][1] = l_cell_wire[687];							inform_L[688][1] = l_cell_wire[688];							inform_L[690][1] = l_cell_wire[689];							inform_L[689][1] = l_cell_wire[690];							inform_L[691][1] = l_cell_wire[691];							inform_L[692][1] = l_cell_wire[692];							inform_L[694][1] = l_cell_wire[693];							inform_L[693][1] = l_cell_wire[694];							inform_L[695][1] = l_cell_wire[695];							inform_L[696][1] = l_cell_wire[696];							inform_L[698][1] = l_cell_wire[697];							inform_L[697][1] = l_cell_wire[698];							inform_L[699][1] = l_cell_wire[699];							inform_L[700][1] = l_cell_wire[700];							inform_L[702][1] = l_cell_wire[701];							inform_L[701][1] = l_cell_wire[702];							inform_L[703][1] = l_cell_wire[703];							inform_L[704][1] = l_cell_wire[704];							inform_L[706][1] = l_cell_wire[705];							inform_L[705][1] = l_cell_wire[706];							inform_L[707][1] = l_cell_wire[707];							inform_L[708][1] = l_cell_wire[708];							inform_L[710][1] = l_cell_wire[709];							inform_L[709][1] = l_cell_wire[710];							inform_L[711][1] = l_cell_wire[711];							inform_L[712][1] = l_cell_wire[712];							inform_L[714][1] = l_cell_wire[713];							inform_L[713][1] = l_cell_wire[714];							inform_L[715][1] = l_cell_wire[715];							inform_L[716][1] = l_cell_wire[716];							inform_L[718][1] = l_cell_wire[717];							inform_L[717][1] = l_cell_wire[718];							inform_L[719][1] = l_cell_wire[719];							inform_L[720][1] = l_cell_wire[720];							inform_L[722][1] = l_cell_wire[721];							inform_L[721][1] = l_cell_wire[722];							inform_L[723][1] = l_cell_wire[723];							inform_L[724][1] = l_cell_wire[724];							inform_L[726][1] = l_cell_wire[725];							inform_L[725][1] = l_cell_wire[726];							inform_L[727][1] = l_cell_wire[727];							inform_L[728][1] = l_cell_wire[728];							inform_L[730][1] = l_cell_wire[729];							inform_L[729][1] = l_cell_wire[730];							inform_L[731][1] = l_cell_wire[731];							inform_L[732][1] = l_cell_wire[732];							inform_L[734][1] = l_cell_wire[733];							inform_L[733][1] = l_cell_wire[734];							inform_L[735][1] = l_cell_wire[735];							inform_L[736][1] = l_cell_wire[736];							inform_L[738][1] = l_cell_wire[737];							inform_L[737][1] = l_cell_wire[738];							inform_L[739][1] = l_cell_wire[739];							inform_L[740][1] = l_cell_wire[740];							inform_L[742][1] = l_cell_wire[741];							inform_L[741][1] = l_cell_wire[742];							inform_L[743][1] = l_cell_wire[743];							inform_L[744][1] = l_cell_wire[744];							inform_L[746][1] = l_cell_wire[745];							inform_L[745][1] = l_cell_wire[746];							inform_L[747][1] = l_cell_wire[747];							inform_L[748][1] = l_cell_wire[748];							inform_L[750][1] = l_cell_wire[749];							inform_L[749][1] = l_cell_wire[750];							inform_L[751][1] = l_cell_wire[751];							inform_L[752][1] = l_cell_wire[752];							inform_L[754][1] = l_cell_wire[753];							inform_L[753][1] = l_cell_wire[754];							inform_L[755][1] = l_cell_wire[755];							inform_L[756][1] = l_cell_wire[756];							inform_L[758][1] = l_cell_wire[757];							inform_L[757][1] = l_cell_wire[758];							inform_L[759][1] = l_cell_wire[759];							inform_L[760][1] = l_cell_wire[760];							inform_L[762][1] = l_cell_wire[761];							inform_L[761][1] = l_cell_wire[762];							inform_L[763][1] = l_cell_wire[763];							inform_L[764][1] = l_cell_wire[764];							inform_L[766][1] = l_cell_wire[765];							inform_L[765][1] = l_cell_wire[766];							inform_L[767][1] = l_cell_wire[767];							inform_L[768][1] = l_cell_wire[768];							inform_L[770][1] = l_cell_wire[769];							inform_L[769][1] = l_cell_wire[770];							inform_L[771][1] = l_cell_wire[771];							inform_L[772][1] = l_cell_wire[772];							inform_L[774][1] = l_cell_wire[773];							inform_L[773][1] = l_cell_wire[774];							inform_L[775][1] = l_cell_wire[775];							inform_L[776][1] = l_cell_wire[776];							inform_L[778][1] = l_cell_wire[777];							inform_L[777][1] = l_cell_wire[778];							inform_L[779][1] = l_cell_wire[779];							inform_L[780][1] = l_cell_wire[780];							inform_L[782][1] = l_cell_wire[781];							inform_L[781][1] = l_cell_wire[782];							inform_L[783][1] = l_cell_wire[783];							inform_L[784][1] = l_cell_wire[784];							inform_L[786][1] = l_cell_wire[785];							inform_L[785][1] = l_cell_wire[786];							inform_L[787][1] = l_cell_wire[787];							inform_L[788][1] = l_cell_wire[788];							inform_L[790][1] = l_cell_wire[789];							inform_L[789][1] = l_cell_wire[790];							inform_L[791][1] = l_cell_wire[791];							inform_L[792][1] = l_cell_wire[792];							inform_L[794][1] = l_cell_wire[793];							inform_L[793][1] = l_cell_wire[794];							inform_L[795][1] = l_cell_wire[795];							inform_L[796][1] = l_cell_wire[796];							inform_L[798][1] = l_cell_wire[797];							inform_L[797][1] = l_cell_wire[798];							inform_L[799][1] = l_cell_wire[799];							inform_L[800][1] = l_cell_wire[800];							inform_L[802][1] = l_cell_wire[801];							inform_L[801][1] = l_cell_wire[802];							inform_L[803][1] = l_cell_wire[803];							inform_L[804][1] = l_cell_wire[804];							inform_L[806][1] = l_cell_wire[805];							inform_L[805][1] = l_cell_wire[806];							inform_L[807][1] = l_cell_wire[807];							inform_L[808][1] = l_cell_wire[808];							inform_L[810][1] = l_cell_wire[809];							inform_L[809][1] = l_cell_wire[810];							inform_L[811][1] = l_cell_wire[811];							inform_L[812][1] = l_cell_wire[812];							inform_L[814][1] = l_cell_wire[813];							inform_L[813][1] = l_cell_wire[814];							inform_L[815][1] = l_cell_wire[815];							inform_L[816][1] = l_cell_wire[816];							inform_L[818][1] = l_cell_wire[817];							inform_L[817][1] = l_cell_wire[818];							inform_L[819][1] = l_cell_wire[819];							inform_L[820][1] = l_cell_wire[820];							inform_L[822][1] = l_cell_wire[821];							inform_L[821][1] = l_cell_wire[822];							inform_L[823][1] = l_cell_wire[823];							inform_L[824][1] = l_cell_wire[824];							inform_L[826][1] = l_cell_wire[825];							inform_L[825][1] = l_cell_wire[826];							inform_L[827][1] = l_cell_wire[827];							inform_L[828][1] = l_cell_wire[828];							inform_L[830][1] = l_cell_wire[829];							inform_L[829][1] = l_cell_wire[830];							inform_L[831][1] = l_cell_wire[831];							inform_L[832][1] = l_cell_wire[832];							inform_L[834][1] = l_cell_wire[833];							inform_L[833][1] = l_cell_wire[834];							inform_L[835][1] = l_cell_wire[835];							inform_L[836][1] = l_cell_wire[836];							inform_L[838][1] = l_cell_wire[837];							inform_L[837][1] = l_cell_wire[838];							inform_L[839][1] = l_cell_wire[839];							inform_L[840][1] = l_cell_wire[840];							inform_L[842][1] = l_cell_wire[841];							inform_L[841][1] = l_cell_wire[842];							inform_L[843][1] = l_cell_wire[843];							inform_L[844][1] = l_cell_wire[844];							inform_L[846][1] = l_cell_wire[845];							inform_L[845][1] = l_cell_wire[846];							inform_L[847][1] = l_cell_wire[847];							inform_L[848][1] = l_cell_wire[848];							inform_L[850][1] = l_cell_wire[849];							inform_L[849][1] = l_cell_wire[850];							inform_L[851][1] = l_cell_wire[851];							inform_L[852][1] = l_cell_wire[852];							inform_L[854][1] = l_cell_wire[853];							inform_L[853][1] = l_cell_wire[854];							inform_L[855][1] = l_cell_wire[855];							inform_L[856][1] = l_cell_wire[856];							inform_L[858][1] = l_cell_wire[857];							inform_L[857][1] = l_cell_wire[858];							inform_L[859][1] = l_cell_wire[859];							inform_L[860][1] = l_cell_wire[860];							inform_L[862][1] = l_cell_wire[861];							inform_L[861][1] = l_cell_wire[862];							inform_L[863][1] = l_cell_wire[863];							inform_L[864][1] = l_cell_wire[864];							inform_L[866][1] = l_cell_wire[865];							inform_L[865][1] = l_cell_wire[866];							inform_L[867][1] = l_cell_wire[867];							inform_L[868][1] = l_cell_wire[868];							inform_L[870][1] = l_cell_wire[869];							inform_L[869][1] = l_cell_wire[870];							inform_L[871][1] = l_cell_wire[871];							inform_L[872][1] = l_cell_wire[872];							inform_L[874][1] = l_cell_wire[873];							inform_L[873][1] = l_cell_wire[874];							inform_L[875][1] = l_cell_wire[875];							inform_L[876][1] = l_cell_wire[876];							inform_L[878][1] = l_cell_wire[877];							inform_L[877][1] = l_cell_wire[878];							inform_L[879][1] = l_cell_wire[879];							inform_L[880][1] = l_cell_wire[880];							inform_L[882][1] = l_cell_wire[881];							inform_L[881][1] = l_cell_wire[882];							inform_L[883][1] = l_cell_wire[883];							inform_L[884][1] = l_cell_wire[884];							inform_L[886][1] = l_cell_wire[885];							inform_L[885][1] = l_cell_wire[886];							inform_L[887][1] = l_cell_wire[887];							inform_L[888][1] = l_cell_wire[888];							inform_L[890][1] = l_cell_wire[889];							inform_L[889][1] = l_cell_wire[890];							inform_L[891][1] = l_cell_wire[891];							inform_L[892][1] = l_cell_wire[892];							inform_L[894][1] = l_cell_wire[893];							inform_L[893][1] = l_cell_wire[894];							inform_L[895][1] = l_cell_wire[895];							inform_L[896][1] = l_cell_wire[896];							inform_L[898][1] = l_cell_wire[897];							inform_L[897][1] = l_cell_wire[898];							inform_L[899][1] = l_cell_wire[899];							inform_L[900][1] = l_cell_wire[900];							inform_L[902][1] = l_cell_wire[901];							inform_L[901][1] = l_cell_wire[902];							inform_L[903][1] = l_cell_wire[903];							inform_L[904][1] = l_cell_wire[904];							inform_L[906][1] = l_cell_wire[905];							inform_L[905][1] = l_cell_wire[906];							inform_L[907][1] = l_cell_wire[907];							inform_L[908][1] = l_cell_wire[908];							inform_L[910][1] = l_cell_wire[909];							inform_L[909][1] = l_cell_wire[910];							inform_L[911][1] = l_cell_wire[911];							inform_L[912][1] = l_cell_wire[912];							inform_L[914][1] = l_cell_wire[913];							inform_L[913][1] = l_cell_wire[914];							inform_L[915][1] = l_cell_wire[915];							inform_L[916][1] = l_cell_wire[916];							inform_L[918][1] = l_cell_wire[917];							inform_L[917][1] = l_cell_wire[918];							inform_L[919][1] = l_cell_wire[919];							inform_L[920][1] = l_cell_wire[920];							inform_L[922][1] = l_cell_wire[921];							inform_L[921][1] = l_cell_wire[922];							inform_L[923][1] = l_cell_wire[923];							inform_L[924][1] = l_cell_wire[924];							inform_L[926][1] = l_cell_wire[925];							inform_L[925][1] = l_cell_wire[926];							inform_L[927][1] = l_cell_wire[927];							inform_L[928][1] = l_cell_wire[928];							inform_L[930][1] = l_cell_wire[929];							inform_L[929][1] = l_cell_wire[930];							inform_L[931][1] = l_cell_wire[931];							inform_L[932][1] = l_cell_wire[932];							inform_L[934][1] = l_cell_wire[933];							inform_L[933][1] = l_cell_wire[934];							inform_L[935][1] = l_cell_wire[935];							inform_L[936][1] = l_cell_wire[936];							inform_L[938][1] = l_cell_wire[937];							inform_L[937][1] = l_cell_wire[938];							inform_L[939][1] = l_cell_wire[939];							inform_L[940][1] = l_cell_wire[940];							inform_L[942][1] = l_cell_wire[941];							inform_L[941][1] = l_cell_wire[942];							inform_L[943][1] = l_cell_wire[943];							inform_L[944][1] = l_cell_wire[944];							inform_L[946][1] = l_cell_wire[945];							inform_L[945][1] = l_cell_wire[946];							inform_L[947][1] = l_cell_wire[947];							inform_L[948][1] = l_cell_wire[948];							inform_L[950][1] = l_cell_wire[949];							inform_L[949][1] = l_cell_wire[950];							inform_L[951][1] = l_cell_wire[951];							inform_L[952][1] = l_cell_wire[952];							inform_L[954][1] = l_cell_wire[953];							inform_L[953][1] = l_cell_wire[954];							inform_L[955][1] = l_cell_wire[955];							inform_L[956][1] = l_cell_wire[956];							inform_L[958][1] = l_cell_wire[957];							inform_L[957][1] = l_cell_wire[958];							inform_L[959][1] = l_cell_wire[959];							inform_L[960][1] = l_cell_wire[960];							inform_L[962][1] = l_cell_wire[961];							inform_L[961][1] = l_cell_wire[962];							inform_L[963][1] = l_cell_wire[963];							inform_L[964][1] = l_cell_wire[964];							inform_L[966][1] = l_cell_wire[965];							inform_L[965][1] = l_cell_wire[966];							inform_L[967][1] = l_cell_wire[967];							inform_L[968][1] = l_cell_wire[968];							inform_L[970][1] = l_cell_wire[969];							inform_L[969][1] = l_cell_wire[970];							inform_L[971][1] = l_cell_wire[971];							inform_L[972][1] = l_cell_wire[972];							inform_L[974][1] = l_cell_wire[973];							inform_L[973][1] = l_cell_wire[974];							inform_L[975][1] = l_cell_wire[975];							inform_L[976][1] = l_cell_wire[976];							inform_L[978][1] = l_cell_wire[977];							inform_L[977][1] = l_cell_wire[978];							inform_L[979][1] = l_cell_wire[979];							inform_L[980][1] = l_cell_wire[980];							inform_L[982][1] = l_cell_wire[981];							inform_L[981][1] = l_cell_wire[982];							inform_L[983][1] = l_cell_wire[983];							inform_L[984][1] = l_cell_wire[984];							inform_L[986][1] = l_cell_wire[985];							inform_L[985][1] = l_cell_wire[986];							inform_L[987][1] = l_cell_wire[987];							inform_L[988][1] = l_cell_wire[988];							inform_L[990][1] = l_cell_wire[989];							inform_L[989][1] = l_cell_wire[990];							inform_L[991][1] = l_cell_wire[991];							inform_L[992][1] = l_cell_wire[992];							inform_L[994][1] = l_cell_wire[993];							inform_L[993][1] = l_cell_wire[994];							inform_L[995][1] = l_cell_wire[995];							inform_L[996][1] = l_cell_wire[996];							inform_L[998][1] = l_cell_wire[997];							inform_L[997][1] = l_cell_wire[998];							inform_L[999][1] = l_cell_wire[999];							inform_L[1000][1] = l_cell_wire[1000];							inform_L[1002][1] = l_cell_wire[1001];							inform_L[1001][1] = l_cell_wire[1002];							inform_L[1003][1] = l_cell_wire[1003];							inform_L[1004][1] = l_cell_wire[1004];							inform_L[1006][1] = l_cell_wire[1005];							inform_L[1005][1] = l_cell_wire[1006];							inform_L[1007][1] = l_cell_wire[1007];							inform_L[1008][1] = l_cell_wire[1008];							inform_L[1010][1] = l_cell_wire[1009];							inform_L[1009][1] = l_cell_wire[1010];							inform_L[1011][1] = l_cell_wire[1011];							inform_L[1012][1] = l_cell_wire[1012];							inform_L[1014][1] = l_cell_wire[1013];							inform_L[1013][1] = l_cell_wire[1014];							inform_L[1015][1] = l_cell_wire[1015];							inform_L[1016][1] = l_cell_wire[1016];							inform_L[1018][1] = l_cell_wire[1017];							inform_L[1017][1] = l_cell_wire[1018];							inform_L[1019][1] = l_cell_wire[1019];							inform_L[1020][1] = l_cell_wire[1020];							inform_L[1022][1] = l_cell_wire[1021];							inform_L[1021][1] = l_cell_wire[1022];							inform_L[1023][1] = l_cell_wire[1023];						end
						3:						begin							inform_R[0][3] = r_cell_wire[0];							inform_R[4][3] = r_cell_wire[1];							inform_R[1][3] = r_cell_wire[2];							inform_R[5][3] = r_cell_wire[3];							inform_R[2][3] = r_cell_wire[4];							inform_R[6][3] = r_cell_wire[5];							inform_R[3][3] = r_cell_wire[6];							inform_R[7][3] = r_cell_wire[7];							inform_R[8][3] = r_cell_wire[8];							inform_R[12][3] = r_cell_wire[9];							inform_R[9][3] = r_cell_wire[10];							inform_R[13][3] = r_cell_wire[11];							inform_R[10][3] = r_cell_wire[12];							inform_R[14][3] = r_cell_wire[13];							inform_R[11][3] = r_cell_wire[14];							inform_R[15][3] = r_cell_wire[15];							inform_R[16][3] = r_cell_wire[16];							inform_R[20][3] = r_cell_wire[17];							inform_R[17][3] = r_cell_wire[18];							inform_R[21][3] = r_cell_wire[19];							inform_R[18][3] = r_cell_wire[20];							inform_R[22][3] = r_cell_wire[21];							inform_R[19][3] = r_cell_wire[22];							inform_R[23][3] = r_cell_wire[23];							inform_R[24][3] = r_cell_wire[24];							inform_R[28][3] = r_cell_wire[25];							inform_R[25][3] = r_cell_wire[26];							inform_R[29][3] = r_cell_wire[27];							inform_R[26][3] = r_cell_wire[28];							inform_R[30][3] = r_cell_wire[29];							inform_R[27][3] = r_cell_wire[30];							inform_R[31][3] = r_cell_wire[31];							inform_R[32][3] = r_cell_wire[32];							inform_R[36][3] = r_cell_wire[33];							inform_R[33][3] = r_cell_wire[34];							inform_R[37][3] = r_cell_wire[35];							inform_R[34][3] = r_cell_wire[36];							inform_R[38][3] = r_cell_wire[37];							inform_R[35][3] = r_cell_wire[38];							inform_R[39][3] = r_cell_wire[39];							inform_R[40][3] = r_cell_wire[40];							inform_R[44][3] = r_cell_wire[41];							inform_R[41][3] = r_cell_wire[42];							inform_R[45][3] = r_cell_wire[43];							inform_R[42][3] = r_cell_wire[44];							inform_R[46][3] = r_cell_wire[45];							inform_R[43][3] = r_cell_wire[46];							inform_R[47][3] = r_cell_wire[47];							inform_R[48][3] = r_cell_wire[48];							inform_R[52][3] = r_cell_wire[49];							inform_R[49][3] = r_cell_wire[50];							inform_R[53][3] = r_cell_wire[51];							inform_R[50][3] = r_cell_wire[52];							inform_R[54][3] = r_cell_wire[53];							inform_R[51][3] = r_cell_wire[54];							inform_R[55][3] = r_cell_wire[55];							inform_R[56][3] = r_cell_wire[56];							inform_R[60][3] = r_cell_wire[57];							inform_R[57][3] = r_cell_wire[58];							inform_R[61][3] = r_cell_wire[59];							inform_R[58][3] = r_cell_wire[60];							inform_R[62][3] = r_cell_wire[61];							inform_R[59][3] = r_cell_wire[62];							inform_R[63][3] = r_cell_wire[63];							inform_R[64][3] = r_cell_wire[64];							inform_R[68][3] = r_cell_wire[65];							inform_R[65][3] = r_cell_wire[66];							inform_R[69][3] = r_cell_wire[67];							inform_R[66][3] = r_cell_wire[68];							inform_R[70][3] = r_cell_wire[69];							inform_R[67][3] = r_cell_wire[70];							inform_R[71][3] = r_cell_wire[71];							inform_R[72][3] = r_cell_wire[72];							inform_R[76][3] = r_cell_wire[73];							inform_R[73][3] = r_cell_wire[74];							inform_R[77][3] = r_cell_wire[75];							inform_R[74][3] = r_cell_wire[76];							inform_R[78][3] = r_cell_wire[77];							inform_R[75][3] = r_cell_wire[78];							inform_R[79][3] = r_cell_wire[79];							inform_R[80][3] = r_cell_wire[80];							inform_R[84][3] = r_cell_wire[81];							inform_R[81][3] = r_cell_wire[82];							inform_R[85][3] = r_cell_wire[83];							inform_R[82][3] = r_cell_wire[84];							inform_R[86][3] = r_cell_wire[85];							inform_R[83][3] = r_cell_wire[86];							inform_R[87][3] = r_cell_wire[87];							inform_R[88][3] = r_cell_wire[88];							inform_R[92][3] = r_cell_wire[89];							inform_R[89][3] = r_cell_wire[90];							inform_R[93][3] = r_cell_wire[91];							inform_R[90][3] = r_cell_wire[92];							inform_R[94][3] = r_cell_wire[93];							inform_R[91][3] = r_cell_wire[94];							inform_R[95][3] = r_cell_wire[95];							inform_R[96][3] = r_cell_wire[96];							inform_R[100][3] = r_cell_wire[97];							inform_R[97][3] = r_cell_wire[98];							inform_R[101][3] = r_cell_wire[99];							inform_R[98][3] = r_cell_wire[100];							inform_R[102][3] = r_cell_wire[101];							inform_R[99][3] = r_cell_wire[102];							inform_R[103][3] = r_cell_wire[103];							inform_R[104][3] = r_cell_wire[104];							inform_R[108][3] = r_cell_wire[105];							inform_R[105][3] = r_cell_wire[106];							inform_R[109][3] = r_cell_wire[107];							inform_R[106][3] = r_cell_wire[108];							inform_R[110][3] = r_cell_wire[109];							inform_R[107][3] = r_cell_wire[110];							inform_R[111][3] = r_cell_wire[111];							inform_R[112][3] = r_cell_wire[112];							inform_R[116][3] = r_cell_wire[113];							inform_R[113][3] = r_cell_wire[114];							inform_R[117][3] = r_cell_wire[115];							inform_R[114][3] = r_cell_wire[116];							inform_R[118][3] = r_cell_wire[117];							inform_R[115][3] = r_cell_wire[118];							inform_R[119][3] = r_cell_wire[119];							inform_R[120][3] = r_cell_wire[120];							inform_R[124][3] = r_cell_wire[121];							inform_R[121][3] = r_cell_wire[122];							inform_R[125][3] = r_cell_wire[123];							inform_R[122][3] = r_cell_wire[124];							inform_R[126][3] = r_cell_wire[125];							inform_R[123][3] = r_cell_wire[126];							inform_R[127][3] = r_cell_wire[127];							inform_R[128][3] = r_cell_wire[128];							inform_R[132][3] = r_cell_wire[129];							inform_R[129][3] = r_cell_wire[130];							inform_R[133][3] = r_cell_wire[131];							inform_R[130][3] = r_cell_wire[132];							inform_R[134][3] = r_cell_wire[133];							inform_R[131][3] = r_cell_wire[134];							inform_R[135][3] = r_cell_wire[135];							inform_R[136][3] = r_cell_wire[136];							inform_R[140][3] = r_cell_wire[137];							inform_R[137][3] = r_cell_wire[138];							inform_R[141][3] = r_cell_wire[139];							inform_R[138][3] = r_cell_wire[140];							inform_R[142][3] = r_cell_wire[141];							inform_R[139][3] = r_cell_wire[142];							inform_R[143][3] = r_cell_wire[143];							inform_R[144][3] = r_cell_wire[144];							inform_R[148][3] = r_cell_wire[145];							inform_R[145][3] = r_cell_wire[146];							inform_R[149][3] = r_cell_wire[147];							inform_R[146][3] = r_cell_wire[148];							inform_R[150][3] = r_cell_wire[149];							inform_R[147][3] = r_cell_wire[150];							inform_R[151][3] = r_cell_wire[151];							inform_R[152][3] = r_cell_wire[152];							inform_R[156][3] = r_cell_wire[153];							inform_R[153][3] = r_cell_wire[154];							inform_R[157][3] = r_cell_wire[155];							inform_R[154][3] = r_cell_wire[156];							inform_R[158][3] = r_cell_wire[157];							inform_R[155][3] = r_cell_wire[158];							inform_R[159][3] = r_cell_wire[159];							inform_R[160][3] = r_cell_wire[160];							inform_R[164][3] = r_cell_wire[161];							inform_R[161][3] = r_cell_wire[162];							inform_R[165][3] = r_cell_wire[163];							inform_R[162][3] = r_cell_wire[164];							inform_R[166][3] = r_cell_wire[165];							inform_R[163][3] = r_cell_wire[166];							inform_R[167][3] = r_cell_wire[167];							inform_R[168][3] = r_cell_wire[168];							inform_R[172][3] = r_cell_wire[169];							inform_R[169][3] = r_cell_wire[170];							inform_R[173][3] = r_cell_wire[171];							inform_R[170][3] = r_cell_wire[172];							inform_R[174][3] = r_cell_wire[173];							inform_R[171][3] = r_cell_wire[174];							inform_R[175][3] = r_cell_wire[175];							inform_R[176][3] = r_cell_wire[176];							inform_R[180][3] = r_cell_wire[177];							inform_R[177][3] = r_cell_wire[178];							inform_R[181][3] = r_cell_wire[179];							inform_R[178][3] = r_cell_wire[180];							inform_R[182][3] = r_cell_wire[181];							inform_R[179][3] = r_cell_wire[182];							inform_R[183][3] = r_cell_wire[183];							inform_R[184][3] = r_cell_wire[184];							inform_R[188][3] = r_cell_wire[185];							inform_R[185][3] = r_cell_wire[186];							inform_R[189][3] = r_cell_wire[187];							inform_R[186][3] = r_cell_wire[188];							inform_R[190][3] = r_cell_wire[189];							inform_R[187][3] = r_cell_wire[190];							inform_R[191][3] = r_cell_wire[191];							inform_R[192][3] = r_cell_wire[192];							inform_R[196][3] = r_cell_wire[193];							inform_R[193][3] = r_cell_wire[194];							inform_R[197][3] = r_cell_wire[195];							inform_R[194][3] = r_cell_wire[196];							inform_R[198][3] = r_cell_wire[197];							inform_R[195][3] = r_cell_wire[198];							inform_R[199][3] = r_cell_wire[199];							inform_R[200][3] = r_cell_wire[200];							inform_R[204][3] = r_cell_wire[201];							inform_R[201][3] = r_cell_wire[202];							inform_R[205][3] = r_cell_wire[203];							inform_R[202][3] = r_cell_wire[204];							inform_R[206][3] = r_cell_wire[205];							inform_R[203][3] = r_cell_wire[206];							inform_R[207][3] = r_cell_wire[207];							inform_R[208][3] = r_cell_wire[208];							inform_R[212][3] = r_cell_wire[209];							inform_R[209][3] = r_cell_wire[210];							inform_R[213][3] = r_cell_wire[211];							inform_R[210][3] = r_cell_wire[212];							inform_R[214][3] = r_cell_wire[213];							inform_R[211][3] = r_cell_wire[214];							inform_R[215][3] = r_cell_wire[215];							inform_R[216][3] = r_cell_wire[216];							inform_R[220][3] = r_cell_wire[217];							inform_R[217][3] = r_cell_wire[218];							inform_R[221][3] = r_cell_wire[219];							inform_R[218][3] = r_cell_wire[220];							inform_R[222][3] = r_cell_wire[221];							inform_R[219][3] = r_cell_wire[222];							inform_R[223][3] = r_cell_wire[223];							inform_R[224][3] = r_cell_wire[224];							inform_R[228][3] = r_cell_wire[225];							inform_R[225][3] = r_cell_wire[226];							inform_R[229][3] = r_cell_wire[227];							inform_R[226][3] = r_cell_wire[228];							inform_R[230][3] = r_cell_wire[229];							inform_R[227][3] = r_cell_wire[230];							inform_R[231][3] = r_cell_wire[231];							inform_R[232][3] = r_cell_wire[232];							inform_R[236][3] = r_cell_wire[233];							inform_R[233][3] = r_cell_wire[234];							inform_R[237][3] = r_cell_wire[235];							inform_R[234][3] = r_cell_wire[236];							inform_R[238][3] = r_cell_wire[237];							inform_R[235][3] = r_cell_wire[238];							inform_R[239][3] = r_cell_wire[239];							inform_R[240][3] = r_cell_wire[240];							inform_R[244][3] = r_cell_wire[241];							inform_R[241][3] = r_cell_wire[242];							inform_R[245][3] = r_cell_wire[243];							inform_R[242][3] = r_cell_wire[244];							inform_R[246][3] = r_cell_wire[245];							inform_R[243][3] = r_cell_wire[246];							inform_R[247][3] = r_cell_wire[247];							inform_R[248][3] = r_cell_wire[248];							inform_R[252][3] = r_cell_wire[249];							inform_R[249][3] = r_cell_wire[250];							inform_R[253][3] = r_cell_wire[251];							inform_R[250][3] = r_cell_wire[252];							inform_R[254][3] = r_cell_wire[253];							inform_R[251][3] = r_cell_wire[254];							inform_R[255][3] = r_cell_wire[255];							inform_R[256][3] = r_cell_wire[256];							inform_R[260][3] = r_cell_wire[257];							inform_R[257][3] = r_cell_wire[258];							inform_R[261][3] = r_cell_wire[259];							inform_R[258][3] = r_cell_wire[260];							inform_R[262][3] = r_cell_wire[261];							inform_R[259][3] = r_cell_wire[262];							inform_R[263][3] = r_cell_wire[263];							inform_R[264][3] = r_cell_wire[264];							inform_R[268][3] = r_cell_wire[265];							inform_R[265][3] = r_cell_wire[266];							inform_R[269][3] = r_cell_wire[267];							inform_R[266][3] = r_cell_wire[268];							inform_R[270][3] = r_cell_wire[269];							inform_R[267][3] = r_cell_wire[270];							inform_R[271][3] = r_cell_wire[271];							inform_R[272][3] = r_cell_wire[272];							inform_R[276][3] = r_cell_wire[273];							inform_R[273][3] = r_cell_wire[274];							inform_R[277][3] = r_cell_wire[275];							inform_R[274][3] = r_cell_wire[276];							inform_R[278][3] = r_cell_wire[277];							inform_R[275][3] = r_cell_wire[278];							inform_R[279][3] = r_cell_wire[279];							inform_R[280][3] = r_cell_wire[280];							inform_R[284][3] = r_cell_wire[281];							inform_R[281][3] = r_cell_wire[282];							inform_R[285][3] = r_cell_wire[283];							inform_R[282][3] = r_cell_wire[284];							inform_R[286][3] = r_cell_wire[285];							inform_R[283][3] = r_cell_wire[286];							inform_R[287][3] = r_cell_wire[287];							inform_R[288][3] = r_cell_wire[288];							inform_R[292][3] = r_cell_wire[289];							inform_R[289][3] = r_cell_wire[290];							inform_R[293][3] = r_cell_wire[291];							inform_R[290][3] = r_cell_wire[292];							inform_R[294][3] = r_cell_wire[293];							inform_R[291][3] = r_cell_wire[294];							inform_R[295][3] = r_cell_wire[295];							inform_R[296][3] = r_cell_wire[296];							inform_R[300][3] = r_cell_wire[297];							inform_R[297][3] = r_cell_wire[298];							inform_R[301][3] = r_cell_wire[299];							inform_R[298][3] = r_cell_wire[300];							inform_R[302][3] = r_cell_wire[301];							inform_R[299][3] = r_cell_wire[302];							inform_R[303][3] = r_cell_wire[303];							inform_R[304][3] = r_cell_wire[304];							inform_R[308][3] = r_cell_wire[305];							inform_R[305][3] = r_cell_wire[306];							inform_R[309][3] = r_cell_wire[307];							inform_R[306][3] = r_cell_wire[308];							inform_R[310][3] = r_cell_wire[309];							inform_R[307][3] = r_cell_wire[310];							inform_R[311][3] = r_cell_wire[311];							inform_R[312][3] = r_cell_wire[312];							inform_R[316][3] = r_cell_wire[313];							inform_R[313][3] = r_cell_wire[314];							inform_R[317][3] = r_cell_wire[315];							inform_R[314][3] = r_cell_wire[316];							inform_R[318][3] = r_cell_wire[317];							inform_R[315][3] = r_cell_wire[318];							inform_R[319][3] = r_cell_wire[319];							inform_R[320][3] = r_cell_wire[320];							inform_R[324][3] = r_cell_wire[321];							inform_R[321][3] = r_cell_wire[322];							inform_R[325][3] = r_cell_wire[323];							inform_R[322][3] = r_cell_wire[324];							inform_R[326][3] = r_cell_wire[325];							inform_R[323][3] = r_cell_wire[326];							inform_R[327][3] = r_cell_wire[327];							inform_R[328][3] = r_cell_wire[328];							inform_R[332][3] = r_cell_wire[329];							inform_R[329][3] = r_cell_wire[330];							inform_R[333][3] = r_cell_wire[331];							inform_R[330][3] = r_cell_wire[332];							inform_R[334][3] = r_cell_wire[333];							inform_R[331][3] = r_cell_wire[334];							inform_R[335][3] = r_cell_wire[335];							inform_R[336][3] = r_cell_wire[336];							inform_R[340][3] = r_cell_wire[337];							inform_R[337][3] = r_cell_wire[338];							inform_R[341][3] = r_cell_wire[339];							inform_R[338][3] = r_cell_wire[340];							inform_R[342][3] = r_cell_wire[341];							inform_R[339][3] = r_cell_wire[342];							inform_R[343][3] = r_cell_wire[343];							inform_R[344][3] = r_cell_wire[344];							inform_R[348][3] = r_cell_wire[345];							inform_R[345][3] = r_cell_wire[346];							inform_R[349][3] = r_cell_wire[347];							inform_R[346][3] = r_cell_wire[348];							inform_R[350][3] = r_cell_wire[349];							inform_R[347][3] = r_cell_wire[350];							inform_R[351][3] = r_cell_wire[351];							inform_R[352][3] = r_cell_wire[352];							inform_R[356][3] = r_cell_wire[353];							inform_R[353][3] = r_cell_wire[354];							inform_R[357][3] = r_cell_wire[355];							inform_R[354][3] = r_cell_wire[356];							inform_R[358][3] = r_cell_wire[357];							inform_R[355][3] = r_cell_wire[358];							inform_R[359][3] = r_cell_wire[359];							inform_R[360][3] = r_cell_wire[360];							inform_R[364][3] = r_cell_wire[361];							inform_R[361][3] = r_cell_wire[362];							inform_R[365][3] = r_cell_wire[363];							inform_R[362][3] = r_cell_wire[364];							inform_R[366][3] = r_cell_wire[365];							inform_R[363][3] = r_cell_wire[366];							inform_R[367][3] = r_cell_wire[367];							inform_R[368][3] = r_cell_wire[368];							inform_R[372][3] = r_cell_wire[369];							inform_R[369][3] = r_cell_wire[370];							inform_R[373][3] = r_cell_wire[371];							inform_R[370][3] = r_cell_wire[372];							inform_R[374][3] = r_cell_wire[373];							inform_R[371][3] = r_cell_wire[374];							inform_R[375][3] = r_cell_wire[375];							inform_R[376][3] = r_cell_wire[376];							inform_R[380][3] = r_cell_wire[377];							inform_R[377][3] = r_cell_wire[378];							inform_R[381][3] = r_cell_wire[379];							inform_R[378][3] = r_cell_wire[380];							inform_R[382][3] = r_cell_wire[381];							inform_R[379][3] = r_cell_wire[382];							inform_R[383][3] = r_cell_wire[383];							inform_R[384][3] = r_cell_wire[384];							inform_R[388][3] = r_cell_wire[385];							inform_R[385][3] = r_cell_wire[386];							inform_R[389][3] = r_cell_wire[387];							inform_R[386][3] = r_cell_wire[388];							inform_R[390][3] = r_cell_wire[389];							inform_R[387][3] = r_cell_wire[390];							inform_R[391][3] = r_cell_wire[391];							inform_R[392][3] = r_cell_wire[392];							inform_R[396][3] = r_cell_wire[393];							inform_R[393][3] = r_cell_wire[394];							inform_R[397][3] = r_cell_wire[395];							inform_R[394][3] = r_cell_wire[396];							inform_R[398][3] = r_cell_wire[397];							inform_R[395][3] = r_cell_wire[398];							inform_R[399][3] = r_cell_wire[399];							inform_R[400][3] = r_cell_wire[400];							inform_R[404][3] = r_cell_wire[401];							inform_R[401][3] = r_cell_wire[402];							inform_R[405][3] = r_cell_wire[403];							inform_R[402][3] = r_cell_wire[404];							inform_R[406][3] = r_cell_wire[405];							inform_R[403][3] = r_cell_wire[406];							inform_R[407][3] = r_cell_wire[407];							inform_R[408][3] = r_cell_wire[408];							inform_R[412][3] = r_cell_wire[409];							inform_R[409][3] = r_cell_wire[410];							inform_R[413][3] = r_cell_wire[411];							inform_R[410][3] = r_cell_wire[412];							inform_R[414][3] = r_cell_wire[413];							inform_R[411][3] = r_cell_wire[414];							inform_R[415][3] = r_cell_wire[415];							inform_R[416][3] = r_cell_wire[416];							inform_R[420][3] = r_cell_wire[417];							inform_R[417][3] = r_cell_wire[418];							inform_R[421][3] = r_cell_wire[419];							inform_R[418][3] = r_cell_wire[420];							inform_R[422][3] = r_cell_wire[421];							inform_R[419][3] = r_cell_wire[422];							inform_R[423][3] = r_cell_wire[423];							inform_R[424][3] = r_cell_wire[424];							inform_R[428][3] = r_cell_wire[425];							inform_R[425][3] = r_cell_wire[426];							inform_R[429][3] = r_cell_wire[427];							inform_R[426][3] = r_cell_wire[428];							inform_R[430][3] = r_cell_wire[429];							inform_R[427][3] = r_cell_wire[430];							inform_R[431][3] = r_cell_wire[431];							inform_R[432][3] = r_cell_wire[432];							inform_R[436][3] = r_cell_wire[433];							inform_R[433][3] = r_cell_wire[434];							inform_R[437][3] = r_cell_wire[435];							inform_R[434][3] = r_cell_wire[436];							inform_R[438][3] = r_cell_wire[437];							inform_R[435][3] = r_cell_wire[438];							inform_R[439][3] = r_cell_wire[439];							inform_R[440][3] = r_cell_wire[440];							inform_R[444][3] = r_cell_wire[441];							inform_R[441][3] = r_cell_wire[442];							inform_R[445][3] = r_cell_wire[443];							inform_R[442][3] = r_cell_wire[444];							inform_R[446][3] = r_cell_wire[445];							inform_R[443][3] = r_cell_wire[446];							inform_R[447][3] = r_cell_wire[447];							inform_R[448][3] = r_cell_wire[448];							inform_R[452][3] = r_cell_wire[449];							inform_R[449][3] = r_cell_wire[450];							inform_R[453][3] = r_cell_wire[451];							inform_R[450][3] = r_cell_wire[452];							inform_R[454][3] = r_cell_wire[453];							inform_R[451][3] = r_cell_wire[454];							inform_R[455][3] = r_cell_wire[455];							inform_R[456][3] = r_cell_wire[456];							inform_R[460][3] = r_cell_wire[457];							inform_R[457][3] = r_cell_wire[458];							inform_R[461][3] = r_cell_wire[459];							inform_R[458][3] = r_cell_wire[460];							inform_R[462][3] = r_cell_wire[461];							inform_R[459][3] = r_cell_wire[462];							inform_R[463][3] = r_cell_wire[463];							inform_R[464][3] = r_cell_wire[464];							inform_R[468][3] = r_cell_wire[465];							inform_R[465][3] = r_cell_wire[466];							inform_R[469][3] = r_cell_wire[467];							inform_R[466][3] = r_cell_wire[468];							inform_R[470][3] = r_cell_wire[469];							inform_R[467][3] = r_cell_wire[470];							inform_R[471][3] = r_cell_wire[471];							inform_R[472][3] = r_cell_wire[472];							inform_R[476][3] = r_cell_wire[473];							inform_R[473][3] = r_cell_wire[474];							inform_R[477][3] = r_cell_wire[475];							inform_R[474][3] = r_cell_wire[476];							inform_R[478][3] = r_cell_wire[477];							inform_R[475][3] = r_cell_wire[478];							inform_R[479][3] = r_cell_wire[479];							inform_R[480][3] = r_cell_wire[480];							inform_R[484][3] = r_cell_wire[481];							inform_R[481][3] = r_cell_wire[482];							inform_R[485][3] = r_cell_wire[483];							inform_R[482][3] = r_cell_wire[484];							inform_R[486][3] = r_cell_wire[485];							inform_R[483][3] = r_cell_wire[486];							inform_R[487][3] = r_cell_wire[487];							inform_R[488][3] = r_cell_wire[488];							inform_R[492][3] = r_cell_wire[489];							inform_R[489][3] = r_cell_wire[490];							inform_R[493][3] = r_cell_wire[491];							inform_R[490][3] = r_cell_wire[492];							inform_R[494][3] = r_cell_wire[493];							inform_R[491][3] = r_cell_wire[494];							inform_R[495][3] = r_cell_wire[495];							inform_R[496][3] = r_cell_wire[496];							inform_R[500][3] = r_cell_wire[497];							inform_R[497][3] = r_cell_wire[498];							inform_R[501][3] = r_cell_wire[499];							inform_R[498][3] = r_cell_wire[500];							inform_R[502][3] = r_cell_wire[501];							inform_R[499][3] = r_cell_wire[502];							inform_R[503][3] = r_cell_wire[503];							inform_R[504][3] = r_cell_wire[504];							inform_R[508][3] = r_cell_wire[505];							inform_R[505][3] = r_cell_wire[506];							inform_R[509][3] = r_cell_wire[507];							inform_R[506][3] = r_cell_wire[508];							inform_R[510][3] = r_cell_wire[509];							inform_R[507][3] = r_cell_wire[510];							inform_R[511][3] = r_cell_wire[511];							inform_R[512][3] = r_cell_wire[512];							inform_R[516][3] = r_cell_wire[513];							inform_R[513][3] = r_cell_wire[514];							inform_R[517][3] = r_cell_wire[515];							inform_R[514][3] = r_cell_wire[516];							inform_R[518][3] = r_cell_wire[517];							inform_R[515][3] = r_cell_wire[518];							inform_R[519][3] = r_cell_wire[519];							inform_R[520][3] = r_cell_wire[520];							inform_R[524][3] = r_cell_wire[521];							inform_R[521][3] = r_cell_wire[522];							inform_R[525][3] = r_cell_wire[523];							inform_R[522][3] = r_cell_wire[524];							inform_R[526][3] = r_cell_wire[525];							inform_R[523][3] = r_cell_wire[526];							inform_R[527][3] = r_cell_wire[527];							inform_R[528][3] = r_cell_wire[528];							inform_R[532][3] = r_cell_wire[529];							inform_R[529][3] = r_cell_wire[530];							inform_R[533][3] = r_cell_wire[531];							inform_R[530][3] = r_cell_wire[532];							inform_R[534][3] = r_cell_wire[533];							inform_R[531][3] = r_cell_wire[534];							inform_R[535][3] = r_cell_wire[535];							inform_R[536][3] = r_cell_wire[536];							inform_R[540][3] = r_cell_wire[537];							inform_R[537][3] = r_cell_wire[538];							inform_R[541][3] = r_cell_wire[539];							inform_R[538][3] = r_cell_wire[540];							inform_R[542][3] = r_cell_wire[541];							inform_R[539][3] = r_cell_wire[542];							inform_R[543][3] = r_cell_wire[543];							inform_R[544][3] = r_cell_wire[544];							inform_R[548][3] = r_cell_wire[545];							inform_R[545][3] = r_cell_wire[546];							inform_R[549][3] = r_cell_wire[547];							inform_R[546][3] = r_cell_wire[548];							inform_R[550][3] = r_cell_wire[549];							inform_R[547][3] = r_cell_wire[550];							inform_R[551][3] = r_cell_wire[551];							inform_R[552][3] = r_cell_wire[552];							inform_R[556][3] = r_cell_wire[553];							inform_R[553][3] = r_cell_wire[554];							inform_R[557][3] = r_cell_wire[555];							inform_R[554][3] = r_cell_wire[556];							inform_R[558][3] = r_cell_wire[557];							inform_R[555][3] = r_cell_wire[558];							inform_R[559][3] = r_cell_wire[559];							inform_R[560][3] = r_cell_wire[560];							inform_R[564][3] = r_cell_wire[561];							inform_R[561][3] = r_cell_wire[562];							inform_R[565][3] = r_cell_wire[563];							inform_R[562][3] = r_cell_wire[564];							inform_R[566][3] = r_cell_wire[565];							inform_R[563][3] = r_cell_wire[566];							inform_R[567][3] = r_cell_wire[567];							inform_R[568][3] = r_cell_wire[568];							inform_R[572][3] = r_cell_wire[569];							inform_R[569][3] = r_cell_wire[570];							inform_R[573][3] = r_cell_wire[571];							inform_R[570][3] = r_cell_wire[572];							inform_R[574][3] = r_cell_wire[573];							inform_R[571][3] = r_cell_wire[574];							inform_R[575][3] = r_cell_wire[575];							inform_R[576][3] = r_cell_wire[576];							inform_R[580][3] = r_cell_wire[577];							inform_R[577][3] = r_cell_wire[578];							inform_R[581][3] = r_cell_wire[579];							inform_R[578][3] = r_cell_wire[580];							inform_R[582][3] = r_cell_wire[581];							inform_R[579][3] = r_cell_wire[582];							inform_R[583][3] = r_cell_wire[583];							inform_R[584][3] = r_cell_wire[584];							inform_R[588][3] = r_cell_wire[585];							inform_R[585][3] = r_cell_wire[586];							inform_R[589][3] = r_cell_wire[587];							inform_R[586][3] = r_cell_wire[588];							inform_R[590][3] = r_cell_wire[589];							inform_R[587][3] = r_cell_wire[590];							inform_R[591][3] = r_cell_wire[591];							inform_R[592][3] = r_cell_wire[592];							inform_R[596][3] = r_cell_wire[593];							inform_R[593][3] = r_cell_wire[594];							inform_R[597][3] = r_cell_wire[595];							inform_R[594][3] = r_cell_wire[596];							inform_R[598][3] = r_cell_wire[597];							inform_R[595][3] = r_cell_wire[598];							inform_R[599][3] = r_cell_wire[599];							inform_R[600][3] = r_cell_wire[600];							inform_R[604][3] = r_cell_wire[601];							inform_R[601][3] = r_cell_wire[602];							inform_R[605][3] = r_cell_wire[603];							inform_R[602][3] = r_cell_wire[604];							inform_R[606][3] = r_cell_wire[605];							inform_R[603][3] = r_cell_wire[606];							inform_R[607][3] = r_cell_wire[607];							inform_R[608][3] = r_cell_wire[608];							inform_R[612][3] = r_cell_wire[609];							inform_R[609][3] = r_cell_wire[610];							inform_R[613][3] = r_cell_wire[611];							inform_R[610][3] = r_cell_wire[612];							inform_R[614][3] = r_cell_wire[613];							inform_R[611][3] = r_cell_wire[614];							inform_R[615][3] = r_cell_wire[615];							inform_R[616][3] = r_cell_wire[616];							inform_R[620][3] = r_cell_wire[617];							inform_R[617][3] = r_cell_wire[618];							inform_R[621][3] = r_cell_wire[619];							inform_R[618][3] = r_cell_wire[620];							inform_R[622][3] = r_cell_wire[621];							inform_R[619][3] = r_cell_wire[622];							inform_R[623][3] = r_cell_wire[623];							inform_R[624][3] = r_cell_wire[624];							inform_R[628][3] = r_cell_wire[625];							inform_R[625][3] = r_cell_wire[626];							inform_R[629][3] = r_cell_wire[627];							inform_R[626][3] = r_cell_wire[628];							inform_R[630][3] = r_cell_wire[629];							inform_R[627][3] = r_cell_wire[630];							inform_R[631][3] = r_cell_wire[631];							inform_R[632][3] = r_cell_wire[632];							inform_R[636][3] = r_cell_wire[633];							inform_R[633][3] = r_cell_wire[634];							inform_R[637][3] = r_cell_wire[635];							inform_R[634][3] = r_cell_wire[636];							inform_R[638][3] = r_cell_wire[637];							inform_R[635][3] = r_cell_wire[638];							inform_R[639][3] = r_cell_wire[639];							inform_R[640][3] = r_cell_wire[640];							inform_R[644][3] = r_cell_wire[641];							inform_R[641][3] = r_cell_wire[642];							inform_R[645][3] = r_cell_wire[643];							inform_R[642][3] = r_cell_wire[644];							inform_R[646][3] = r_cell_wire[645];							inform_R[643][3] = r_cell_wire[646];							inform_R[647][3] = r_cell_wire[647];							inform_R[648][3] = r_cell_wire[648];							inform_R[652][3] = r_cell_wire[649];							inform_R[649][3] = r_cell_wire[650];							inform_R[653][3] = r_cell_wire[651];							inform_R[650][3] = r_cell_wire[652];							inform_R[654][3] = r_cell_wire[653];							inform_R[651][3] = r_cell_wire[654];							inform_R[655][3] = r_cell_wire[655];							inform_R[656][3] = r_cell_wire[656];							inform_R[660][3] = r_cell_wire[657];							inform_R[657][3] = r_cell_wire[658];							inform_R[661][3] = r_cell_wire[659];							inform_R[658][3] = r_cell_wire[660];							inform_R[662][3] = r_cell_wire[661];							inform_R[659][3] = r_cell_wire[662];							inform_R[663][3] = r_cell_wire[663];							inform_R[664][3] = r_cell_wire[664];							inform_R[668][3] = r_cell_wire[665];							inform_R[665][3] = r_cell_wire[666];							inform_R[669][3] = r_cell_wire[667];							inform_R[666][3] = r_cell_wire[668];							inform_R[670][3] = r_cell_wire[669];							inform_R[667][3] = r_cell_wire[670];							inform_R[671][3] = r_cell_wire[671];							inform_R[672][3] = r_cell_wire[672];							inform_R[676][3] = r_cell_wire[673];							inform_R[673][3] = r_cell_wire[674];							inform_R[677][3] = r_cell_wire[675];							inform_R[674][3] = r_cell_wire[676];							inform_R[678][3] = r_cell_wire[677];							inform_R[675][3] = r_cell_wire[678];							inform_R[679][3] = r_cell_wire[679];							inform_R[680][3] = r_cell_wire[680];							inform_R[684][3] = r_cell_wire[681];							inform_R[681][3] = r_cell_wire[682];							inform_R[685][3] = r_cell_wire[683];							inform_R[682][3] = r_cell_wire[684];							inform_R[686][3] = r_cell_wire[685];							inform_R[683][3] = r_cell_wire[686];							inform_R[687][3] = r_cell_wire[687];							inform_R[688][3] = r_cell_wire[688];							inform_R[692][3] = r_cell_wire[689];							inform_R[689][3] = r_cell_wire[690];							inform_R[693][3] = r_cell_wire[691];							inform_R[690][3] = r_cell_wire[692];							inform_R[694][3] = r_cell_wire[693];							inform_R[691][3] = r_cell_wire[694];							inform_R[695][3] = r_cell_wire[695];							inform_R[696][3] = r_cell_wire[696];							inform_R[700][3] = r_cell_wire[697];							inform_R[697][3] = r_cell_wire[698];							inform_R[701][3] = r_cell_wire[699];							inform_R[698][3] = r_cell_wire[700];							inform_R[702][3] = r_cell_wire[701];							inform_R[699][3] = r_cell_wire[702];							inform_R[703][3] = r_cell_wire[703];							inform_R[704][3] = r_cell_wire[704];							inform_R[708][3] = r_cell_wire[705];							inform_R[705][3] = r_cell_wire[706];							inform_R[709][3] = r_cell_wire[707];							inform_R[706][3] = r_cell_wire[708];							inform_R[710][3] = r_cell_wire[709];							inform_R[707][3] = r_cell_wire[710];							inform_R[711][3] = r_cell_wire[711];							inform_R[712][3] = r_cell_wire[712];							inform_R[716][3] = r_cell_wire[713];							inform_R[713][3] = r_cell_wire[714];							inform_R[717][3] = r_cell_wire[715];							inform_R[714][3] = r_cell_wire[716];							inform_R[718][3] = r_cell_wire[717];							inform_R[715][3] = r_cell_wire[718];							inform_R[719][3] = r_cell_wire[719];							inform_R[720][3] = r_cell_wire[720];							inform_R[724][3] = r_cell_wire[721];							inform_R[721][3] = r_cell_wire[722];							inform_R[725][3] = r_cell_wire[723];							inform_R[722][3] = r_cell_wire[724];							inform_R[726][3] = r_cell_wire[725];							inform_R[723][3] = r_cell_wire[726];							inform_R[727][3] = r_cell_wire[727];							inform_R[728][3] = r_cell_wire[728];							inform_R[732][3] = r_cell_wire[729];							inform_R[729][3] = r_cell_wire[730];							inform_R[733][3] = r_cell_wire[731];							inform_R[730][3] = r_cell_wire[732];							inform_R[734][3] = r_cell_wire[733];							inform_R[731][3] = r_cell_wire[734];							inform_R[735][3] = r_cell_wire[735];							inform_R[736][3] = r_cell_wire[736];							inform_R[740][3] = r_cell_wire[737];							inform_R[737][3] = r_cell_wire[738];							inform_R[741][3] = r_cell_wire[739];							inform_R[738][3] = r_cell_wire[740];							inform_R[742][3] = r_cell_wire[741];							inform_R[739][3] = r_cell_wire[742];							inform_R[743][3] = r_cell_wire[743];							inform_R[744][3] = r_cell_wire[744];							inform_R[748][3] = r_cell_wire[745];							inform_R[745][3] = r_cell_wire[746];							inform_R[749][3] = r_cell_wire[747];							inform_R[746][3] = r_cell_wire[748];							inform_R[750][3] = r_cell_wire[749];							inform_R[747][3] = r_cell_wire[750];							inform_R[751][3] = r_cell_wire[751];							inform_R[752][3] = r_cell_wire[752];							inform_R[756][3] = r_cell_wire[753];							inform_R[753][3] = r_cell_wire[754];							inform_R[757][3] = r_cell_wire[755];							inform_R[754][3] = r_cell_wire[756];							inform_R[758][3] = r_cell_wire[757];							inform_R[755][3] = r_cell_wire[758];							inform_R[759][3] = r_cell_wire[759];							inform_R[760][3] = r_cell_wire[760];							inform_R[764][3] = r_cell_wire[761];							inform_R[761][3] = r_cell_wire[762];							inform_R[765][3] = r_cell_wire[763];							inform_R[762][3] = r_cell_wire[764];							inform_R[766][3] = r_cell_wire[765];							inform_R[763][3] = r_cell_wire[766];							inform_R[767][3] = r_cell_wire[767];							inform_R[768][3] = r_cell_wire[768];							inform_R[772][3] = r_cell_wire[769];							inform_R[769][3] = r_cell_wire[770];							inform_R[773][3] = r_cell_wire[771];							inform_R[770][3] = r_cell_wire[772];							inform_R[774][3] = r_cell_wire[773];							inform_R[771][3] = r_cell_wire[774];							inform_R[775][3] = r_cell_wire[775];							inform_R[776][3] = r_cell_wire[776];							inform_R[780][3] = r_cell_wire[777];							inform_R[777][3] = r_cell_wire[778];							inform_R[781][3] = r_cell_wire[779];							inform_R[778][3] = r_cell_wire[780];							inform_R[782][3] = r_cell_wire[781];							inform_R[779][3] = r_cell_wire[782];							inform_R[783][3] = r_cell_wire[783];							inform_R[784][3] = r_cell_wire[784];							inform_R[788][3] = r_cell_wire[785];							inform_R[785][3] = r_cell_wire[786];							inform_R[789][3] = r_cell_wire[787];							inform_R[786][3] = r_cell_wire[788];							inform_R[790][3] = r_cell_wire[789];							inform_R[787][3] = r_cell_wire[790];							inform_R[791][3] = r_cell_wire[791];							inform_R[792][3] = r_cell_wire[792];							inform_R[796][3] = r_cell_wire[793];							inform_R[793][3] = r_cell_wire[794];							inform_R[797][3] = r_cell_wire[795];							inform_R[794][3] = r_cell_wire[796];							inform_R[798][3] = r_cell_wire[797];							inform_R[795][3] = r_cell_wire[798];							inform_R[799][3] = r_cell_wire[799];							inform_R[800][3] = r_cell_wire[800];							inform_R[804][3] = r_cell_wire[801];							inform_R[801][3] = r_cell_wire[802];							inform_R[805][3] = r_cell_wire[803];							inform_R[802][3] = r_cell_wire[804];							inform_R[806][3] = r_cell_wire[805];							inform_R[803][3] = r_cell_wire[806];							inform_R[807][3] = r_cell_wire[807];							inform_R[808][3] = r_cell_wire[808];							inform_R[812][3] = r_cell_wire[809];							inform_R[809][3] = r_cell_wire[810];							inform_R[813][3] = r_cell_wire[811];							inform_R[810][3] = r_cell_wire[812];							inform_R[814][3] = r_cell_wire[813];							inform_R[811][3] = r_cell_wire[814];							inform_R[815][3] = r_cell_wire[815];							inform_R[816][3] = r_cell_wire[816];							inform_R[820][3] = r_cell_wire[817];							inform_R[817][3] = r_cell_wire[818];							inform_R[821][3] = r_cell_wire[819];							inform_R[818][3] = r_cell_wire[820];							inform_R[822][3] = r_cell_wire[821];							inform_R[819][3] = r_cell_wire[822];							inform_R[823][3] = r_cell_wire[823];							inform_R[824][3] = r_cell_wire[824];							inform_R[828][3] = r_cell_wire[825];							inform_R[825][3] = r_cell_wire[826];							inform_R[829][3] = r_cell_wire[827];							inform_R[826][3] = r_cell_wire[828];							inform_R[830][3] = r_cell_wire[829];							inform_R[827][3] = r_cell_wire[830];							inform_R[831][3] = r_cell_wire[831];							inform_R[832][3] = r_cell_wire[832];							inform_R[836][3] = r_cell_wire[833];							inform_R[833][3] = r_cell_wire[834];							inform_R[837][3] = r_cell_wire[835];							inform_R[834][3] = r_cell_wire[836];							inform_R[838][3] = r_cell_wire[837];							inform_R[835][3] = r_cell_wire[838];							inform_R[839][3] = r_cell_wire[839];							inform_R[840][3] = r_cell_wire[840];							inform_R[844][3] = r_cell_wire[841];							inform_R[841][3] = r_cell_wire[842];							inform_R[845][3] = r_cell_wire[843];							inform_R[842][3] = r_cell_wire[844];							inform_R[846][3] = r_cell_wire[845];							inform_R[843][3] = r_cell_wire[846];							inform_R[847][3] = r_cell_wire[847];							inform_R[848][3] = r_cell_wire[848];							inform_R[852][3] = r_cell_wire[849];							inform_R[849][3] = r_cell_wire[850];							inform_R[853][3] = r_cell_wire[851];							inform_R[850][3] = r_cell_wire[852];							inform_R[854][3] = r_cell_wire[853];							inform_R[851][3] = r_cell_wire[854];							inform_R[855][3] = r_cell_wire[855];							inform_R[856][3] = r_cell_wire[856];							inform_R[860][3] = r_cell_wire[857];							inform_R[857][3] = r_cell_wire[858];							inform_R[861][3] = r_cell_wire[859];							inform_R[858][3] = r_cell_wire[860];							inform_R[862][3] = r_cell_wire[861];							inform_R[859][3] = r_cell_wire[862];							inform_R[863][3] = r_cell_wire[863];							inform_R[864][3] = r_cell_wire[864];							inform_R[868][3] = r_cell_wire[865];							inform_R[865][3] = r_cell_wire[866];							inform_R[869][3] = r_cell_wire[867];							inform_R[866][3] = r_cell_wire[868];							inform_R[870][3] = r_cell_wire[869];							inform_R[867][3] = r_cell_wire[870];							inform_R[871][3] = r_cell_wire[871];							inform_R[872][3] = r_cell_wire[872];							inform_R[876][3] = r_cell_wire[873];							inform_R[873][3] = r_cell_wire[874];							inform_R[877][3] = r_cell_wire[875];							inform_R[874][3] = r_cell_wire[876];							inform_R[878][3] = r_cell_wire[877];							inform_R[875][3] = r_cell_wire[878];							inform_R[879][3] = r_cell_wire[879];							inform_R[880][3] = r_cell_wire[880];							inform_R[884][3] = r_cell_wire[881];							inform_R[881][3] = r_cell_wire[882];							inform_R[885][3] = r_cell_wire[883];							inform_R[882][3] = r_cell_wire[884];							inform_R[886][3] = r_cell_wire[885];							inform_R[883][3] = r_cell_wire[886];							inform_R[887][3] = r_cell_wire[887];							inform_R[888][3] = r_cell_wire[888];							inform_R[892][3] = r_cell_wire[889];							inform_R[889][3] = r_cell_wire[890];							inform_R[893][3] = r_cell_wire[891];							inform_R[890][3] = r_cell_wire[892];							inform_R[894][3] = r_cell_wire[893];							inform_R[891][3] = r_cell_wire[894];							inform_R[895][3] = r_cell_wire[895];							inform_R[896][3] = r_cell_wire[896];							inform_R[900][3] = r_cell_wire[897];							inform_R[897][3] = r_cell_wire[898];							inform_R[901][3] = r_cell_wire[899];							inform_R[898][3] = r_cell_wire[900];							inform_R[902][3] = r_cell_wire[901];							inform_R[899][3] = r_cell_wire[902];							inform_R[903][3] = r_cell_wire[903];							inform_R[904][3] = r_cell_wire[904];							inform_R[908][3] = r_cell_wire[905];							inform_R[905][3] = r_cell_wire[906];							inform_R[909][3] = r_cell_wire[907];							inform_R[906][3] = r_cell_wire[908];							inform_R[910][3] = r_cell_wire[909];							inform_R[907][3] = r_cell_wire[910];							inform_R[911][3] = r_cell_wire[911];							inform_R[912][3] = r_cell_wire[912];							inform_R[916][3] = r_cell_wire[913];							inform_R[913][3] = r_cell_wire[914];							inform_R[917][3] = r_cell_wire[915];							inform_R[914][3] = r_cell_wire[916];							inform_R[918][3] = r_cell_wire[917];							inform_R[915][3] = r_cell_wire[918];							inform_R[919][3] = r_cell_wire[919];							inform_R[920][3] = r_cell_wire[920];							inform_R[924][3] = r_cell_wire[921];							inform_R[921][3] = r_cell_wire[922];							inform_R[925][3] = r_cell_wire[923];							inform_R[922][3] = r_cell_wire[924];							inform_R[926][3] = r_cell_wire[925];							inform_R[923][3] = r_cell_wire[926];							inform_R[927][3] = r_cell_wire[927];							inform_R[928][3] = r_cell_wire[928];							inform_R[932][3] = r_cell_wire[929];							inform_R[929][3] = r_cell_wire[930];							inform_R[933][3] = r_cell_wire[931];							inform_R[930][3] = r_cell_wire[932];							inform_R[934][3] = r_cell_wire[933];							inform_R[931][3] = r_cell_wire[934];							inform_R[935][3] = r_cell_wire[935];							inform_R[936][3] = r_cell_wire[936];							inform_R[940][3] = r_cell_wire[937];							inform_R[937][3] = r_cell_wire[938];							inform_R[941][3] = r_cell_wire[939];							inform_R[938][3] = r_cell_wire[940];							inform_R[942][3] = r_cell_wire[941];							inform_R[939][3] = r_cell_wire[942];							inform_R[943][3] = r_cell_wire[943];							inform_R[944][3] = r_cell_wire[944];							inform_R[948][3] = r_cell_wire[945];							inform_R[945][3] = r_cell_wire[946];							inform_R[949][3] = r_cell_wire[947];							inform_R[946][3] = r_cell_wire[948];							inform_R[950][3] = r_cell_wire[949];							inform_R[947][3] = r_cell_wire[950];							inform_R[951][3] = r_cell_wire[951];							inform_R[952][3] = r_cell_wire[952];							inform_R[956][3] = r_cell_wire[953];							inform_R[953][3] = r_cell_wire[954];							inform_R[957][3] = r_cell_wire[955];							inform_R[954][3] = r_cell_wire[956];							inform_R[958][3] = r_cell_wire[957];							inform_R[955][3] = r_cell_wire[958];							inform_R[959][3] = r_cell_wire[959];							inform_R[960][3] = r_cell_wire[960];							inform_R[964][3] = r_cell_wire[961];							inform_R[961][3] = r_cell_wire[962];							inform_R[965][3] = r_cell_wire[963];							inform_R[962][3] = r_cell_wire[964];							inform_R[966][3] = r_cell_wire[965];							inform_R[963][3] = r_cell_wire[966];							inform_R[967][3] = r_cell_wire[967];							inform_R[968][3] = r_cell_wire[968];							inform_R[972][3] = r_cell_wire[969];							inform_R[969][3] = r_cell_wire[970];							inform_R[973][3] = r_cell_wire[971];							inform_R[970][3] = r_cell_wire[972];							inform_R[974][3] = r_cell_wire[973];							inform_R[971][3] = r_cell_wire[974];							inform_R[975][3] = r_cell_wire[975];							inform_R[976][3] = r_cell_wire[976];							inform_R[980][3] = r_cell_wire[977];							inform_R[977][3] = r_cell_wire[978];							inform_R[981][3] = r_cell_wire[979];							inform_R[978][3] = r_cell_wire[980];							inform_R[982][3] = r_cell_wire[981];							inform_R[979][3] = r_cell_wire[982];							inform_R[983][3] = r_cell_wire[983];							inform_R[984][3] = r_cell_wire[984];							inform_R[988][3] = r_cell_wire[985];							inform_R[985][3] = r_cell_wire[986];							inform_R[989][3] = r_cell_wire[987];							inform_R[986][3] = r_cell_wire[988];							inform_R[990][3] = r_cell_wire[989];							inform_R[987][3] = r_cell_wire[990];							inform_R[991][3] = r_cell_wire[991];							inform_R[992][3] = r_cell_wire[992];							inform_R[996][3] = r_cell_wire[993];							inform_R[993][3] = r_cell_wire[994];							inform_R[997][3] = r_cell_wire[995];							inform_R[994][3] = r_cell_wire[996];							inform_R[998][3] = r_cell_wire[997];							inform_R[995][3] = r_cell_wire[998];							inform_R[999][3] = r_cell_wire[999];							inform_R[1000][3] = r_cell_wire[1000];							inform_R[1004][3] = r_cell_wire[1001];							inform_R[1001][3] = r_cell_wire[1002];							inform_R[1005][3] = r_cell_wire[1003];							inform_R[1002][3] = r_cell_wire[1004];							inform_R[1006][3] = r_cell_wire[1005];							inform_R[1003][3] = r_cell_wire[1006];							inform_R[1007][3] = r_cell_wire[1007];							inform_R[1008][3] = r_cell_wire[1008];							inform_R[1012][3] = r_cell_wire[1009];							inform_R[1009][3] = r_cell_wire[1010];							inform_R[1013][3] = r_cell_wire[1011];							inform_R[1010][3] = r_cell_wire[1012];							inform_R[1014][3] = r_cell_wire[1013];							inform_R[1011][3] = r_cell_wire[1014];							inform_R[1015][3] = r_cell_wire[1015];							inform_R[1016][3] = r_cell_wire[1016];							inform_R[1020][3] = r_cell_wire[1017];							inform_R[1017][3] = r_cell_wire[1018];							inform_R[1021][3] = r_cell_wire[1019];							inform_R[1018][3] = r_cell_wire[1020];							inform_R[1022][3] = r_cell_wire[1021];							inform_R[1019][3] = r_cell_wire[1022];							inform_R[1023][3] = r_cell_wire[1023];							inform_L[0][2] = l_cell_wire[0];							inform_L[4][2] = l_cell_wire[1];							inform_L[1][2] = l_cell_wire[2];							inform_L[5][2] = l_cell_wire[3];							inform_L[2][2] = l_cell_wire[4];							inform_L[6][2] = l_cell_wire[5];							inform_L[3][2] = l_cell_wire[6];							inform_L[7][2] = l_cell_wire[7];							inform_L[8][2] = l_cell_wire[8];							inform_L[12][2] = l_cell_wire[9];							inform_L[9][2] = l_cell_wire[10];							inform_L[13][2] = l_cell_wire[11];							inform_L[10][2] = l_cell_wire[12];							inform_L[14][2] = l_cell_wire[13];							inform_L[11][2] = l_cell_wire[14];							inform_L[15][2] = l_cell_wire[15];							inform_L[16][2] = l_cell_wire[16];							inform_L[20][2] = l_cell_wire[17];							inform_L[17][2] = l_cell_wire[18];							inform_L[21][2] = l_cell_wire[19];							inform_L[18][2] = l_cell_wire[20];							inform_L[22][2] = l_cell_wire[21];							inform_L[19][2] = l_cell_wire[22];							inform_L[23][2] = l_cell_wire[23];							inform_L[24][2] = l_cell_wire[24];							inform_L[28][2] = l_cell_wire[25];							inform_L[25][2] = l_cell_wire[26];							inform_L[29][2] = l_cell_wire[27];							inform_L[26][2] = l_cell_wire[28];							inform_L[30][2] = l_cell_wire[29];							inform_L[27][2] = l_cell_wire[30];							inform_L[31][2] = l_cell_wire[31];							inform_L[32][2] = l_cell_wire[32];							inform_L[36][2] = l_cell_wire[33];							inform_L[33][2] = l_cell_wire[34];							inform_L[37][2] = l_cell_wire[35];							inform_L[34][2] = l_cell_wire[36];							inform_L[38][2] = l_cell_wire[37];							inform_L[35][2] = l_cell_wire[38];							inform_L[39][2] = l_cell_wire[39];							inform_L[40][2] = l_cell_wire[40];							inform_L[44][2] = l_cell_wire[41];							inform_L[41][2] = l_cell_wire[42];							inform_L[45][2] = l_cell_wire[43];							inform_L[42][2] = l_cell_wire[44];							inform_L[46][2] = l_cell_wire[45];							inform_L[43][2] = l_cell_wire[46];							inform_L[47][2] = l_cell_wire[47];							inform_L[48][2] = l_cell_wire[48];							inform_L[52][2] = l_cell_wire[49];							inform_L[49][2] = l_cell_wire[50];							inform_L[53][2] = l_cell_wire[51];							inform_L[50][2] = l_cell_wire[52];							inform_L[54][2] = l_cell_wire[53];							inform_L[51][2] = l_cell_wire[54];							inform_L[55][2] = l_cell_wire[55];							inform_L[56][2] = l_cell_wire[56];							inform_L[60][2] = l_cell_wire[57];							inform_L[57][2] = l_cell_wire[58];							inform_L[61][2] = l_cell_wire[59];							inform_L[58][2] = l_cell_wire[60];							inform_L[62][2] = l_cell_wire[61];							inform_L[59][2] = l_cell_wire[62];							inform_L[63][2] = l_cell_wire[63];							inform_L[64][2] = l_cell_wire[64];							inform_L[68][2] = l_cell_wire[65];							inform_L[65][2] = l_cell_wire[66];							inform_L[69][2] = l_cell_wire[67];							inform_L[66][2] = l_cell_wire[68];							inform_L[70][2] = l_cell_wire[69];							inform_L[67][2] = l_cell_wire[70];							inform_L[71][2] = l_cell_wire[71];							inform_L[72][2] = l_cell_wire[72];							inform_L[76][2] = l_cell_wire[73];							inform_L[73][2] = l_cell_wire[74];							inform_L[77][2] = l_cell_wire[75];							inform_L[74][2] = l_cell_wire[76];							inform_L[78][2] = l_cell_wire[77];							inform_L[75][2] = l_cell_wire[78];							inform_L[79][2] = l_cell_wire[79];							inform_L[80][2] = l_cell_wire[80];							inform_L[84][2] = l_cell_wire[81];							inform_L[81][2] = l_cell_wire[82];							inform_L[85][2] = l_cell_wire[83];							inform_L[82][2] = l_cell_wire[84];							inform_L[86][2] = l_cell_wire[85];							inform_L[83][2] = l_cell_wire[86];							inform_L[87][2] = l_cell_wire[87];							inform_L[88][2] = l_cell_wire[88];							inform_L[92][2] = l_cell_wire[89];							inform_L[89][2] = l_cell_wire[90];							inform_L[93][2] = l_cell_wire[91];							inform_L[90][2] = l_cell_wire[92];							inform_L[94][2] = l_cell_wire[93];							inform_L[91][2] = l_cell_wire[94];							inform_L[95][2] = l_cell_wire[95];							inform_L[96][2] = l_cell_wire[96];							inform_L[100][2] = l_cell_wire[97];							inform_L[97][2] = l_cell_wire[98];							inform_L[101][2] = l_cell_wire[99];							inform_L[98][2] = l_cell_wire[100];							inform_L[102][2] = l_cell_wire[101];							inform_L[99][2] = l_cell_wire[102];							inform_L[103][2] = l_cell_wire[103];							inform_L[104][2] = l_cell_wire[104];							inform_L[108][2] = l_cell_wire[105];							inform_L[105][2] = l_cell_wire[106];							inform_L[109][2] = l_cell_wire[107];							inform_L[106][2] = l_cell_wire[108];							inform_L[110][2] = l_cell_wire[109];							inform_L[107][2] = l_cell_wire[110];							inform_L[111][2] = l_cell_wire[111];							inform_L[112][2] = l_cell_wire[112];							inform_L[116][2] = l_cell_wire[113];							inform_L[113][2] = l_cell_wire[114];							inform_L[117][2] = l_cell_wire[115];							inform_L[114][2] = l_cell_wire[116];							inform_L[118][2] = l_cell_wire[117];							inform_L[115][2] = l_cell_wire[118];							inform_L[119][2] = l_cell_wire[119];							inform_L[120][2] = l_cell_wire[120];							inform_L[124][2] = l_cell_wire[121];							inform_L[121][2] = l_cell_wire[122];							inform_L[125][2] = l_cell_wire[123];							inform_L[122][2] = l_cell_wire[124];							inform_L[126][2] = l_cell_wire[125];							inform_L[123][2] = l_cell_wire[126];							inform_L[127][2] = l_cell_wire[127];							inform_L[128][2] = l_cell_wire[128];							inform_L[132][2] = l_cell_wire[129];							inform_L[129][2] = l_cell_wire[130];							inform_L[133][2] = l_cell_wire[131];							inform_L[130][2] = l_cell_wire[132];							inform_L[134][2] = l_cell_wire[133];							inform_L[131][2] = l_cell_wire[134];							inform_L[135][2] = l_cell_wire[135];							inform_L[136][2] = l_cell_wire[136];							inform_L[140][2] = l_cell_wire[137];							inform_L[137][2] = l_cell_wire[138];							inform_L[141][2] = l_cell_wire[139];							inform_L[138][2] = l_cell_wire[140];							inform_L[142][2] = l_cell_wire[141];							inform_L[139][2] = l_cell_wire[142];							inform_L[143][2] = l_cell_wire[143];							inform_L[144][2] = l_cell_wire[144];							inform_L[148][2] = l_cell_wire[145];							inform_L[145][2] = l_cell_wire[146];							inform_L[149][2] = l_cell_wire[147];							inform_L[146][2] = l_cell_wire[148];							inform_L[150][2] = l_cell_wire[149];							inform_L[147][2] = l_cell_wire[150];							inform_L[151][2] = l_cell_wire[151];							inform_L[152][2] = l_cell_wire[152];							inform_L[156][2] = l_cell_wire[153];							inform_L[153][2] = l_cell_wire[154];							inform_L[157][2] = l_cell_wire[155];							inform_L[154][2] = l_cell_wire[156];							inform_L[158][2] = l_cell_wire[157];							inform_L[155][2] = l_cell_wire[158];							inform_L[159][2] = l_cell_wire[159];							inform_L[160][2] = l_cell_wire[160];							inform_L[164][2] = l_cell_wire[161];							inform_L[161][2] = l_cell_wire[162];							inform_L[165][2] = l_cell_wire[163];							inform_L[162][2] = l_cell_wire[164];							inform_L[166][2] = l_cell_wire[165];							inform_L[163][2] = l_cell_wire[166];							inform_L[167][2] = l_cell_wire[167];							inform_L[168][2] = l_cell_wire[168];							inform_L[172][2] = l_cell_wire[169];							inform_L[169][2] = l_cell_wire[170];							inform_L[173][2] = l_cell_wire[171];							inform_L[170][2] = l_cell_wire[172];							inform_L[174][2] = l_cell_wire[173];							inform_L[171][2] = l_cell_wire[174];							inform_L[175][2] = l_cell_wire[175];							inform_L[176][2] = l_cell_wire[176];							inform_L[180][2] = l_cell_wire[177];							inform_L[177][2] = l_cell_wire[178];							inform_L[181][2] = l_cell_wire[179];							inform_L[178][2] = l_cell_wire[180];							inform_L[182][2] = l_cell_wire[181];							inform_L[179][2] = l_cell_wire[182];							inform_L[183][2] = l_cell_wire[183];							inform_L[184][2] = l_cell_wire[184];							inform_L[188][2] = l_cell_wire[185];							inform_L[185][2] = l_cell_wire[186];							inform_L[189][2] = l_cell_wire[187];							inform_L[186][2] = l_cell_wire[188];							inform_L[190][2] = l_cell_wire[189];							inform_L[187][2] = l_cell_wire[190];							inform_L[191][2] = l_cell_wire[191];							inform_L[192][2] = l_cell_wire[192];							inform_L[196][2] = l_cell_wire[193];							inform_L[193][2] = l_cell_wire[194];							inform_L[197][2] = l_cell_wire[195];							inform_L[194][2] = l_cell_wire[196];							inform_L[198][2] = l_cell_wire[197];							inform_L[195][2] = l_cell_wire[198];							inform_L[199][2] = l_cell_wire[199];							inform_L[200][2] = l_cell_wire[200];							inform_L[204][2] = l_cell_wire[201];							inform_L[201][2] = l_cell_wire[202];							inform_L[205][2] = l_cell_wire[203];							inform_L[202][2] = l_cell_wire[204];							inform_L[206][2] = l_cell_wire[205];							inform_L[203][2] = l_cell_wire[206];							inform_L[207][2] = l_cell_wire[207];							inform_L[208][2] = l_cell_wire[208];							inform_L[212][2] = l_cell_wire[209];							inform_L[209][2] = l_cell_wire[210];							inform_L[213][2] = l_cell_wire[211];							inform_L[210][2] = l_cell_wire[212];							inform_L[214][2] = l_cell_wire[213];							inform_L[211][2] = l_cell_wire[214];							inform_L[215][2] = l_cell_wire[215];							inform_L[216][2] = l_cell_wire[216];							inform_L[220][2] = l_cell_wire[217];							inform_L[217][2] = l_cell_wire[218];							inform_L[221][2] = l_cell_wire[219];							inform_L[218][2] = l_cell_wire[220];							inform_L[222][2] = l_cell_wire[221];							inform_L[219][2] = l_cell_wire[222];							inform_L[223][2] = l_cell_wire[223];							inform_L[224][2] = l_cell_wire[224];							inform_L[228][2] = l_cell_wire[225];							inform_L[225][2] = l_cell_wire[226];							inform_L[229][2] = l_cell_wire[227];							inform_L[226][2] = l_cell_wire[228];							inform_L[230][2] = l_cell_wire[229];							inform_L[227][2] = l_cell_wire[230];							inform_L[231][2] = l_cell_wire[231];							inform_L[232][2] = l_cell_wire[232];							inform_L[236][2] = l_cell_wire[233];							inform_L[233][2] = l_cell_wire[234];							inform_L[237][2] = l_cell_wire[235];							inform_L[234][2] = l_cell_wire[236];							inform_L[238][2] = l_cell_wire[237];							inform_L[235][2] = l_cell_wire[238];							inform_L[239][2] = l_cell_wire[239];							inform_L[240][2] = l_cell_wire[240];							inform_L[244][2] = l_cell_wire[241];							inform_L[241][2] = l_cell_wire[242];							inform_L[245][2] = l_cell_wire[243];							inform_L[242][2] = l_cell_wire[244];							inform_L[246][2] = l_cell_wire[245];							inform_L[243][2] = l_cell_wire[246];							inform_L[247][2] = l_cell_wire[247];							inform_L[248][2] = l_cell_wire[248];							inform_L[252][2] = l_cell_wire[249];							inform_L[249][2] = l_cell_wire[250];							inform_L[253][2] = l_cell_wire[251];							inform_L[250][2] = l_cell_wire[252];							inform_L[254][2] = l_cell_wire[253];							inform_L[251][2] = l_cell_wire[254];							inform_L[255][2] = l_cell_wire[255];							inform_L[256][2] = l_cell_wire[256];							inform_L[260][2] = l_cell_wire[257];							inform_L[257][2] = l_cell_wire[258];							inform_L[261][2] = l_cell_wire[259];							inform_L[258][2] = l_cell_wire[260];							inform_L[262][2] = l_cell_wire[261];							inform_L[259][2] = l_cell_wire[262];							inform_L[263][2] = l_cell_wire[263];							inform_L[264][2] = l_cell_wire[264];							inform_L[268][2] = l_cell_wire[265];							inform_L[265][2] = l_cell_wire[266];							inform_L[269][2] = l_cell_wire[267];							inform_L[266][2] = l_cell_wire[268];							inform_L[270][2] = l_cell_wire[269];							inform_L[267][2] = l_cell_wire[270];							inform_L[271][2] = l_cell_wire[271];							inform_L[272][2] = l_cell_wire[272];							inform_L[276][2] = l_cell_wire[273];							inform_L[273][2] = l_cell_wire[274];							inform_L[277][2] = l_cell_wire[275];							inform_L[274][2] = l_cell_wire[276];							inform_L[278][2] = l_cell_wire[277];							inform_L[275][2] = l_cell_wire[278];							inform_L[279][2] = l_cell_wire[279];							inform_L[280][2] = l_cell_wire[280];							inform_L[284][2] = l_cell_wire[281];							inform_L[281][2] = l_cell_wire[282];							inform_L[285][2] = l_cell_wire[283];							inform_L[282][2] = l_cell_wire[284];							inform_L[286][2] = l_cell_wire[285];							inform_L[283][2] = l_cell_wire[286];							inform_L[287][2] = l_cell_wire[287];							inform_L[288][2] = l_cell_wire[288];							inform_L[292][2] = l_cell_wire[289];							inform_L[289][2] = l_cell_wire[290];							inform_L[293][2] = l_cell_wire[291];							inform_L[290][2] = l_cell_wire[292];							inform_L[294][2] = l_cell_wire[293];							inform_L[291][2] = l_cell_wire[294];							inform_L[295][2] = l_cell_wire[295];							inform_L[296][2] = l_cell_wire[296];							inform_L[300][2] = l_cell_wire[297];							inform_L[297][2] = l_cell_wire[298];							inform_L[301][2] = l_cell_wire[299];							inform_L[298][2] = l_cell_wire[300];							inform_L[302][2] = l_cell_wire[301];							inform_L[299][2] = l_cell_wire[302];							inform_L[303][2] = l_cell_wire[303];							inform_L[304][2] = l_cell_wire[304];							inform_L[308][2] = l_cell_wire[305];							inform_L[305][2] = l_cell_wire[306];							inform_L[309][2] = l_cell_wire[307];							inform_L[306][2] = l_cell_wire[308];							inform_L[310][2] = l_cell_wire[309];							inform_L[307][2] = l_cell_wire[310];							inform_L[311][2] = l_cell_wire[311];							inform_L[312][2] = l_cell_wire[312];							inform_L[316][2] = l_cell_wire[313];							inform_L[313][2] = l_cell_wire[314];							inform_L[317][2] = l_cell_wire[315];							inform_L[314][2] = l_cell_wire[316];							inform_L[318][2] = l_cell_wire[317];							inform_L[315][2] = l_cell_wire[318];							inform_L[319][2] = l_cell_wire[319];							inform_L[320][2] = l_cell_wire[320];							inform_L[324][2] = l_cell_wire[321];							inform_L[321][2] = l_cell_wire[322];							inform_L[325][2] = l_cell_wire[323];							inform_L[322][2] = l_cell_wire[324];							inform_L[326][2] = l_cell_wire[325];							inform_L[323][2] = l_cell_wire[326];							inform_L[327][2] = l_cell_wire[327];							inform_L[328][2] = l_cell_wire[328];							inform_L[332][2] = l_cell_wire[329];							inform_L[329][2] = l_cell_wire[330];							inform_L[333][2] = l_cell_wire[331];							inform_L[330][2] = l_cell_wire[332];							inform_L[334][2] = l_cell_wire[333];							inform_L[331][2] = l_cell_wire[334];							inform_L[335][2] = l_cell_wire[335];							inform_L[336][2] = l_cell_wire[336];							inform_L[340][2] = l_cell_wire[337];							inform_L[337][2] = l_cell_wire[338];							inform_L[341][2] = l_cell_wire[339];							inform_L[338][2] = l_cell_wire[340];							inform_L[342][2] = l_cell_wire[341];							inform_L[339][2] = l_cell_wire[342];							inform_L[343][2] = l_cell_wire[343];							inform_L[344][2] = l_cell_wire[344];							inform_L[348][2] = l_cell_wire[345];							inform_L[345][2] = l_cell_wire[346];							inform_L[349][2] = l_cell_wire[347];							inform_L[346][2] = l_cell_wire[348];							inform_L[350][2] = l_cell_wire[349];							inform_L[347][2] = l_cell_wire[350];							inform_L[351][2] = l_cell_wire[351];							inform_L[352][2] = l_cell_wire[352];							inform_L[356][2] = l_cell_wire[353];							inform_L[353][2] = l_cell_wire[354];							inform_L[357][2] = l_cell_wire[355];							inform_L[354][2] = l_cell_wire[356];							inform_L[358][2] = l_cell_wire[357];							inform_L[355][2] = l_cell_wire[358];							inform_L[359][2] = l_cell_wire[359];							inform_L[360][2] = l_cell_wire[360];							inform_L[364][2] = l_cell_wire[361];							inform_L[361][2] = l_cell_wire[362];							inform_L[365][2] = l_cell_wire[363];							inform_L[362][2] = l_cell_wire[364];							inform_L[366][2] = l_cell_wire[365];							inform_L[363][2] = l_cell_wire[366];							inform_L[367][2] = l_cell_wire[367];							inform_L[368][2] = l_cell_wire[368];							inform_L[372][2] = l_cell_wire[369];							inform_L[369][2] = l_cell_wire[370];							inform_L[373][2] = l_cell_wire[371];							inform_L[370][2] = l_cell_wire[372];							inform_L[374][2] = l_cell_wire[373];							inform_L[371][2] = l_cell_wire[374];							inform_L[375][2] = l_cell_wire[375];							inform_L[376][2] = l_cell_wire[376];							inform_L[380][2] = l_cell_wire[377];							inform_L[377][2] = l_cell_wire[378];							inform_L[381][2] = l_cell_wire[379];							inform_L[378][2] = l_cell_wire[380];							inform_L[382][2] = l_cell_wire[381];							inform_L[379][2] = l_cell_wire[382];							inform_L[383][2] = l_cell_wire[383];							inform_L[384][2] = l_cell_wire[384];							inform_L[388][2] = l_cell_wire[385];							inform_L[385][2] = l_cell_wire[386];							inform_L[389][2] = l_cell_wire[387];							inform_L[386][2] = l_cell_wire[388];							inform_L[390][2] = l_cell_wire[389];							inform_L[387][2] = l_cell_wire[390];							inform_L[391][2] = l_cell_wire[391];							inform_L[392][2] = l_cell_wire[392];							inform_L[396][2] = l_cell_wire[393];							inform_L[393][2] = l_cell_wire[394];							inform_L[397][2] = l_cell_wire[395];							inform_L[394][2] = l_cell_wire[396];							inform_L[398][2] = l_cell_wire[397];							inform_L[395][2] = l_cell_wire[398];							inform_L[399][2] = l_cell_wire[399];							inform_L[400][2] = l_cell_wire[400];							inform_L[404][2] = l_cell_wire[401];							inform_L[401][2] = l_cell_wire[402];							inform_L[405][2] = l_cell_wire[403];							inform_L[402][2] = l_cell_wire[404];							inform_L[406][2] = l_cell_wire[405];							inform_L[403][2] = l_cell_wire[406];							inform_L[407][2] = l_cell_wire[407];							inform_L[408][2] = l_cell_wire[408];							inform_L[412][2] = l_cell_wire[409];							inform_L[409][2] = l_cell_wire[410];							inform_L[413][2] = l_cell_wire[411];							inform_L[410][2] = l_cell_wire[412];							inform_L[414][2] = l_cell_wire[413];							inform_L[411][2] = l_cell_wire[414];							inform_L[415][2] = l_cell_wire[415];							inform_L[416][2] = l_cell_wire[416];							inform_L[420][2] = l_cell_wire[417];							inform_L[417][2] = l_cell_wire[418];							inform_L[421][2] = l_cell_wire[419];							inform_L[418][2] = l_cell_wire[420];							inform_L[422][2] = l_cell_wire[421];							inform_L[419][2] = l_cell_wire[422];							inform_L[423][2] = l_cell_wire[423];							inform_L[424][2] = l_cell_wire[424];							inform_L[428][2] = l_cell_wire[425];							inform_L[425][2] = l_cell_wire[426];							inform_L[429][2] = l_cell_wire[427];							inform_L[426][2] = l_cell_wire[428];							inform_L[430][2] = l_cell_wire[429];							inform_L[427][2] = l_cell_wire[430];							inform_L[431][2] = l_cell_wire[431];							inform_L[432][2] = l_cell_wire[432];							inform_L[436][2] = l_cell_wire[433];							inform_L[433][2] = l_cell_wire[434];							inform_L[437][2] = l_cell_wire[435];							inform_L[434][2] = l_cell_wire[436];							inform_L[438][2] = l_cell_wire[437];							inform_L[435][2] = l_cell_wire[438];							inform_L[439][2] = l_cell_wire[439];							inform_L[440][2] = l_cell_wire[440];							inform_L[444][2] = l_cell_wire[441];							inform_L[441][2] = l_cell_wire[442];							inform_L[445][2] = l_cell_wire[443];							inform_L[442][2] = l_cell_wire[444];							inform_L[446][2] = l_cell_wire[445];							inform_L[443][2] = l_cell_wire[446];							inform_L[447][2] = l_cell_wire[447];							inform_L[448][2] = l_cell_wire[448];							inform_L[452][2] = l_cell_wire[449];							inform_L[449][2] = l_cell_wire[450];							inform_L[453][2] = l_cell_wire[451];							inform_L[450][2] = l_cell_wire[452];							inform_L[454][2] = l_cell_wire[453];							inform_L[451][2] = l_cell_wire[454];							inform_L[455][2] = l_cell_wire[455];							inform_L[456][2] = l_cell_wire[456];							inform_L[460][2] = l_cell_wire[457];							inform_L[457][2] = l_cell_wire[458];							inform_L[461][2] = l_cell_wire[459];							inform_L[458][2] = l_cell_wire[460];							inform_L[462][2] = l_cell_wire[461];							inform_L[459][2] = l_cell_wire[462];							inform_L[463][2] = l_cell_wire[463];							inform_L[464][2] = l_cell_wire[464];							inform_L[468][2] = l_cell_wire[465];							inform_L[465][2] = l_cell_wire[466];							inform_L[469][2] = l_cell_wire[467];							inform_L[466][2] = l_cell_wire[468];							inform_L[470][2] = l_cell_wire[469];							inform_L[467][2] = l_cell_wire[470];							inform_L[471][2] = l_cell_wire[471];							inform_L[472][2] = l_cell_wire[472];							inform_L[476][2] = l_cell_wire[473];							inform_L[473][2] = l_cell_wire[474];							inform_L[477][2] = l_cell_wire[475];							inform_L[474][2] = l_cell_wire[476];							inform_L[478][2] = l_cell_wire[477];							inform_L[475][2] = l_cell_wire[478];							inform_L[479][2] = l_cell_wire[479];							inform_L[480][2] = l_cell_wire[480];							inform_L[484][2] = l_cell_wire[481];							inform_L[481][2] = l_cell_wire[482];							inform_L[485][2] = l_cell_wire[483];							inform_L[482][2] = l_cell_wire[484];							inform_L[486][2] = l_cell_wire[485];							inform_L[483][2] = l_cell_wire[486];							inform_L[487][2] = l_cell_wire[487];							inform_L[488][2] = l_cell_wire[488];							inform_L[492][2] = l_cell_wire[489];							inform_L[489][2] = l_cell_wire[490];							inform_L[493][2] = l_cell_wire[491];							inform_L[490][2] = l_cell_wire[492];							inform_L[494][2] = l_cell_wire[493];							inform_L[491][2] = l_cell_wire[494];							inform_L[495][2] = l_cell_wire[495];							inform_L[496][2] = l_cell_wire[496];							inform_L[500][2] = l_cell_wire[497];							inform_L[497][2] = l_cell_wire[498];							inform_L[501][2] = l_cell_wire[499];							inform_L[498][2] = l_cell_wire[500];							inform_L[502][2] = l_cell_wire[501];							inform_L[499][2] = l_cell_wire[502];							inform_L[503][2] = l_cell_wire[503];							inform_L[504][2] = l_cell_wire[504];							inform_L[508][2] = l_cell_wire[505];							inform_L[505][2] = l_cell_wire[506];							inform_L[509][2] = l_cell_wire[507];							inform_L[506][2] = l_cell_wire[508];							inform_L[510][2] = l_cell_wire[509];							inform_L[507][2] = l_cell_wire[510];							inform_L[511][2] = l_cell_wire[511];							inform_L[512][2] = l_cell_wire[512];							inform_L[516][2] = l_cell_wire[513];							inform_L[513][2] = l_cell_wire[514];							inform_L[517][2] = l_cell_wire[515];							inform_L[514][2] = l_cell_wire[516];							inform_L[518][2] = l_cell_wire[517];							inform_L[515][2] = l_cell_wire[518];							inform_L[519][2] = l_cell_wire[519];							inform_L[520][2] = l_cell_wire[520];							inform_L[524][2] = l_cell_wire[521];							inform_L[521][2] = l_cell_wire[522];							inform_L[525][2] = l_cell_wire[523];							inform_L[522][2] = l_cell_wire[524];							inform_L[526][2] = l_cell_wire[525];							inform_L[523][2] = l_cell_wire[526];							inform_L[527][2] = l_cell_wire[527];							inform_L[528][2] = l_cell_wire[528];							inform_L[532][2] = l_cell_wire[529];							inform_L[529][2] = l_cell_wire[530];							inform_L[533][2] = l_cell_wire[531];							inform_L[530][2] = l_cell_wire[532];							inform_L[534][2] = l_cell_wire[533];							inform_L[531][2] = l_cell_wire[534];							inform_L[535][2] = l_cell_wire[535];							inform_L[536][2] = l_cell_wire[536];							inform_L[540][2] = l_cell_wire[537];							inform_L[537][2] = l_cell_wire[538];							inform_L[541][2] = l_cell_wire[539];							inform_L[538][2] = l_cell_wire[540];							inform_L[542][2] = l_cell_wire[541];							inform_L[539][2] = l_cell_wire[542];							inform_L[543][2] = l_cell_wire[543];							inform_L[544][2] = l_cell_wire[544];							inform_L[548][2] = l_cell_wire[545];							inform_L[545][2] = l_cell_wire[546];							inform_L[549][2] = l_cell_wire[547];							inform_L[546][2] = l_cell_wire[548];							inform_L[550][2] = l_cell_wire[549];							inform_L[547][2] = l_cell_wire[550];							inform_L[551][2] = l_cell_wire[551];							inform_L[552][2] = l_cell_wire[552];							inform_L[556][2] = l_cell_wire[553];							inform_L[553][2] = l_cell_wire[554];							inform_L[557][2] = l_cell_wire[555];							inform_L[554][2] = l_cell_wire[556];							inform_L[558][2] = l_cell_wire[557];							inform_L[555][2] = l_cell_wire[558];							inform_L[559][2] = l_cell_wire[559];							inform_L[560][2] = l_cell_wire[560];							inform_L[564][2] = l_cell_wire[561];							inform_L[561][2] = l_cell_wire[562];							inform_L[565][2] = l_cell_wire[563];							inform_L[562][2] = l_cell_wire[564];							inform_L[566][2] = l_cell_wire[565];							inform_L[563][2] = l_cell_wire[566];							inform_L[567][2] = l_cell_wire[567];							inform_L[568][2] = l_cell_wire[568];							inform_L[572][2] = l_cell_wire[569];							inform_L[569][2] = l_cell_wire[570];							inform_L[573][2] = l_cell_wire[571];							inform_L[570][2] = l_cell_wire[572];							inform_L[574][2] = l_cell_wire[573];							inform_L[571][2] = l_cell_wire[574];							inform_L[575][2] = l_cell_wire[575];							inform_L[576][2] = l_cell_wire[576];							inform_L[580][2] = l_cell_wire[577];							inform_L[577][2] = l_cell_wire[578];							inform_L[581][2] = l_cell_wire[579];							inform_L[578][2] = l_cell_wire[580];							inform_L[582][2] = l_cell_wire[581];							inform_L[579][2] = l_cell_wire[582];							inform_L[583][2] = l_cell_wire[583];							inform_L[584][2] = l_cell_wire[584];							inform_L[588][2] = l_cell_wire[585];							inform_L[585][2] = l_cell_wire[586];							inform_L[589][2] = l_cell_wire[587];							inform_L[586][2] = l_cell_wire[588];							inform_L[590][2] = l_cell_wire[589];							inform_L[587][2] = l_cell_wire[590];							inform_L[591][2] = l_cell_wire[591];							inform_L[592][2] = l_cell_wire[592];							inform_L[596][2] = l_cell_wire[593];							inform_L[593][2] = l_cell_wire[594];							inform_L[597][2] = l_cell_wire[595];							inform_L[594][2] = l_cell_wire[596];							inform_L[598][2] = l_cell_wire[597];							inform_L[595][2] = l_cell_wire[598];							inform_L[599][2] = l_cell_wire[599];							inform_L[600][2] = l_cell_wire[600];							inform_L[604][2] = l_cell_wire[601];							inform_L[601][2] = l_cell_wire[602];							inform_L[605][2] = l_cell_wire[603];							inform_L[602][2] = l_cell_wire[604];							inform_L[606][2] = l_cell_wire[605];							inform_L[603][2] = l_cell_wire[606];							inform_L[607][2] = l_cell_wire[607];							inform_L[608][2] = l_cell_wire[608];							inform_L[612][2] = l_cell_wire[609];							inform_L[609][2] = l_cell_wire[610];							inform_L[613][2] = l_cell_wire[611];							inform_L[610][2] = l_cell_wire[612];							inform_L[614][2] = l_cell_wire[613];							inform_L[611][2] = l_cell_wire[614];							inform_L[615][2] = l_cell_wire[615];							inform_L[616][2] = l_cell_wire[616];							inform_L[620][2] = l_cell_wire[617];							inform_L[617][2] = l_cell_wire[618];							inform_L[621][2] = l_cell_wire[619];							inform_L[618][2] = l_cell_wire[620];							inform_L[622][2] = l_cell_wire[621];							inform_L[619][2] = l_cell_wire[622];							inform_L[623][2] = l_cell_wire[623];							inform_L[624][2] = l_cell_wire[624];							inform_L[628][2] = l_cell_wire[625];							inform_L[625][2] = l_cell_wire[626];							inform_L[629][2] = l_cell_wire[627];							inform_L[626][2] = l_cell_wire[628];							inform_L[630][2] = l_cell_wire[629];							inform_L[627][2] = l_cell_wire[630];							inform_L[631][2] = l_cell_wire[631];							inform_L[632][2] = l_cell_wire[632];							inform_L[636][2] = l_cell_wire[633];							inform_L[633][2] = l_cell_wire[634];							inform_L[637][2] = l_cell_wire[635];							inform_L[634][2] = l_cell_wire[636];							inform_L[638][2] = l_cell_wire[637];							inform_L[635][2] = l_cell_wire[638];							inform_L[639][2] = l_cell_wire[639];							inform_L[640][2] = l_cell_wire[640];							inform_L[644][2] = l_cell_wire[641];							inform_L[641][2] = l_cell_wire[642];							inform_L[645][2] = l_cell_wire[643];							inform_L[642][2] = l_cell_wire[644];							inform_L[646][2] = l_cell_wire[645];							inform_L[643][2] = l_cell_wire[646];							inform_L[647][2] = l_cell_wire[647];							inform_L[648][2] = l_cell_wire[648];							inform_L[652][2] = l_cell_wire[649];							inform_L[649][2] = l_cell_wire[650];							inform_L[653][2] = l_cell_wire[651];							inform_L[650][2] = l_cell_wire[652];							inform_L[654][2] = l_cell_wire[653];							inform_L[651][2] = l_cell_wire[654];							inform_L[655][2] = l_cell_wire[655];							inform_L[656][2] = l_cell_wire[656];							inform_L[660][2] = l_cell_wire[657];							inform_L[657][2] = l_cell_wire[658];							inform_L[661][2] = l_cell_wire[659];							inform_L[658][2] = l_cell_wire[660];							inform_L[662][2] = l_cell_wire[661];							inform_L[659][2] = l_cell_wire[662];							inform_L[663][2] = l_cell_wire[663];							inform_L[664][2] = l_cell_wire[664];							inform_L[668][2] = l_cell_wire[665];							inform_L[665][2] = l_cell_wire[666];							inform_L[669][2] = l_cell_wire[667];							inform_L[666][2] = l_cell_wire[668];							inform_L[670][2] = l_cell_wire[669];							inform_L[667][2] = l_cell_wire[670];							inform_L[671][2] = l_cell_wire[671];							inform_L[672][2] = l_cell_wire[672];							inform_L[676][2] = l_cell_wire[673];							inform_L[673][2] = l_cell_wire[674];							inform_L[677][2] = l_cell_wire[675];							inform_L[674][2] = l_cell_wire[676];							inform_L[678][2] = l_cell_wire[677];							inform_L[675][2] = l_cell_wire[678];							inform_L[679][2] = l_cell_wire[679];							inform_L[680][2] = l_cell_wire[680];							inform_L[684][2] = l_cell_wire[681];							inform_L[681][2] = l_cell_wire[682];							inform_L[685][2] = l_cell_wire[683];							inform_L[682][2] = l_cell_wire[684];							inform_L[686][2] = l_cell_wire[685];							inform_L[683][2] = l_cell_wire[686];							inform_L[687][2] = l_cell_wire[687];							inform_L[688][2] = l_cell_wire[688];							inform_L[692][2] = l_cell_wire[689];							inform_L[689][2] = l_cell_wire[690];							inform_L[693][2] = l_cell_wire[691];							inform_L[690][2] = l_cell_wire[692];							inform_L[694][2] = l_cell_wire[693];							inform_L[691][2] = l_cell_wire[694];							inform_L[695][2] = l_cell_wire[695];							inform_L[696][2] = l_cell_wire[696];							inform_L[700][2] = l_cell_wire[697];							inform_L[697][2] = l_cell_wire[698];							inform_L[701][2] = l_cell_wire[699];							inform_L[698][2] = l_cell_wire[700];							inform_L[702][2] = l_cell_wire[701];							inform_L[699][2] = l_cell_wire[702];							inform_L[703][2] = l_cell_wire[703];							inform_L[704][2] = l_cell_wire[704];							inform_L[708][2] = l_cell_wire[705];							inform_L[705][2] = l_cell_wire[706];							inform_L[709][2] = l_cell_wire[707];							inform_L[706][2] = l_cell_wire[708];							inform_L[710][2] = l_cell_wire[709];							inform_L[707][2] = l_cell_wire[710];							inform_L[711][2] = l_cell_wire[711];							inform_L[712][2] = l_cell_wire[712];							inform_L[716][2] = l_cell_wire[713];							inform_L[713][2] = l_cell_wire[714];							inform_L[717][2] = l_cell_wire[715];							inform_L[714][2] = l_cell_wire[716];							inform_L[718][2] = l_cell_wire[717];							inform_L[715][2] = l_cell_wire[718];							inform_L[719][2] = l_cell_wire[719];							inform_L[720][2] = l_cell_wire[720];							inform_L[724][2] = l_cell_wire[721];							inform_L[721][2] = l_cell_wire[722];							inform_L[725][2] = l_cell_wire[723];							inform_L[722][2] = l_cell_wire[724];							inform_L[726][2] = l_cell_wire[725];							inform_L[723][2] = l_cell_wire[726];							inform_L[727][2] = l_cell_wire[727];							inform_L[728][2] = l_cell_wire[728];							inform_L[732][2] = l_cell_wire[729];							inform_L[729][2] = l_cell_wire[730];							inform_L[733][2] = l_cell_wire[731];							inform_L[730][2] = l_cell_wire[732];							inform_L[734][2] = l_cell_wire[733];							inform_L[731][2] = l_cell_wire[734];							inform_L[735][2] = l_cell_wire[735];							inform_L[736][2] = l_cell_wire[736];							inform_L[740][2] = l_cell_wire[737];							inform_L[737][2] = l_cell_wire[738];							inform_L[741][2] = l_cell_wire[739];							inform_L[738][2] = l_cell_wire[740];							inform_L[742][2] = l_cell_wire[741];							inform_L[739][2] = l_cell_wire[742];							inform_L[743][2] = l_cell_wire[743];							inform_L[744][2] = l_cell_wire[744];							inform_L[748][2] = l_cell_wire[745];							inform_L[745][2] = l_cell_wire[746];							inform_L[749][2] = l_cell_wire[747];							inform_L[746][2] = l_cell_wire[748];							inform_L[750][2] = l_cell_wire[749];							inform_L[747][2] = l_cell_wire[750];							inform_L[751][2] = l_cell_wire[751];							inform_L[752][2] = l_cell_wire[752];							inform_L[756][2] = l_cell_wire[753];							inform_L[753][2] = l_cell_wire[754];							inform_L[757][2] = l_cell_wire[755];							inform_L[754][2] = l_cell_wire[756];							inform_L[758][2] = l_cell_wire[757];							inform_L[755][2] = l_cell_wire[758];							inform_L[759][2] = l_cell_wire[759];							inform_L[760][2] = l_cell_wire[760];							inform_L[764][2] = l_cell_wire[761];							inform_L[761][2] = l_cell_wire[762];							inform_L[765][2] = l_cell_wire[763];							inform_L[762][2] = l_cell_wire[764];							inform_L[766][2] = l_cell_wire[765];							inform_L[763][2] = l_cell_wire[766];							inform_L[767][2] = l_cell_wire[767];							inform_L[768][2] = l_cell_wire[768];							inform_L[772][2] = l_cell_wire[769];							inform_L[769][2] = l_cell_wire[770];							inform_L[773][2] = l_cell_wire[771];							inform_L[770][2] = l_cell_wire[772];							inform_L[774][2] = l_cell_wire[773];							inform_L[771][2] = l_cell_wire[774];							inform_L[775][2] = l_cell_wire[775];							inform_L[776][2] = l_cell_wire[776];							inform_L[780][2] = l_cell_wire[777];							inform_L[777][2] = l_cell_wire[778];							inform_L[781][2] = l_cell_wire[779];							inform_L[778][2] = l_cell_wire[780];							inform_L[782][2] = l_cell_wire[781];							inform_L[779][2] = l_cell_wire[782];							inform_L[783][2] = l_cell_wire[783];							inform_L[784][2] = l_cell_wire[784];							inform_L[788][2] = l_cell_wire[785];							inform_L[785][2] = l_cell_wire[786];							inform_L[789][2] = l_cell_wire[787];							inform_L[786][2] = l_cell_wire[788];							inform_L[790][2] = l_cell_wire[789];							inform_L[787][2] = l_cell_wire[790];							inform_L[791][2] = l_cell_wire[791];							inform_L[792][2] = l_cell_wire[792];							inform_L[796][2] = l_cell_wire[793];							inform_L[793][2] = l_cell_wire[794];							inform_L[797][2] = l_cell_wire[795];							inform_L[794][2] = l_cell_wire[796];							inform_L[798][2] = l_cell_wire[797];							inform_L[795][2] = l_cell_wire[798];							inform_L[799][2] = l_cell_wire[799];							inform_L[800][2] = l_cell_wire[800];							inform_L[804][2] = l_cell_wire[801];							inform_L[801][2] = l_cell_wire[802];							inform_L[805][2] = l_cell_wire[803];							inform_L[802][2] = l_cell_wire[804];							inform_L[806][2] = l_cell_wire[805];							inform_L[803][2] = l_cell_wire[806];							inform_L[807][2] = l_cell_wire[807];							inform_L[808][2] = l_cell_wire[808];							inform_L[812][2] = l_cell_wire[809];							inform_L[809][2] = l_cell_wire[810];							inform_L[813][2] = l_cell_wire[811];							inform_L[810][2] = l_cell_wire[812];							inform_L[814][2] = l_cell_wire[813];							inform_L[811][2] = l_cell_wire[814];							inform_L[815][2] = l_cell_wire[815];							inform_L[816][2] = l_cell_wire[816];							inform_L[820][2] = l_cell_wire[817];							inform_L[817][2] = l_cell_wire[818];							inform_L[821][2] = l_cell_wire[819];							inform_L[818][2] = l_cell_wire[820];							inform_L[822][2] = l_cell_wire[821];							inform_L[819][2] = l_cell_wire[822];							inform_L[823][2] = l_cell_wire[823];							inform_L[824][2] = l_cell_wire[824];							inform_L[828][2] = l_cell_wire[825];							inform_L[825][2] = l_cell_wire[826];							inform_L[829][2] = l_cell_wire[827];							inform_L[826][2] = l_cell_wire[828];							inform_L[830][2] = l_cell_wire[829];							inform_L[827][2] = l_cell_wire[830];							inform_L[831][2] = l_cell_wire[831];							inform_L[832][2] = l_cell_wire[832];							inform_L[836][2] = l_cell_wire[833];							inform_L[833][2] = l_cell_wire[834];							inform_L[837][2] = l_cell_wire[835];							inform_L[834][2] = l_cell_wire[836];							inform_L[838][2] = l_cell_wire[837];							inform_L[835][2] = l_cell_wire[838];							inform_L[839][2] = l_cell_wire[839];							inform_L[840][2] = l_cell_wire[840];							inform_L[844][2] = l_cell_wire[841];							inform_L[841][2] = l_cell_wire[842];							inform_L[845][2] = l_cell_wire[843];							inform_L[842][2] = l_cell_wire[844];							inform_L[846][2] = l_cell_wire[845];							inform_L[843][2] = l_cell_wire[846];							inform_L[847][2] = l_cell_wire[847];							inform_L[848][2] = l_cell_wire[848];							inform_L[852][2] = l_cell_wire[849];							inform_L[849][2] = l_cell_wire[850];							inform_L[853][2] = l_cell_wire[851];							inform_L[850][2] = l_cell_wire[852];							inform_L[854][2] = l_cell_wire[853];							inform_L[851][2] = l_cell_wire[854];							inform_L[855][2] = l_cell_wire[855];							inform_L[856][2] = l_cell_wire[856];							inform_L[860][2] = l_cell_wire[857];							inform_L[857][2] = l_cell_wire[858];							inform_L[861][2] = l_cell_wire[859];							inform_L[858][2] = l_cell_wire[860];							inform_L[862][2] = l_cell_wire[861];							inform_L[859][2] = l_cell_wire[862];							inform_L[863][2] = l_cell_wire[863];							inform_L[864][2] = l_cell_wire[864];							inform_L[868][2] = l_cell_wire[865];							inform_L[865][2] = l_cell_wire[866];							inform_L[869][2] = l_cell_wire[867];							inform_L[866][2] = l_cell_wire[868];							inform_L[870][2] = l_cell_wire[869];							inform_L[867][2] = l_cell_wire[870];							inform_L[871][2] = l_cell_wire[871];							inform_L[872][2] = l_cell_wire[872];							inform_L[876][2] = l_cell_wire[873];							inform_L[873][2] = l_cell_wire[874];							inform_L[877][2] = l_cell_wire[875];							inform_L[874][2] = l_cell_wire[876];							inform_L[878][2] = l_cell_wire[877];							inform_L[875][2] = l_cell_wire[878];							inform_L[879][2] = l_cell_wire[879];							inform_L[880][2] = l_cell_wire[880];							inform_L[884][2] = l_cell_wire[881];							inform_L[881][2] = l_cell_wire[882];							inform_L[885][2] = l_cell_wire[883];							inform_L[882][2] = l_cell_wire[884];							inform_L[886][2] = l_cell_wire[885];							inform_L[883][2] = l_cell_wire[886];							inform_L[887][2] = l_cell_wire[887];							inform_L[888][2] = l_cell_wire[888];							inform_L[892][2] = l_cell_wire[889];							inform_L[889][2] = l_cell_wire[890];							inform_L[893][2] = l_cell_wire[891];							inform_L[890][2] = l_cell_wire[892];							inform_L[894][2] = l_cell_wire[893];							inform_L[891][2] = l_cell_wire[894];							inform_L[895][2] = l_cell_wire[895];							inform_L[896][2] = l_cell_wire[896];							inform_L[900][2] = l_cell_wire[897];							inform_L[897][2] = l_cell_wire[898];							inform_L[901][2] = l_cell_wire[899];							inform_L[898][2] = l_cell_wire[900];							inform_L[902][2] = l_cell_wire[901];							inform_L[899][2] = l_cell_wire[902];							inform_L[903][2] = l_cell_wire[903];							inform_L[904][2] = l_cell_wire[904];							inform_L[908][2] = l_cell_wire[905];							inform_L[905][2] = l_cell_wire[906];							inform_L[909][2] = l_cell_wire[907];							inform_L[906][2] = l_cell_wire[908];							inform_L[910][2] = l_cell_wire[909];							inform_L[907][2] = l_cell_wire[910];							inform_L[911][2] = l_cell_wire[911];							inform_L[912][2] = l_cell_wire[912];							inform_L[916][2] = l_cell_wire[913];							inform_L[913][2] = l_cell_wire[914];							inform_L[917][2] = l_cell_wire[915];							inform_L[914][2] = l_cell_wire[916];							inform_L[918][2] = l_cell_wire[917];							inform_L[915][2] = l_cell_wire[918];							inform_L[919][2] = l_cell_wire[919];							inform_L[920][2] = l_cell_wire[920];							inform_L[924][2] = l_cell_wire[921];							inform_L[921][2] = l_cell_wire[922];							inform_L[925][2] = l_cell_wire[923];							inform_L[922][2] = l_cell_wire[924];							inform_L[926][2] = l_cell_wire[925];							inform_L[923][2] = l_cell_wire[926];							inform_L[927][2] = l_cell_wire[927];							inform_L[928][2] = l_cell_wire[928];							inform_L[932][2] = l_cell_wire[929];							inform_L[929][2] = l_cell_wire[930];							inform_L[933][2] = l_cell_wire[931];							inform_L[930][2] = l_cell_wire[932];							inform_L[934][2] = l_cell_wire[933];							inform_L[931][2] = l_cell_wire[934];							inform_L[935][2] = l_cell_wire[935];							inform_L[936][2] = l_cell_wire[936];							inform_L[940][2] = l_cell_wire[937];							inform_L[937][2] = l_cell_wire[938];							inform_L[941][2] = l_cell_wire[939];							inform_L[938][2] = l_cell_wire[940];							inform_L[942][2] = l_cell_wire[941];							inform_L[939][2] = l_cell_wire[942];							inform_L[943][2] = l_cell_wire[943];							inform_L[944][2] = l_cell_wire[944];							inform_L[948][2] = l_cell_wire[945];							inform_L[945][2] = l_cell_wire[946];							inform_L[949][2] = l_cell_wire[947];							inform_L[946][2] = l_cell_wire[948];							inform_L[950][2] = l_cell_wire[949];							inform_L[947][2] = l_cell_wire[950];							inform_L[951][2] = l_cell_wire[951];							inform_L[952][2] = l_cell_wire[952];							inform_L[956][2] = l_cell_wire[953];							inform_L[953][2] = l_cell_wire[954];							inform_L[957][2] = l_cell_wire[955];							inform_L[954][2] = l_cell_wire[956];							inform_L[958][2] = l_cell_wire[957];							inform_L[955][2] = l_cell_wire[958];							inform_L[959][2] = l_cell_wire[959];							inform_L[960][2] = l_cell_wire[960];							inform_L[964][2] = l_cell_wire[961];							inform_L[961][2] = l_cell_wire[962];							inform_L[965][2] = l_cell_wire[963];							inform_L[962][2] = l_cell_wire[964];							inform_L[966][2] = l_cell_wire[965];							inform_L[963][2] = l_cell_wire[966];							inform_L[967][2] = l_cell_wire[967];							inform_L[968][2] = l_cell_wire[968];							inform_L[972][2] = l_cell_wire[969];							inform_L[969][2] = l_cell_wire[970];							inform_L[973][2] = l_cell_wire[971];							inform_L[970][2] = l_cell_wire[972];							inform_L[974][2] = l_cell_wire[973];							inform_L[971][2] = l_cell_wire[974];							inform_L[975][2] = l_cell_wire[975];							inform_L[976][2] = l_cell_wire[976];							inform_L[980][2] = l_cell_wire[977];							inform_L[977][2] = l_cell_wire[978];							inform_L[981][2] = l_cell_wire[979];							inform_L[978][2] = l_cell_wire[980];							inform_L[982][2] = l_cell_wire[981];							inform_L[979][2] = l_cell_wire[982];							inform_L[983][2] = l_cell_wire[983];							inform_L[984][2] = l_cell_wire[984];							inform_L[988][2] = l_cell_wire[985];							inform_L[985][2] = l_cell_wire[986];							inform_L[989][2] = l_cell_wire[987];							inform_L[986][2] = l_cell_wire[988];							inform_L[990][2] = l_cell_wire[989];							inform_L[987][2] = l_cell_wire[990];							inform_L[991][2] = l_cell_wire[991];							inform_L[992][2] = l_cell_wire[992];							inform_L[996][2] = l_cell_wire[993];							inform_L[993][2] = l_cell_wire[994];							inform_L[997][2] = l_cell_wire[995];							inform_L[994][2] = l_cell_wire[996];							inform_L[998][2] = l_cell_wire[997];							inform_L[995][2] = l_cell_wire[998];							inform_L[999][2] = l_cell_wire[999];							inform_L[1000][2] = l_cell_wire[1000];							inform_L[1004][2] = l_cell_wire[1001];							inform_L[1001][2] = l_cell_wire[1002];							inform_L[1005][2] = l_cell_wire[1003];							inform_L[1002][2] = l_cell_wire[1004];							inform_L[1006][2] = l_cell_wire[1005];							inform_L[1003][2] = l_cell_wire[1006];							inform_L[1007][2] = l_cell_wire[1007];							inform_L[1008][2] = l_cell_wire[1008];							inform_L[1012][2] = l_cell_wire[1009];							inform_L[1009][2] = l_cell_wire[1010];							inform_L[1013][2] = l_cell_wire[1011];							inform_L[1010][2] = l_cell_wire[1012];							inform_L[1014][2] = l_cell_wire[1013];							inform_L[1011][2] = l_cell_wire[1014];							inform_L[1015][2] = l_cell_wire[1015];							inform_L[1016][2] = l_cell_wire[1016];							inform_L[1020][2] = l_cell_wire[1017];							inform_L[1017][2] = l_cell_wire[1018];							inform_L[1021][2] = l_cell_wire[1019];							inform_L[1018][2] = l_cell_wire[1020];							inform_L[1022][2] = l_cell_wire[1021];							inform_L[1019][2] = l_cell_wire[1022];							inform_L[1023][2] = l_cell_wire[1023];						end
						4:						begin							inform_R[0][4] = r_cell_wire[0];							inform_R[8][4] = r_cell_wire[1];							inform_R[1][4] = r_cell_wire[2];							inform_R[9][4] = r_cell_wire[3];							inform_R[2][4] = r_cell_wire[4];							inform_R[10][4] = r_cell_wire[5];							inform_R[3][4] = r_cell_wire[6];							inform_R[11][4] = r_cell_wire[7];							inform_R[4][4] = r_cell_wire[8];							inform_R[12][4] = r_cell_wire[9];							inform_R[5][4] = r_cell_wire[10];							inform_R[13][4] = r_cell_wire[11];							inform_R[6][4] = r_cell_wire[12];							inform_R[14][4] = r_cell_wire[13];							inform_R[7][4] = r_cell_wire[14];							inform_R[15][4] = r_cell_wire[15];							inform_R[16][4] = r_cell_wire[16];							inform_R[24][4] = r_cell_wire[17];							inform_R[17][4] = r_cell_wire[18];							inform_R[25][4] = r_cell_wire[19];							inform_R[18][4] = r_cell_wire[20];							inform_R[26][4] = r_cell_wire[21];							inform_R[19][4] = r_cell_wire[22];							inform_R[27][4] = r_cell_wire[23];							inform_R[20][4] = r_cell_wire[24];							inform_R[28][4] = r_cell_wire[25];							inform_R[21][4] = r_cell_wire[26];							inform_R[29][4] = r_cell_wire[27];							inform_R[22][4] = r_cell_wire[28];							inform_R[30][4] = r_cell_wire[29];							inform_R[23][4] = r_cell_wire[30];							inform_R[31][4] = r_cell_wire[31];							inform_R[32][4] = r_cell_wire[32];							inform_R[40][4] = r_cell_wire[33];							inform_R[33][4] = r_cell_wire[34];							inform_R[41][4] = r_cell_wire[35];							inform_R[34][4] = r_cell_wire[36];							inform_R[42][4] = r_cell_wire[37];							inform_R[35][4] = r_cell_wire[38];							inform_R[43][4] = r_cell_wire[39];							inform_R[36][4] = r_cell_wire[40];							inform_R[44][4] = r_cell_wire[41];							inform_R[37][4] = r_cell_wire[42];							inform_R[45][4] = r_cell_wire[43];							inform_R[38][4] = r_cell_wire[44];							inform_R[46][4] = r_cell_wire[45];							inform_R[39][4] = r_cell_wire[46];							inform_R[47][4] = r_cell_wire[47];							inform_R[48][4] = r_cell_wire[48];							inform_R[56][4] = r_cell_wire[49];							inform_R[49][4] = r_cell_wire[50];							inform_R[57][4] = r_cell_wire[51];							inform_R[50][4] = r_cell_wire[52];							inform_R[58][4] = r_cell_wire[53];							inform_R[51][4] = r_cell_wire[54];							inform_R[59][4] = r_cell_wire[55];							inform_R[52][4] = r_cell_wire[56];							inform_R[60][4] = r_cell_wire[57];							inform_R[53][4] = r_cell_wire[58];							inform_R[61][4] = r_cell_wire[59];							inform_R[54][4] = r_cell_wire[60];							inform_R[62][4] = r_cell_wire[61];							inform_R[55][4] = r_cell_wire[62];							inform_R[63][4] = r_cell_wire[63];							inform_R[64][4] = r_cell_wire[64];							inform_R[72][4] = r_cell_wire[65];							inform_R[65][4] = r_cell_wire[66];							inform_R[73][4] = r_cell_wire[67];							inform_R[66][4] = r_cell_wire[68];							inform_R[74][4] = r_cell_wire[69];							inform_R[67][4] = r_cell_wire[70];							inform_R[75][4] = r_cell_wire[71];							inform_R[68][4] = r_cell_wire[72];							inform_R[76][4] = r_cell_wire[73];							inform_R[69][4] = r_cell_wire[74];							inform_R[77][4] = r_cell_wire[75];							inform_R[70][4] = r_cell_wire[76];							inform_R[78][4] = r_cell_wire[77];							inform_R[71][4] = r_cell_wire[78];							inform_R[79][4] = r_cell_wire[79];							inform_R[80][4] = r_cell_wire[80];							inform_R[88][4] = r_cell_wire[81];							inform_R[81][4] = r_cell_wire[82];							inform_R[89][4] = r_cell_wire[83];							inform_R[82][4] = r_cell_wire[84];							inform_R[90][4] = r_cell_wire[85];							inform_R[83][4] = r_cell_wire[86];							inform_R[91][4] = r_cell_wire[87];							inform_R[84][4] = r_cell_wire[88];							inform_R[92][4] = r_cell_wire[89];							inform_R[85][4] = r_cell_wire[90];							inform_R[93][4] = r_cell_wire[91];							inform_R[86][4] = r_cell_wire[92];							inform_R[94][4] = r_cell_wire[93];							inform_R[87][4] = r_cell_wire[94];							inform_R[95][4] = r_cell_wire[95];							inform_R[96][4] = r_cell_wire[96];							inform_R[104][4] = r_cell_wire[97];							inform_R[97][4] = r_cell_wire[98];							inform_R[105][4] = r_cell_wire[99];							inform_R[98][4] = r_cell_wire[100];							inform_R[106][4] = r_cell_wire[101];							inform_R[99][4] = r_cell_wire[102];							inform_R[107][4] = r_cell_wire[103];							inform_R[100][4] = r_cell_wire[104];							inform_R[108][4] = r_cell_wire[105];							inform_R[101][4] = r_cell_wire[106];							inform_R[109][4] = r_cell_wire[107];							inform_R[102][4] = r_cell_wire[108];							inform_R[110][4] = r_cell_wire[109];							inform_R[103][4] = r_cell_wire[110];							inform_R[111][4] = r_cell_wire[111];							inform_R[112][4] = r_cell_wire[112];							inform_R[120][4] = r_cell_wire[113];							inform_R[113][4] = r_cell_wire[114];							inform_R[121][4] = r_cell_wire[115];							inform_R[114][4] = r_cell_wire[116];							inform_R[122][4] = r_cell_wire[117];							inform_R[115][4] = r_cell_wire[118];							inform_R[123][4] = r_cell_wire[119];							inform_R[116][4] = r_cell_wire[120];							inform_R[124][4] = r_cell_wire[121];							inform_R[117][4] = r_cell_wire[122];							inform_R[125][4] = r_cell_wire[123];							inform_R[118][4] = r_cell_wire[124];							inform_R[126][4] = r_cell_wire[125];							inform_R[119][4] = r_cell_wire[126];							inform_R[127][4] = r_cell_wire[127];							inform_R[128][4] = r_cell_wire[128];							inform_R[136][4] = r_cell_wire[129];							inform_R[129][4] = r_cell_wire[130];							inform_R[137][4] = r_cell_wire[131];							inform_R[130][4] = r_cell_wire[132];							inform_R[138][4] = r_cell_wire[133];							inform_R[131][4] = r_cell_wire[134];							inform_R[139][4] = r_cell_wire[135];							inform_R[132][4] = r_cell_wire[136];							inform_R[140][4] = r_cell_wire[137];							inform_R[133][4] = r_cell_wire[138];							inform_R[141][4] = r_cell_wire[139];							inform_R[134][4] = r_cell_wire[140];							inform_R[142][4] = r_cell_wire[141];							inform_R[135][4] = r_cell_wire[142];							inform_R[143][4] = r_cell_wire[143];							inform_R[144][4] = r_cell_wire[144];							inform_R[152][4] = r_cell_wire[145];							inform_R[145][4] = r_cell_wire[146];							inform_R[153][4] = r_cell_wire[147];							inform_R[146][4] = r_cell_wire[148];							inform_R[154][4] = r_cell_wire[149];							inform_R[147][4] = r_cell_wire[150];							inform_R[155][4] = r_cell_wire[151];							inform_R[148][4] = r_cell_wire[152];							inform_R[156][4] = r_cell_wire[153];							inform_R[149][4] = r_cell_wire[154];							inform_R[157][4] = r_cell_wire[155];							inform_R[150][4] = r_cell_wire[156];							inform_R[158][4] = r_cell_wire[157];							inform_R[151][4] = r_cell_wire[158];							inform_R[159][4] = r_cell_wire[159];							inform_R[160][4] = r_cell_wire[160];							inform_R[168][4] = r_cell_wire[161];							inform_R[161][4] = r_cell_wire[162];							inform_R[169][4] = r_cell_wire[163];							inform_R[162][4] = r_cell_wire[164];							inform_R[170][4] = r_cell_wire[165];							inform_R[163][4] = r_cell_wire[166];							inform_R[171][4] = r_cell_wire[167];							inform_R[164][4] = r_cell_wire[168];							inform_R[172][4] = r_cell_wire[169];							inform_R[165][4] = r_cell_wire[170];							inform_R[173][4] = r_cell_wire[171];							inform_R[166][4] = r_cell_wire[172];							inform_R[174][4] = r_cell_wire[173];							inform_R[167][4] = r_cell_wire[174];							inform_R[175][4] = r_cell_wire[175];							inform_R[176][4] = r_cell_wire[176];							inform_R[184][4] = r_cell_wire[177];							inform_R[177][4] = r_cell_wire[178];							inform_R[185][4] = r_cell_wire[179];							inform_R[178][4] = r_cell_wire[180];							inform_R[186][4] = r_cell_wire[181];							inform_R[179][4] = r_cell_wire[182];							inform_R[187][4] = r_cell_wire[183];							inform_R[180][4] = r_cell_wire[184];							inform_R[188][4] = r_cell_wire[185];							inform_R[181][4] = r_cell_wire[186];							inform_R[189][4] = r_cell_wire[187];							inform_R[182][4] = r_cell_wire[188];							inform_R[190][4] = r_cell_wire[189];							inform_R[183][4] = r_cell_wire[190];							inform_R[191][4] = r_cell_wire[191];							inform_R[192][4] = r_cell_wire[192];							inform_R[200][4] = r_cell_wire[193];							inform_R[193][4] = r_cell_wire[194];							inform_R[201][4] = r_cell_wire[195];							inform_R[194][4] = r_cell_wire[196];							inform_R[202][4] = r_cell_wire[197];							inform_R[195][4] = r_cell_wire[198];							inform_R[203][4] = r_cell_wire[199];							inform_R[196][4] = r_cell_wire[200];							inform_R[204][4] = r_cell_wire[201];							inform_R[197][4] = r_cell_wire[202];							inform_R[205][4] = r_cell_wire[203];							inform_R[198][4] = r_cell_wire[204];							inform_R[206][4] = r_cell_wire[205];							inform_R[199][4] = r_cell_wire[206];							inform_R[207][4] = r_cell_wire[207];							inform_R[208][4] = r_cell_wire[208];							inform_R[216][4] = r_cell_wire[209];							inform_R[209][4] = r_cell_wire[210];							inform_R[217][4] = r_cell_wire[211];							inform_R[210][4] = r_cell_wire[212];							inform_R[218][4] = r_cell_wire[213];							inform_R[211][4] = r_cell_wire[214];							inform_R[219][4] = r_cell_wire[215];							inform_R[212][4] = r_cell_wire[216];							inform_R[220][4] = r_cell_wire[217];							inform_R[213][4] = r_cell_wire[218];							inform_R[221][4] = r_cell_wire[219];							inform_R[214][4] = r_cell_wire[220];							inform_R[222][4] = r_cell_wire[221];							inform_R[215][4] = r_cell_wire[222];							inform_R[223][4] = r_cell_wire[223];							inform_R[224][4] = r_cell_wire[224];							inform_R[232][4] = r_cell_wire[225];							inform_R[225][4] = r_cell_wire[226];							inform_R[233][4] = r_cell_wire[227];							inform_R[226][4] = r_cell_wire[228];							inform_R[234][4] = r_cell_wire[229];							inform_R[227][4] = r_cell_wire[230];							inform_R[235][4] = r_cell_wire[231];							inform_R[228][4] = r_cell_wire[232];							inform_R[236][4] = r_cell_wire[233];							inform_R[229][4] = r_cell_wire[234];							inform_R[237][4] = r_cell_wire[235];							inform_R[230][4] = r_cell_wire[236];							inform_R[238][4] = r_cell_wire[237];							inform_R[231][4] = r_cell_wire[238];							inform_R[239][4] = r_cell_wire[239];							inform_R[240][4] = r_cell_wire[240];							inform_R[248][4] = r_cell_wire[241];							inform_R[241][4] = r_cell_wire[242];							inform_R[249][4] = r_cell_wire[243];							inform_R[242][4] = r_cell_wire[244];							inform_R[250][4] = r_cell_wire[245];							inform_R[243][4] = r_cell_wire[246];							inform_R[251][4] = r_cell_wire[247];							inform_R[244][4] = r_cell_wire[248];							inform_R[252][4] = r_cell_wire[249];							inform_R[245][4] = r_cell_wire[250];							inform_R[253][4] = r_cell_wire[251];							inform_R[246][4] = r_cell_wire[252];							inform_R[254][4] = r_cell_wire[253];							inform_R[247][4] = r_cell_wire[254];							inform_R[255][4] = r_cell_wire[255];							inform_R[256][4] = r_cell_wire[256];							inform_R[264][4] = r_cell_wire[257];							inform_R[257][4] = r_cell_wire[258];							inform_R[265][4] = r_cell_wire[259];							inform_R[258][4] = r_cell_wire[260];							inform_R[266][4] = r_cell_wire[261];							inform_R[259][4] = r_cell_wire[262];							inform_R[267][4] = r_cell_wire[263];							inform_R[260][4] = r_cell_wire[264];							inform_R[268][4] = r_cell_wire[265];							inform_R[261][4] = r_cell_wire[266];							inform_R[269][4] = r_cell_wire[267];							inform_R[262][4] = r_cell_wire[268];							inform_R[270][4] = r_cell_wire[269];							inform_R[263][4] = r_cell_wire[270];							inform_R[271][4] = r_cell_wire[271];							inform_R[272][4] = r_cell_wire[272];							inform_R[280][4] = r_cell_wire[273];							inform_R[273][4] = r_cell_wire[274];							inform_R[281][4] = r_cell_wire[275];							inform_R[274][4] = r_cell_wire[276];							inform_R[282][4] = r_cell_wire[277];							inform_R[275][4] = r_cell_wire[278];							inform_R[283][4] = r_cell_wire[279];							inform_R[276][4] = r_cell_wire[280];							inform_R[284][4] = r_cell_wire[281];							inform_R[277][4] = r_cell_wire[282];							inform_R[285][4] = r_cell_wire[283];							inform_R[278][4] = r_cell_wire[284];							inform_R[286][4] = r_cell_wire[285];							inform_R[279][4] = r_cell_wire[286];							inform_R[287][4] = r_cell_wire[287];							inform_R[288][4] = r_cell_wire[288];							inform_R[296][4] = r_cell_wire[289];							inform_R[289][4] = r_cell_wire[290];							inform_R[297][4] = r_cell_wire[291];							inform_R[290][4] = r_cell_wire[292];							inform_R[298][4] = r_cell_wire[293];							inform_R[291][4] = r_cell_wire[294];							inform_R[299][4] = r_cell_wire[295];							inform_R[292][4] = r_cell_wire[296];							inform_R[300][4] = r_cell_wire[297];							inform_R[293][4] = r_cell_wire[298];							inform_R[301][4] = r_cell_wire[299];							inform_R[294][4] = r_cell_wire[300];							inform_R[302][4] = r_cell_wire[301];							inform_R[295][4] = r_cell_wire[302];							inform_R[303][4] = r_cell_wire[303];							inform_R[304][4] = r_cell_wire[304];							inform_R[312][4] = r_cell_wire[305];							inform_R[305][4] = r_cell_wire[306];							inform_R[313][4] = r_cell_wire[307];							inform_R[306][4] = r_cell_wire[308];							inform_R[314][4] = r_cell_wire[309];							inform_R[307][4] = r_cell_wire[310];							inform_R[315][4] = r_cell_wire[311];							inform_R[308][4] = r_cell_wire[312];							inform_R[316][4] = r_cell_wire[313];							inform_R[309][4] = r_cell_wire[314];							inform_R[317][4] = r_cell_wire[315];							inform_R[310][4] = r_cell_wire[316];							inform_R[318][4] = r_cell_wire[317];							inform_R[311][4] = r_cell_wire[318];							inform_R[319][4] = r_cell_wire[319];							inform_R[320][4] = r_cell_wire[320];							inform_R[328][4] = r_cell_wire[321];							inform_R[321][4] = r_cell_wire[322];							inform_R[329][4] = r_cell_wire[323];							inform_R[322][4] = r_cell_wire[324];							inform_R[330][4] = r_cell_wire[325];							inform_R[323][4] = r_cell_wire[326];							inform_R[331][4] = r_cell_wire[327];							inform_R[324][4] = r_cell_wire[328];							inform_R[332][4] = r_cell_wire[329];							inform_R[325][4] = r_cell_wire[330];							inform_R[333][4] = r_cell_wire[331];							inform_R[326][4] = r_cell_wire[332];							inform_R[334][4] = r_cell_wire[333];							inform_R[327][4] = r_cell_wire[334];							inform_R[335][4] = r_cell_wire[335];							inform_R[336][4] = r_cell_wire[336];							inform_R[344][4] = r_cell_wire[337];							inform_R[337][4] = r_cell_wire[338];							inform_R[345][4] = r_cell_wire[339];							inform_R[338][4] = r_cell_wire[340];							inform_R[346][4] = r_cell_wire[341];							inform_R[339][4] = r_cell_wire[342];							inform_R[347][4] = r_cell_wire[343];							inform_R[340][4] = r_cell_wire[344];							inform_R[348][4] = r_cell_wire[345];							inform_R[341][4] = r_cell_wire[346];							inform_R[349][4] = r_cell_wire[347];							inform_R[342][4] = r_cell_wire[348];							inform_R[350][4] = r_cell_wire[349];							inform_R[343][4] = r_cell_wire[350];							inform_R[351][4] = r_cell_wire[351];							inform_R[352][4] = r_cell_wire[352];							inform_R[360][4] = r_cell_wire[353];							inform_R[353][4] = r_cell_wire[354];							inform_R[361][4] = r_cell_wire[355];							inform_R[354][4] = r_cell_wire[356];							inform_R[362][4] = r_cell_wire[357];							inform_R[355][4] = r_cell_wire[358];							inform_R[363][4] = r_cell_wire[359];							inform_R[356][4] = r_cell_wire[360];							inform_R[364][4] = r_cell_wire[361];							inform_R[357][4] = r_cell_wire[362];							inform_R[365][4] = r_cell_wire[363];							inform_R[358][4] = r_cell_wire[364];							inform_R[366][4] = r_cell_wire[365];							inform_R[359][4] = r_cell_wire[366];							inform_R[367][4] = r_cell_wire[367];							inform_R[368][4] = r_cell_wire[368];							inform_R[376][4] = r_cell_wire[369];							inform_R[369][4] = r_cell_wire[370];							inform_R[377][4] = r_cell_wire[371];							inform_R[370][4] = r_cell_wire[372];							inform_R[378][4] = r_cell_wire[373];							inform_R[371][4] = r_cell_wire[374];							inform_R[379][4] = r_cell_wire[375];							inform_R[372][4] = r_cell_wire[376];							inform_R[380][4] = r_cell_wire[377];							inform_R[373][4] = r_cell_wire[378];							inform_R[381][4] = r_cell_wire[379];							inform_R[374][4] = r_cell_wire[380];							inform_R[382][4] = r_cell_wire[381];							inform_R[375][4] = r_cell_wire[382];							inform_R[383][4] = r_cell_wire[383];							inform_R[384][4] = r_cell_wire[384];							inform_R[392][4] = r_cell_wire[385];							inform_R[385][4] = r_cell_wire[386];							inform_R[393][4] = r_cell_wire[387];							inform_R[386][4] = r_cell_wire[388];							inform_R[394][4] = r_cell_wire[389];							inform_R[387][4] = r_cell_wire[390];							inform_R[395][4] = r_cell_wire[391];							inform_R[388][4] = r_cell_wire[392];							inform_R[396][4] = r_cell_wire[393];							inform_R[389][4] = r_cell_wire[394];							inform_R[397][4] = r_cell_wire[395];							inform_R[390][4] = r_cell_wire[396];							inform_R[398][4] = r_cell_wire[397];							inform_R[391][4] = r_cell_wire[398];							inform_R[399][4] = r_cell_wire[399];							inform_R[400][4] = r_cell_wire[400];							inform_R[408][4] = r_cell_wire[401];							inform_R[401][4] = r_cell_wire[402];							inform_R[409][4] = r_cell_wire[403];							inform_R[402][4] = r_cell_wire[404];							inform_R[410][4] = r_cell_wire[405];							inform_R[403][4] = r_cell_wire[406];							inform_R[411][4] = r_cell_wire[407];							inform_R[404][4] = r_cell_wire[408];							inform_R[412][4] = r_cell_wire[409];							inform_R[405][4] = r_cell_wire[410];							inform_R[413][4] = r_cell_wire[411];							inform_R[406][4] = r_cell_wire[412];							inform_R[414][4] = r_cell_wire[413];							inform_R[407][4] = r_cell_wire[414];							inform_R[415][4] = r_cell_wire[415];							inform_R[416][4] = r_cell_wire[416];							inform_R[424][4] = r_cell_wire[417];							inform_R[417][4] = r_cell_wire[418];							inform_R[425][4] = r_cell_wire[419];							inform_R[418][4] = r_cell_wire[420];							inform_R[426][4] = r_cell_wire[421];							inform_R[419][4] = r_cell_wire[422];							inform_R[427][4] = r_cell_wire[423];							inform_R[420][4] = r_cell_wire[424];							inform_R[428][4] = r_cell_wire[425];							inform_R[421][4] = r_cell_wire[426];							inform_R[429][4] = r_cell_wire[427];							inform_R[422][4] = r_cell_wire[428];							inform_R[430][4] = r_cell_wire[429];							inform_R[423][4] = r_cell_wire[430];							inform_R[431][4] = r_cell_wire[431];							inform_R[432][4] = r_cell_wire[432];							inform_R[440][4] = r_cell_wire[433];							inform_R[433][4] = r_cell_wire[434];							inform_R[441][4] = r_cell_wire[435];							inform_R[434][4] = r_cell_wire[436];							inform_R[442][4] = r_cell_wire[437];							inform_R[435][4] = r_cell_wire[438];							inform_R[443][4] = r_cell_wire[439];							inform_R[436][4] = r_cell_wire[440];							inform_R[444][4] = r_cell_wire[441];							inform_R[437][4] = r_cell_wire[442];							inform_R[445][4] = r_cell_wire[443];							inform_R[438][4] = r_cell_wire[444];							inform_R[446][4] = r_cell_wire[445];							inform_R[439][4] = r_cell_wire[446];							inform_R[447][4] = r_cell_wire[447];							inform_R[448][4] = r_cell_wire[448];							inform_R[456][4] = r_cell_wire[449];							inform_R[449][4] = r_cell_wire[450];							inform_R[457][4] = r_cell_wire[451];							inform_R[450][4] = r_cell_wire[452];							inform_R[458][4] = r_cell_wire[453];							inform_R[451][4] = r_cell_wire[454];							inform_R[459][4] = r_cell_wire[455];							inform_R[452][4] = r_cell_wire[456];							inform_R[460][4] = r_cell_wire[457];							inform_R[453][4] = r_cell_wire[458];							inform_R[461][4] = r_cell_wire[459];							inform_R[454][4] = r_cell_wire[460];							inform_R[462][4] = r_cell_wire[461];							inform_R[455][4] = r_cell_wire[462];							inform_R[463][4] = r_cell_wire[463];							inform_R[464][4] = r_cell_wire[464];							inform_R[472][4] = r_cell_wire[465];							inform_R[465][4] = r_cell_wire[466];							inform_R[473][4] = r_cell_wire[467];							inform_R[466][4] = r_cell_wire[468];							inform_R[474][4] = r_cell_wire[469];							inform_R[467][4] = r_cell_wire[470];							inform_R[475][4] = r_cell_wire[471];							inform_R[468][4] = r_cell_wire[472];							inform_R[476][4] = r_cell_wire[473];							inform_R[469][4] = r_cell_wire[474];							inform_R[477][4] = r_cell_wire[475];							inform_R[470][4] = r_cell_wire[476];							inform_R[478][4] = r_cell_wire[477];							inform_R[471][4] = r_cell_wire[478];							inform_R[479][4] = r_cell_wire[479];							inform_R[480][4] = r_cell_wire[480];							inform_R[488][4] = r_cell_wire[481];							inform_R[481][4] = r_cell_wire[482];							inform_R[489][4] = r_cell_wire[483];							inform_R[482][4] = r_cell_wire[484];							inform_R[490][4] = r_cell_wire[485];							inform_R[483][4] = r_cell_wire[486];							inform_R[491][4] = r_cell_wire[487];							inform_R[484][4] = r_cell_wire[488];							inform_R[492][4] = r_cell_wire[489];							inform_R[485][4] = r_cell_wire[490];							inform_R[493][4] = r_cell_wire[491];							inform_R[486][4] = r_cell_wire[492];							inform_R[494][4] = r_cell_wire[493];							inform_R[487][4] = r_cell_wire[494];							inform_R[495][4] = r_cell_wire[495];							inform_R[496][4] = r_cell_wire[496];							inform_R[504][4] = r_cell_wire[497];							inform_R[497][4] = r_cell_wire[498];							inform_R[505][4] = r_cell_wire[499];							inform_R[498][4] = r_cell_wire[500];							inform_R[506][4] = r_cell_wire[501];							inform_R[499][4] = r_cell_wire[502];							inform_R[507][4] = r_cell_wire[503];							inform_R[500][4] = r_cell_wire[504];							inform_R[508][4] = r_cell_wire[505];							inform_R[501][4] = r_cell_wire[506];							inform_R[509][4] = r_cell_wire[507];							inform_R[502][4] = r_cell_wire[508];							inform_R[510][4] = r_cell_wire[509];							inform_R[503][4] = r_cell_wire[510];							inform_R[511][4] = r_cell_wire[511];							inform_R[512][4] = r_cell_wire[512];							inform_R[520][4] = r_cell_wire[513];							inform_R[513][4] = r_cell_wire[514];							inform_R[521][4] = r_cell_wire[515];							inform_R[514][4] = r_cell_wire[516];							inform_R[522][4] = r_cell_wire[517];							inform_R[515][4] = r_cell_wire[518];							inform_R[523][4] = r_cell_wire[519];							inform_R[516][4] = r_cell_wire[520];							inform_R[524][4] = r_cell_wire[521];							inform_R[517][4] = r_cell_wire[522];							inform_R[525][4] = r_cell_wire[523];							inform_R[518][4] = r_cell_wire[524];							inform_R[526][4] = r_cell_wire[525];							inform_R[519][4] = r_cell_wire[526];							inform_R[527][4] = r_cell_wire[527];							inform_R[528][4] = r_cell_wire[528];							inform_R[536][4] = r_cell_wire[529];							inform_R[529][4] = r_cell_wire[530];							inform_R[537][4] = r_cell_wire[531];							inform_R[530][4] = r_cell_wire[532];							inform_R[538][4] = r_cell_wire[533];							inform_R[531][4] = r_cell_wire[534];							inform_R[539][4] = r_cell_wire[535];							inform_R[532][4] = r_cell_wire[536];							inform_R[540][4] = r_cell_wire[537];							inform_R[533][4] = r_cell_wire[538];							inform_R[541][4] = r_cell_wire[539];							inform_R[534][4] = r_cell_wire[540];							inform_R[542][4] = r_cell_wire[541];							inform_R[535][4] = r_cell_wire[542];							inform_R[543][4] = r_cell_wire[543];							inform_R[544][4] = r_cell_wire[544];							inform_R[552][4] = r_cell_wire[545];							inform_R[545][4] = r_cell_wire[546];							inform_R[553][4] = r_cell_wire[547];							inform_R[546][4] = r_cell_wire[548];							inform_R[554][4] = r_cell_wire[549];							inform_R[547][4] = r_cell_wire[550];							inform_R[555][4] = r_cell_wire[551];							inform_R[548][4] = r_cell_wire[552];							inform_R[556][4] = r_cell_wire[553];							inform_R[549][4] = r_cell_wire[554];							inform_R[557][4] = r_cell_wire[555];							inform_R[550][4] = r_cell_wire[556];							inform_R[558][4] = r_cell_wire[557];							inform_R[551][4] = r_cell_wire[558];							inform_R[559][4] = r_cell_wire[559];							inform_R[560][4] = r_cell_wire[560];							inform_R[568][4] = r_cell_wire[561];							inform_R[561][4] = r_cell_wire[562];							inform_R[569][4] = r_cell_wire[563];							inform_R[562][4] = r_cell_wire[564];							inform_R[570][4] = r_cell_wire[565];							inform_R[563][4] = r_cell_wire[566];							inform_R[571][4] = r_cell_wire[567];							inform_R[564][4] = r_cell_wire[568];							inform_R[572][4] = r_cell_wire[569];							inform_R[565][4] = r_cell_wire[570];							inform_R[573][4] = r_cell_wire[571];							inform_R[566][4] = r_cell_wire[572];							inform_R[574][4] = r_cell_wire[573];							inform_R[567][4] = r_cell_wire[574];							inform_R[575][4] = r_cell_wire[575];							inform_R[576][4] = r_cell_wire[576];							inform_R[584][4] = r_cell_wire[577];							inform_R[577][4] = r_cell_wire[578];							inform_R[585][4] = r_cell_wire[579];							inform_R[578][4] = r_cell_wire[580];							inform_R[586][4] = r_cell_wire[581];							inform_R[579][4] = r_cell_wire[582];							inform_R[587][4] = r_cell_wire[583];							inform_R[580][4] = r_cell_wire[584];							inform_R[588][4] = r_cell_wire[585];							inform_R[581][4] = r_cell_wire[586];							inform_R[589][4] = r_cell_wire[587];							inform_R[582][4] = r_cell_wire[588];							inform_R[590][4] = r_cell_wire[589];							inform_R[583][4] = r_cell_wire[590];							inform_R[591][4] = r_cell_wire[591];							inform_R[592][4] = r_cell_wire[592];							inform_R[600][4] = r_cell_wire[593];							inform_R[593][4] = r_cell_wire[594];							inform_R[601][4] = r_cell_wire[595];							inform_R[594][4] = r_cell_wire[596];							inform_R[602][4] = r_cell_wire[597];							inform_R[595][4] = r_cell_wire[598];							inform_R[603][4] = r_cell_wire[599];							inform_R[596][4] = r_cell_wire[600];							inform_R[604][4] = r_cell_wire[601];							inform_R[597][4] = r_cell_wire[602];							inform_R[605][4] = r_cell_wire[603];							inform_R[598][4] = r_cell_wire[604];							inform_R[606][4] = r_cell_wire[605];							inform_R[599][4] = r_cell_wire[606];							inform_R[607][4] = r_cell_wire[607];							inform_R[608][4] = r_cell_wire[608];							inform_R[616][4] = r_cell_wire[609];							inform_R[609][4] = r_cell_wire[610];							inform_R[617][4] = r_cell_wire[611];							inform_R[610][4] = r_cell_wire[612];							inform_R[618][4] = r_cell_wire[613];							inform_R[611][4] = r_cell_wire[614];							inform_R[619][4] = r_cell_wire[615];							inform_R[612][4] = r_cell_wire[616];							inform_R[620][4] = r_cell_wire[617];							inform_R[613][4] = r_cell_wire[618];							inform_R[621][4] = r_cell_wire[619];							inform_R[614][4] = r_cell_wire[620];							inform_R[622][4] = r_cell_wire[621];							inform_R[615][4] = r_cell_wire[622];							inform_R[623][4] = r_cell_wire[623];							inform_R[624][4] = r_cell_wire[624];							inform_R[632][4] = r_cell_wire[625];							inform_R[625][4] = r_cell_wire[626];							inform_R[633][4] = r_cell_wire[627];							inform_R[626][4] = r_cell_wire[628];							inform_R[634][4] = r_cell_wire[629];							inform_R[627][4] = r_cell_wire[630];							inform_R[635][4] = r_cell_wire[631];							inform_R[628][4] = r_cell_wire[632];							inform_R[636][4] = r_cell_wire[633];							inform_R[629][4] = r_cell_wire[634];							inform_R[637][4] = r_cell_wire[635];							inform_R[630][4] = r_cell_wire[636];							inform_R[638][4] = r_cell_wire[637];							inform_R[631][4] = r_cell_wire[638];							inform_R[639][4] = r_cell_wire[639];							inform_R[640][4] = r_cell_wire[640];							inform_R[648][4] = r_cell_wire[641];							inform_R[641][4] = r_cell_wire[642];							inform_R[649][4] = r_cell_wire[643];							inform_R[642][4] = r_cell_wire[644];							inform_R[650][4] = r_cell_wire[645];							inform_R[643][4] = r_cell_wire[646];							inform_R[651][4] = r_cell_wire[647];							inform_R[644][4] = r_cell_wire[648];							inform_R[652][4] = r_cell_wire[649];							inform_R[645][4] = r_cell_wire[650];							inform_R[653][4] = r_cell_wire[651];							inform_R[646][4] = r_cell_wire[652];							inform_R[654][4] = r_cell_wire[653];							inform_R[647][4] = r_cell_wire[654];							inform_R[655][4] = r_cell_wire[655];							inform_R[656][4] = r_cell_wire[656];							inform_R[664][4] = r_cell_wire[657];							inform_R[657][4] = r_cell_wire[658];							inform_R[665][4] = r_cell_wire[659];							inform_R[658][4] = r_cell_wire[660];							inform_R[666][4] = r_cell_wire[661];							inform_R[659][4] = r_cell_wire[662];							inform_R[667][4] = r_cell_wire[663];							inform_R[660][4] = r_cell_wire[664];							inform_R[668][4] = r_cell_wire[665];							inform_R[661][4] = r_cell_wire[666];							inform_R[669][4] = r_cell_wire[667];							inform_R[662][4] = r_cell_wire[668];							inform_R[670][4] = r_cell_wire[669];							inform_R[663][4] = r_cell_wire[670];							inform_R[671][4] = r_cell_wire[671];							inform_R[672][4] = r_cell_wire[672];							inform_R[680][4] = r_cell_wire[673];							inform_R[673][4] = r_cell_wire[674];							inform_R[681][4] = r_cell_wire[675];							inform_R[674][4] = r_cell_wire[676];							inform_R[682][4] = r_cell_wire[677];							inform_R[675][4] = r_cell_wire[678];							inform_R[683][4] = r_cell_wire[679];							inform_R[676][4] = r_cell_wire[680];							inform_R[684][4] = r_cell_wire[681];							inform_R[677][4] = r_cell_wire[682];							inform_R[685][4] = r_cell_wire[683];							inform_R[678][4] = r_cell_wire[684];							inform_R[686][4] = r_cell_wire[685];							inform_R[679][4] = r_cell_wire[686];							inform_R[687][4] = r_cell_wire[687];							inform_R[688][4] = r_cell_wire[688];							inform_R[696][4] = r_cell_wire[689];							inform_R[689][4] = r_cell_wire[690];							inform_R[697][4] = r_cell_wire[691];							inform_R[690][4] = r_cell_wire[692];							inform_R[698][4] = r_cell_wire[693];							inform_R[691][4] = r_cell_wire[694];							inform_R[699][4] = r_cell_wire[695];							inform_R[692][4] = r_cell_wire[696];							inform_R[700][4] = r_cell_wire[697];							inform_R[693][4] = r_cell_wire[698];							inform_R[701][4] = r_cell_wire[699];							inform_R[694][4] = r_cell_wire[700];							inform_R[702][4] = r_cell_wire[701];							inform_R[695][4] = r_cell_wire[702];							inform_R[703][4] = r_cell_wire[703];							inform_R[704][4] = r_cell_wire[704];							inform_R[712][4] = r_cell_wire[705];							inform_R[705][4] = r_cell_wire[706];							inform_R[713][4] = r_cell_wire[707];							inform_R[706][4] = r_cell_wire[708];							inform_R[714][4] = r_cell_wire[709];							inform_R[707][4] = r_cell_wire[710];							inform_R[715][4] = r_cell_wire[711];							inform_R[708][4] = r_cell_wire[712];							inform_R[716][4] = r_cell_wire[713];							inform_R[709][4] = r_cell_wire[714];							inform_R[717][4] = r_cell_wire[715];							inform_R[710][4] = r_cell_wire[716];							inform_R[718][4] = r_cell_wire[717];							inform_R[711][4] = r_cell_wire[718];							inform_R[719][4] = r_cell_wire[719];							inform_R[720][4] = r_cell_wire[720];							inform_R[728][4] = r_cell_wire[721];							inform_R[721][4] = r_cell_wire[722];							inform_R[729][4] = r_cell_wire[723];							inform_R[722][4] = r_cell_wire[724];							inform_R[730][4] = r_cell_wire[725];							inform_R[723][4] = r_cell_wire[726];							inform_R[731][4] = r_cell_wire[727];							inform_R[724][4] = r_cell_wire[728];							inform_R[732][4] = r_cell_wire[729];							inform_R[725][4] = r_cell_wire[730];							inform_R[733][4] = r_cell_wire[731];							inform_R[726][4] = r_cell_wire[732];							inform_R[734][4] = r_cell_wire[733];							inform_R[727][4] = r_cell_wire[734];							inform_R[735][4] = r_cell_wire[735];							inform_R[736][4] = r_cell_wire[736];							inform_R[744][4] = r_cell_wire[737];							inform_R[737][4] = r_cell_wire[738];							inform_R[745][4] = r_cell_wire[739];							inform_R[738][4] = r_cell_wire[740];							inform_R[746][4] = r_cell_wire[741];							inform_R[739][4] = r_cell_wire[742];							inform_R[747][4] = r_cell_wire[743];							inform_R[740][4] = r_cell_wire[744];							inform_R[748][4] = r_cell_wire[745];							inform_R[741][4] = r_cell_wire[746];							inform_R[749][4] = r_cell_wire[747];							inform_R[742][4] = r_cell_wire[748];							inform_R[750][4] = r_cell_wire[749];							inform_R[743][4] = r_cell_wire[750];							inform_R[751][4] = r_cell_wire[751];							inform_R[752][4] = r_cell_wire[752];							inform_R[760][4] = r_cell_wire[753];							inform_R[753][4] = r_cell_wire[754];							inform_R[761][4] = r_cell_wire[755];							inform_R[754][4] = r_cell_wire[756];							inform_R[762][4] = r_cell_wire[757];							inform_R[755][4] = r_cell_wire[758];							inform_R[763][4] = r_cell_wire[759];							inform_R[756][4] = r_cell_wire[760];							inform_R[764][4] = r_cell_wire[761];							inform_R[757][4] = r_cell_wire[762];							inform_R[765][4] = r_cell_wire[763];							inform_R[758][4] = r_cell_wire[764];							inform_R[766][4] = r_cell_wire[765];							inform_R[759][4] = r_cell_wire[766];							inform_R[767][4] = r_cell_wire[767];							inform_R[768][4] = r_cell_wire[768];							inform_R[776][4] = r_cell_wire[769];							inform_R[769][4] = r_cell_wire[770];							inform_R[777][4] = r_cell_wire[771];							inform_R[770][4] = r_cell_wire[772];							inform_R[778][4] = r_cell_wire[773];							inform_R[771][4] = r_cell_wire[774];							inform_R[779][4] = r_cell_wire[775];							inform_R[772][4] = r_cell_wire[776];							inform_R[780][4] = r_cell_wire[777];							inform_R[773][4] = r_cell_wire[778];							inform_R[781][4] = r_cell_wire[779];							inform_R[774][4] = r_cell_wire[780];							inform_R[782][4] = r_cell_wire[781];							inform_R[775][4] = r_cell_wire[782];							inform_R[783][4] = r_cell_wire[783];							inform_R[784][4] = r_cell_wire[784];							inform_R[792][4] = r_cell_wire[785];							inform_R[785][4] = r_cell_wire[786];							inform_R[793][4] = r_cell_wire[787];							inform_R[786][4] = r_cell_wire[788];							inform_R[794][4] = r_cell_wire[789];							inform_R[787][4] = r_cell_wire[790];							inform_R[795][4] = r_cell_wire[791];							inform_R[788][4] = r_cell_wire[792];							inform_R[796][4] = r_cell_wire[793];							inform_R[789][4] = r_cell_wire[794];							inform_R[797][4] = r_cell_wire[795];							inform_R[790][4] = r_cell_wire[796];							inform_R[798][4] = r_cell_wire[797];							inform_R[791][4] = r_cell_wire[798];							inform_R[799][4] = r_cell_wire[799];							inform_R[800][4] = r_cell_wire[800];							inform_R[808][4] = r_cell_wire[801];							inform_R[801][4] = r_cell_wire[802];							inform_R[809][4] = r_cell_wire[803];							inform_R[802][4] = r_cell_wire[804];							inform_R[810][4] = r_cell_wire[805];							inform_R[803][4] = r_cell_wire[806];							inform_R[811][4] = r_cell_wire[807];							inform_R[804][4] = r_cell_wire[808];							inform_R[812][4] = r_cell_wire[809];							inform_R[805][4] = r_cell_wire[810];							inform_R[813][4] = r_cell_wire[811];							inform_R[806][4] = r_cell_wire[812];							inform_R[814][4] = r_cell_wire[813];							inform_R[807][4] = r_cell_wire[814];							inform_R[815][4] = r_cell_wire[815];							inform_R[816][4] = r_cell_wire[816];							inform_R[824][4] = r_cell_wire[817];							inform_R[817][4] = r_cell_wire[818];							inform_R[825][4] = r_cell_wire[819];							inform_R[818][4] = r_cell_wire[820];							inform_R[826][4] = r_cell_wire[821];							inform_R[819][4] = r_cell_wire[822];							inform_R[827][4] = r_cell_wire[823];							inform_R[820][4] = r_cell_wire[824];							inform_R[828][4] = r_cell_wire[825];							inform_R[821][4] = r_cell_wire[826];							inform_R[829][4] = r_cell_wire[827];							inform_R[822][4] = r_cell_wire[828];							inform_R[830][4] = r_cell_wire[829];							inform_R[823][4] = r_cell_wire[830];							inform_R[831][4] = r_cell_wire[831];							inform_R[832][4] = r_cell_wire[832];							inform_R[840][4] = r_cell_wire[833];							inform_R[833][4] = r_cell_wire[834];							inform_R[841][4] = r_cell_wire[835];							inform_R[834][4] = r_cell_wire[836];							inform_R[842][4] = r_cell_wire[837];							inform_R[835][4] = r_cell_wire[838];							inform_R[843][4] = r_cell_wire[839];							inform_R[836][4] = r_cell_wire[840];							inform_R[844][4] = r_cell_wire[841];							inform_R[837][4] = r_cell_wire[842];							inform_R[845][4] = r_cell_wire[843];							inform_R[838][4] = r_cell_wire[844];							inform_R[846][4] = r_cell_wire[845];							inform_R[839][4] = r_cell_wire[846];							inform_R[847][4] = r_cell_wire[847];							inform_R[848][4] = r_cell_wire[848];							inform_R[856][4] = r_cell_wire[849];							inform_R[849][4] = r_cell_wire[850];							inform_R[857][4] = r_cell_wire[851];							inform_R[850][4] = r_cell_wire[852];							inform_R[858][4] = r_cell_wire[853];							inform_R[851][4] = r_cell_wire[854];							inform_R[859][4] = r_cell_wire[855];							inform_R[852][4] = r_cell_wire[856];							inform_R[860][4] = r_cell_wire[857];							inform_R[853][4] = r_cell_wire[858];							inform_R[861][4] = r_cell_wire[859];							inform_R[854][4] = r_cell_wire[860];							inform_R[862][4] = r_cell_wire[861];							inform_R[855][4] = r_cell_wire[862];							inform_R[863][4] = r_cell_wire[863];							inform_R[864][4] = r_cell_wire[864];							inform_R[872][4] = r_cell_wire[865];							inform_R[865][4] = r_cell_wire[866];							inform_R[873][4] = r_cell_wire[867];							inform_R[866][4] = r_cell_wire[868];							inform_R[874][4] = r_cell_wire[869];							inform_R[867][4] = r_cell_wire[870];							inform_R[875][4] = r_cell_wire[871];							inform_R[868][4] = r_cell_wire[872];							inform_R[876][4] = r_cell_wire[873];							inform_R[869][4] = r_cell_wire[874];							inform_R[877][4] = r_cell_wire[875];							inform_R[870][4] = r_cell_wire[876];							inform_R[878][4] = r_cell_wire[877];							inform_R[871][4] = r_cell_wire[878];							inform_R[879][4] = r_cell_wire[879];							inform_R[880][4] = r_cell_wire[880];							inform_R[888][4] = r_cell_wire[881];							inform_R[881][4] = r_cell_wire[882];							inform_R[889][4] = r_cell_wire[883];							inform_R[882][4] = r_cell_wire[884];							inform_R[890][4] = r_cell_wire[885];							inform_R[883][4] = r_cell_wire[886];							inform_R[891][4] = r_cell_wire[887];							inform_R[884][4] = r_cell_wire[888];							inform_R[892][4] = r_cell_wire[889];							inform_R[885][4] = r_cell_wire[890];							inform_R[893][4] = r_cell_wire[891];							inform_R[886][4] = r_cell_wire[892];							inform_R[894][4] = r_cell_wire[893];							inform_R[887][4] = r_cell_wire[894];							inform_R[895][4] = r_cell_wire[895];							inform_R[896][4] = r_cell_wire[896];							inform_R[904][4] = r_cell_wire[897];							inform_R[897][4] = r_cell_wire[898];							inform_R[905][4] = r_cell_wire[899];							inform_R[898][4] = r_cell_wire[900];							inform_R[906][4] = r_cell_wire[901];							inform_R[899][4] = r_cell_wire[902];							inform_R[907][4] = r_cell_wire[903];							inform_R[900][4] = r_cell_wire[904];							inform_R[908][4] = r_cell_wire[905];							inform_R[901][4] = r_cell_wire[906];							inform_R[909][4] = r_cell_wire[907];							inform_R[902][4] = r_cell_wire[908];							inform_R[910][4] = r_cell_wire[909];							inform_R[903][4] = r_cell_wire[910];							inform_R[911][4] = r_cell_wire[911];							inform_R[912][4] = r_cell_wire[912];							inform_R[920][4] = r_cell_wire[913];							inform_R[913][4] = r_cell_wire[914];							inform_R[921][4] = r_cell_wire[915];							inform_R[914][4] = r_cell_wire[916];							inform_R[922][4] = r_cell_wire[917];							inform_R[915][4] = r_cell_wire[918];							inform_R[923][4] = r_cell_wire[919];							inform_R[916][4] = r_cell_wire[920];							inform_R[924][4] = r_cell_wire[921];							inform_R[917][4] = r_cell_wire[922];							inform_R[925][4] = r_cell_wire[923];							inform_R[918][4] = r_cell_wire[924];							inform_R[926][4] = r_cell_wire[925];							inform_R[919][4] = r_cell_wire[926];							inform_R[927][4] = r_cell_wire[927];							inform_R[928][4] = r_cell_wire[928];							inform_R[936][4] = r_cell_wire[929];							inform_R[929][4] = r_cell_wire[930];							inform_R[937][4] = r_cell_wire[931];							inform_R[930][4] = r_cell_wire[932];							inform_R[938][4] = r_cell_wire[933];							inform_R[931][4] = r_cell_wire[934];							inform_R[939][4] = r_cell_wire[935];							inform_R[932][4] = r_cell_wire[936];							inform_R[940][4] = r_cell_wire[937];							inform_R[933][4] = r_cell_wire[938];							inform_R[941][4] = r_cell_wire[939];							inform_R[934][4] = r_cell_wire[940];							inform_R[942][4] = r_cell_wire[941];							inform_R[935][4] = r_cell_wire[942];							inform_R[943][4] = r_cell_wire[943];							inform_R[944][4] = r_cell_wire[944];							inform_R[952][4] = r_cell_wire[945];							inform_R[945][4] = r_cell_wire[946];							inform_R[953][4] = r_cell_wire[947];							inform_R[946][4] = r_cell_wire[948];							inform_R[954][4] = r_cell_wire[949];							inform_R[947][4] = r_cell_wire[950];							inform_R[955][4] = r_cell_wire[951];							inform_R[948][4] = r_cell_wire[952];							inform_R[956][4] = r_cell_wire[953];							inform_R[949][4] = r_cell_wire[954];							inform_R[957][4] = r_cell_wire[955];							inform_R[950][4] = r_cell_wire[956];							inform_R[958][4] = r_cell_wire[957];							inform_R[951][4] = r_cell_wire[958];							inform_R[959][4] = r_cell_wire[959];							inform_R[960][4] = r_cell_wire[960];							inform_R[968][4] = r_cell_wire[961];							inform_R[961][4] = r_cell_wire[962];							inform_R[969][4] = r_cell_wire[963];							inform_R[962][4] = r_cell_wire[964];							inform_R[970][4] = r_cell_wire[965];							inform_R[963][4] = r_cell_wire[966];							inform_R[971][4] = r_cell_wire[967];							inform_R[964][4] = r_cell_wire[968];							inform_R[972][4] = r_cell_wire[969];							inform_R[965][4] = r_cell_wire[970];							inform_R[973][4] = r_cell_wire[971];							inform_R[966][4] = r_cell_wire[972];							inform_R[974][4] = r_cell_wire[973];							inform_R[967][4] = r_cell_wire[974];							inform_R[975][4] = r_cell_wire[975];							inform_R[976][4] = r_cell_wire[976];							inform_R[984][4] = r_cell_wire[977];							inform_R[977][4] = r_cell_wire[978];							inform_R[985][4] = r_cell_wire[979];							inform_R[978][4] = r_cell_wire[980];							inform_R[986][4] = r_cell_wire[981];							inform_R[979][4] = r_cell_wire[982];							inform_R[987][4] = r_cell_wire[983];							inform_R[980][4] = r_cell_wire[984];							inform_R[988][4] = r_cell_wire[985];							inform_R[981][4] = r_cell_wire[986];							inform_R[989][4] = r_cell_wire[987];							inform_R[982][4] = r_cell_wire[988];							inform_R[990][4] = r_cell_wire[989];							inform_R[983][4] = r_cell_wire[990];							inform_R[991][4] = r_cell_wire[991];							inform_R[992][4] = r_cell_wire[992];							inform_R[1000][4] = r_cell_wire[993];							inform_R[993][4] = r_cell_wire[994];							inform_R[1001][4] = r_cell_wire[995];							inform_R[994][4] = r_cell_wire[996];							inform_R[1002][4] = r_cell_wire[997];							inform_R[995][4] = r_cell_wire[998];							inform_R[1003][4] = r_cell_wire[999];							inform_R[996][4] = r_cell_wire[1000];							inform_R[1004][4] = r_cell_wire[1001];							inform_R[997][4] = r_cell_wire[1002];							inform_R[1005][4] = r_cell_wire[1003];							inform_R[998][4] = r_cell_wire[1004];							inform_R[1006][4] = r_cell_wire[1005];							inform_R[999][4] = r_cell_wire[1006];							inform_R[1007][4] = r_cell_wire[1007];							inform_R[1008][4] = r_cell_wire[1008];							inform_R[1016][4] = r_cell_wire[1009];							inform_R[1009][4] = r_cell_wire[1010];							inform_R[1017][4] = r_cell_wire[1011];							inform_R[1010][4] = r_cell_wire[1012];							inform_R[1018][4] = r_cell_wire[1013];							inform_R[1011][4] = r_cell_wire[1014];							inform_R[1019][4] = r_cell_wire[1015];							inform_R[1012][4] = r_cell_wire[1016];							inform_R[1020][4] = r_cell_wire[1017];							inform_R[1013][4] = r_cell_wire[1018];							inform_R[1021][4] = r_cell_wire[1019];							inform_R[1014][4] = r_cell_wire[1020];							inform_R[1022][4] = r_cell_wire[1021];							inform_R[1015][4] = r_cell_wire[1022];							inform_R[1023][4] = r_cell_wire[1023];							inform_L[0][3] = l_cell_wire[0];							inform_L[8][3] = l_cell_wire[1];							inform_L[1][3] = l_cell_wire[2];							inform_L[9][3] = l_cell_wire[3];							inform_L[2][3] = l_cell_wire[4];							inform_L[10][3] = l_cell_wire[5];							inform_L[3][3] = l_cell_wire[6];							inform_L[11][3] = l_cell_wire[7];							inform_L[4][3] = l_cell_wire[8];							inform_L[12][3] = l_cell_wire[9];							inform_L[5][3] = l_cell_wire[10];							inform_L[13][3] = l_cell_wire[11];							inform_L[6][3] = l_cell_wire[12];							inform_L[14][3] = l_cell_wire[13];							inform_L[7][3] = l_cell_wire[14];							inform_L[15][3] = l_cell_wire[15];							inform_L[16][3] = l_cell_wire[16];							inform_L[24][3] = l_cell_wire[17];							inform_L[17][3] = l_cell_wire[18];							inform_L[25][3] = l_cell_wire[19];							inform_L[18][3] = l_cell_wire[20];							inform_L[26][3] = l_cell_wire[21];							inform_L[19][3] = l_cell_wire[22];							inform_L[27][3] = l_cell_wire[23];							inform_L[20][3] = l_cell_wire[24];							inform_L[28][3] = l_cell_wire[25];							inform_L[21][3] = l_cell_wire[26];							inform_L[29][3] = l_cell_wire[27];							inform_L[22][3] = l_cell_wire[28];							inform_L[30][3] = l_cell_wire[29];							inform_L[23][3] = l_cell_wire[30];							inform_L[31][3] = l_cell_wire[31];							inform_L[32][3] = l_cell_wire[32];							inform_L[40][3] = l_cell_wire[33];							inform_L[33][3] = l_cell_wire[34];							inform_L[41][3] = l_cell_wire[35];							inform_L[34][3] = l_cell_wire[36];							inform_L[42][3] = l_cell_wire[37];							inform_L[35][3] = l_cell_wire[38];							inform_L[43][3] = l_cell_wire[39];							inform_L[36][3] = l_cell_wire[40];							inform_L[44][3] = l_cell_wire[41];							inform_L[37][3] = l_cell_wire[42];							inform_L[45][3] = l_cell_wire[43];							inform_L[38][3] = l_cell_wire[44];							inform_L[46][3] = l_cell_wire[45];							inform_L[39][3] = l_cell_wire[46];							inform_L[47][3] = l_cell_wire[47];							inform_L[48][3] = l_cell_wire[48];							inform_L[56][3] = l_cell_wire[49];							inform_L[49][3] = l_cell_wire[50];							inform_L[57][3] = l_cell_wire[51];							inform_L[50][3] = l_cell_wire[52];							inform_L[58][3] = l_cell_wire[53];							inform_L[51][3] = l_cell_wire[54];							inform_L[59][3] = l_cell_wire[55];							inform_L[52][3] = l_cell_wire[56];							inform_L[60][3] = l_cell_wire[57];							inform_L[53][3] = l_cell_wire[58];							inform_L[61][3] = l_cell_wire[59];							inform_L[54][3] = l_cell_wire[60];							inform_L[62][3] = l_cell_wire[61];							inform_L[55][3] = l_cell_wire[62];							inform_L[63][3] = l_cell_wire[63];							inform_L[64][3] = l_cell_wire[64];							inform_L[72][3] = l_cell_wire[65];							inform_L[65][3] = l_cell_wire[66];							inform_L[73][3] = l_cell_wire[67];							inform_L[66][3] = l_cell_wire[68];							inform_L[74][3] = l_cell_wire[69];							inform_L[67][3] = l_cell_wire[70];							inform_L[75][3] = l_cell_wire[71];							inform_L[68][3] = l_cell_wire[72];							inform_L[76][3] = l_cell_wire[73];							inform_L[69][3] = l_cell_wire[74];							inform_L[77][3] = l_cell_wire[75];							inform_L[70][3] = l_cell_wire[76];							inform_L[78][3] = l_cell_wire[77];							inform_L[71][3] = l_cell_wire[78];							inform_L[79][3] = l_cell_wire[79];							inform_L[80][3] = l_cell_wire[80];							inform_L[88][3] = l_cell_wire[81];							inform_L[81][3] = l_cell_wire[82];							inform_L[89][3] = l_cell_wire[83];							inform_L[82][3] = l_cell_wire[84];							inform_L[90][3] = l_cell_wire[85];							inform_L[83][3] = l_cell_wire[86];							inform_L[91][3] = l_cell_wire[87];							inform_L[84][3] = l_cell_wire[88];							inform_L[92][3] = l_cell_wire[89];							inform_L[85][3] = l_cell_wire[90];							inform_L[93][3] = l_cell_wire[91];							inform_L[86][3] = l_cell_wire[92];							inform_L[94][3] = l_cell_wire[93];							inform_L[87][3] = l_cell_wire[94];							inform_L[95][3] = l_cell_wire[95];							inform_L[96][3] = l_cell_wire[96];							inform_L[104][3] = l_cell_wire[97];							inform_L[97][3] = l_cell_wire[98];							inform_L[105][3] = l_cell_wire[99];							inform_L[98][3] = l_cell_wire[100];							inform_L[106][3] = l_cell_wire[101];							inform_L[99][3] = l_cell_wire[102];							inform_L[107][3] = l_cell_wire[103];							inform_L[100][3] = l_cell_wire[104];							inform_L[108][3] = l_cell_wire[105];							inform_L[101][3] = l_cell_wire[106];							inform_L[109][3] = l_cell_wire[107];							inform_L[102][3] = l_cell_wire[108];							inform_L[110][3] = l_cell_wire[109];							inform_L[103][3] = l_cell_wire[110];							inform_L[111][3] = l_cell_wire[111];							inform_L[112][3] = l_cell_wire[112];							inform_L[120][3] = l_cell_wire[113];							inform_L[113][3] = l_cell_wire[114];							inform_L[121][3] = l_cell_wire[115];							inform_L[114][3] = l_cell_wire[116];							inform_L[122][3] = l_cell_wire[117];							inform_L[115][3] = l_cell_wire[118];							inform_L[123][3] = l_cell_wire[119];							inform_L[116][3] = l_cell_wire[120];							inform_L[124][3] = l_cell_wire[121];							inform_L[117][3] = l_cell_wire[122];							inform_L[125][3] = l_cell_wire[123];							inform_L[118][3] = l_cell_wire[124];							inform_L[126][3] = l_cell_wire[125];							inform_L[119][3] = l_cell_wire[126];							inform_L[127][3] = l_cell_wire[127];							inform_L[128][3] = l_cell_wire[128];							inform_L[136][3] = l_cell_wire[129];							inform_L[129][3] = l_cell_wire[130];							inform_L[137][3] = l_cell_wire[131];							inform_L[130][3] = l_cell_wire[132];							inform_L[138][3] = l_cell_wire[133];							inform_L[131][3] = l_cell_wire[134];							inform_L[139][3] = l_cell_wire[135];							inform_L[132][3] = l_cell_wire[136];							inform_L[140][3] = l_cell_wire[137];							inform_L[133][3] = l_cell_wire[138];							inform_L[141][3] = l_cell_wire[139];							inform_L[134][3] = l_cell_wire[140];							inform_L[142][3] = l_cell_wire[141];							inform_L[135][3] = l_cell_wire[142];							inform_L[143][3] = l_cell_wire[143];							inform_L[144][3] = l_cell_wire[144];							inform_L[152][3] = l_cell_wire[145];							inform_L[145][3] = l_cell_wire[146];							inform_L[153][3] = l_cell_wire[147];							inform_L[146][3] = l_cell_wire[148];							inform_L[154][3] = l_cell_wire[149];							inform_L[147][3] = l_cell_wire[150];							inform_L[155][3] = l_cell_wire[151];							inform_L[148][3] = l_cell_wire[152];							inform_L[156][3] = l_cell_wire[153];							inform_L[149][3] = l_cell_wire[154];							inform_L[157][3] = l_cell_wire[155];							inform_L[150][3] = l_cell_wire[156];							inform_L[158][3] = l_cell_wire[157];							inform_L[151][3] = l_cell_wire[158];							inform_L[159][3] = l_cell_wire[159];							inform_L[160][3] = l_cell_wire[160];							inform_L[168][3] = l_cell_wire[161];							inform_L[161][3] = l_cell_wire[162];							inform_L[169][3] = l_cell_wire[163];							inform_L[162][3] = l_cell_wire[164];							inform_L[170][3] = l_cell_wire[165];							inform_L[163][3] = l_cell_wire[166];							inform_L[171][3] = l_cell_wire[167];							inform_L[164][3] = l_cell_wire[168];							inform_L[172][3] = l_cell_wire[169];							inform_L[165][3] = l_cell_wire[170];							inform_L[173][3] = l_cell_wire[171];							inform_L[166][3] = l_cell_wire[172];							inform_L[174][3] = l_cell_wire[173];							inform_L[167][3] = l_cell_wire[174];							inform_L[175][3] = l_cell_wire[175];							inform_L[176][3] = l_cell_wire[176];							inform_L[184][3] = l_cell_wire[177];							inform_L[177][3] = l_cell_wire[178];							inform_L[185][3] = l_cell_wire[179];							inform_L[178][3] = l_cell_wire[180];							inform_L[186][3] = l_cell_wire[181];							inform_L[179][3] = l_cell_wire[182];							inform_L[187][3] = l_cell_wire[183];							inform_L[180][3] = l_cell_wire[184];							inform_L[188][3] = l_cell_wire[185];							inform_L[181][3] = l_cell_wire[186];							inform_L[189][3] = l_cell_wire[187];							inform_L[182][3] = l_cell_wire[188];							inform_L[190][3] = l_cell_wire[189];							inform_L[183][3] = l_cell_wire[190];							inform_L[191][3] = l_cell_wire[191];							inform_L[192][3] = l_cell_wire[192];							inform_L[200][3] = l_cell_wire[193];							inform_L[193][3] = l_cell_wire[194];							inform_L[201][3] = l_cell_wire[195];							inform_L[194][3] = l_cell_wire[196];							inform_L[202][3] = l_cell_wire[197];							inform_L[195][3] = l_cell_wire[198];							inform_L[203][3] = l_cell_wire[199];							inform_L[196][3] = l_cell_wire[200];							inform_L[204][3] = l_cell_wire[201];							inform_L[197][3] = l_cell_wire[202];							inform_L[205][3] = l_cell_wire[203];							inform_L[198][3] = l_cell_wire[204];							inform_L[206][3] = l_cell_wire[205];							inform_L[199][3] = l_cell_wire[206];							inform_L[207][3] = l_cell_wire[207];							inform_L[208][3] = l_cell_wire[208];							inform_L[216][3] = l_cell_wire[209];							inform_L[209][3] = l_cell_wire[210];							inform_L[217][3] = l_cell_wire[211];							inform_L[210][3] = l_cell_wire[212];							inform_L[218][3] = l_cell_wire[213];							inform_L[211][3] = l_cell_wire[214];							inform_L[219][3] = l_cell_wire[215];							inform_L[212][3] = l_cell_wire[216];							inform_L[220][3] = l_cell_wire[217];							inform_L[213][3] = l_cell_wire[218];							inform_L[221][3] = l_cell_wire[219];							inform_L[214][3] = l_cell_wire[220];							inform_L[222][3] = l_cell_wire[221];							inform_L[215][3] = l_cell_wire[222];							inform_L[223][3] = l_cell_wire[223];							inform_L[224][3] = l_cell_wire[224];							inform_L[232][3] = l_cell_wire[225];							inform_L[225][3] = l_cell_wire[226];							inform_L[233][3] = l_cell_wire[227];							inform_L[226][3] = l_cell_wire[228];							inform_L[234][3] = l_cell_wire[229];							inform_L[227][3] = l_cell_wire[230];							inform_L[235][3] = l_cell_wire[231];							inform_L[228][3] = l_cell_wire[232];							inform_L[236][3] = l_cell_wire[233];							inform_L[229][3] = l_cell_wire[234];							inform_L[237][3] = l_cell_wire[235];							inform_L[230][3] = l_cell_wire[236];							inform_L[238][3] = l_cell_wire[237];							inform_L[231][3] = l_cell_wire[238];							inform_L[239][3] = l_cell_wire[239];							inform_L[240][3] = l_cell_wire[240];							inform_L[248][3] = l_cell_wire[241];							inform_L[241][3] = l_cell_wire[242];							inform_L[249][3] = l_cell_wire[243];							inform_L[242][3] = l_cell_wire[244];							inform_L[250][3] = l_cell_wire[245];							inform_L[243][3] = l_cell_wire[246];							inform_L[251][3] = l_cell_wire[247];							inform_L[244][3] = l_cell_wire[248];							inform_L[252][3] = l_cell_wire[249];							inform_L[245][3] = l_cell_wire[250];							inform_L[253][3] = l_cell_wire[251];							inform_L[246][3] = l_cell_wire[252];							inform_L[254][3] = l_cell_wire[253];							inform_L[247][3] = l_cell_wire[254];							inform_L[255][3] = l_cell_wire[255];							inform_L[256][3] = l_cell_wire[256];							inform_L[264][3] = l_cell_wire[257];							inform_L[257][3] = l_cell_wire[258];							inform_L[265][3] = l_cell_wire[259];							inform_L[258][3] = l_cell_wire[260];							inform_L[266][3] = l_cell_wire[261];							inform_L[259][3] = l_cell_wire[262];							inform_L[267][3] = l_cell_wire[263];							inform_L[260][3] = l_cell_wire[264];							inform_L[268][3] = l_cell_wire[265];							inform_L[261][3] = l_cell_wire[266];							inform_L[269][3] = l_cell_wire[267];							inform_L[262][3] = l_cell_wire[268];							inform_L[270][3] = l_cell_wire[269];							inform_L[263][3] = l_cell_wire[270];							inform_L[271][3] = l_cell_wire[271];							inform_L[272][3] = l_cell_wire[272];							inform_L[280][3] = l_cell_wire[273];							inform_L[273][3] = l_cell_wire[274];							inform_L[281][3] = l_cell_wire[275];							inform_L[274][3] = l_cell_wire[276];							inform_L[282][3] = l_cell_wire[277];							inform_L[275][3] = l_cell_wire[278];							inform_L[283][3] = l_cell_wire[279];							inform_L[276][3] = l_cell_wire[280];							inform_L[284][3] = l_cell_wire[281];							inform_L[277][3] = l_cell_wire[282];							inform_L[285][3] = l_cell_wire[283];							inform_L[278][3] = l_cell_wire[284];							inform_L[286][3] = l_cell_wire[285];							inform_L[279][3] = l_cell_wire[286];							inform_L[287][3] = l_cell_wire[287];							inform_L[288][3] = l_cell_wire[288];							inform_L[296][3] = l_cell_wire[289];							inform_L[289][3] = l_cell_wire[290];							inform_L[297][3] = l_cell_wire[291];							inform_L[290][3] = l_cell_wire[292];							inform_L[298][3] = l_cell_wire[293];							inform_L[291][3] = l_cell_wire[294];							inform_L[299][3] = l_cell_wire[295];							inform_L[292][3] = l_cell_wire[296];							inform_L[300][3] = l_cell_wire[297];							inform_L[293][3] = l_cell_wire[298];							inform_L[301][3] = l_cell_wire[299];							inform_L[294][3] = l_cell_wire[300];							inform_L[302][3] = l_cell_wire[301];							inform_L[295][3] = l_cell_wire[302];							inform_L[303][3] = l_cell_wire[303];							inform_L[304][3] = l_cell_wire[304];							inform_L[312][3] = l_cell_wire[305];							inform_L[305][3] = l_cell_wire[306];							inform_L[313][3] = l_cell_wire[307];							inform_L[306][3] = l_cell_wire[308];							inform_L[314][3] = l_cell_wire[309];							inform_L[307][3] = l_cell_wire[310];							inform_L[315][3] = l_cell_wire[311];							inform_L[308][3] = l_cell_wire[312];							inform_L[316][3] = l_cell_wire[313];							inform_L[309][3] = l_cell_wire[314];							inform_L[317][3] = l_cell_wire[315];							inform_L[310][3] = l_cell_wire[316];							inform_L[318][3] = l_cell_wire[317];							inform_L[311][3] = l_cell_wire[318];							inform_L[319][3] = l_cell_wire[319];							inform_L[320][3] = l_cell_wire[320];							inform_L[328][3] = l_cell_wire[321];							inform_L[321][3] = l_cell_wire[322];							inform_L[329][3] = l_cell_wire[323];							inform_L[322][3] = l_cell_wire[324];							inform_L[330][3] = l_cell_wire[325];							inform_L[323][3] = l_cell_wire[326];							inform_L[331][3] = l_cell_wire[327];							inform_L[324][3] = l_cell_wire[328];							inform_L[332][3] = l_cell_wire[329];							inform_L[325][3] = l_cell_wire[330];							inform_L[333][3] = l_cell_wire[331];							inform_L[326][3] = l_cell_wire[332];							inform_L[334][3] = l_cell_wire[333];							inform_L[327][3] = l_cell_wire[334];							inform_L[335][3] = l_cell_wire[335];							inform_L[336][3] = l_cell_wire[336];							inform_L[344][3] = l_cell_wire[337];							inform_L[337][3] = l_cell_wire[338];							inform_L[345][3] = l_cell_wire[339];							inform_L[338][3] = l_cell_wire[340];							inform_L[346][3] = l_cell_wire[341];							inform_L[339][3] = l_cell_wire[342];							inform_L[347][3] = l_cell_wire[343];							inform_L[340][3] = l_cell_wire[344];							inform_L[348][3] = l_cell_wire[345];							inform_L[341][3] = l_cell_wire[346];							inform_L[349][3] = l_cell_wire[347];							inform_L[342][3] = l_cell_wire[348];							inform_L[350][3] = l_cell_wire[349];							inform_L[343][3] = l_cell_wire[350];							inform_L[351][3] = l_cell_wire[351];							inform_L[352][3] = l_cell_wire[352];							inform_L[360][3] = l_cell_wire[353];							inform_L[353][3] = l_cell_wire[354];							inform_L[361][3] = l_cell_wire[355];							inform_L[354][3] = l_cell_wire[356];							inform_L[362][3] = l_cell_wire[357];							inform_L[355][3] = l_cell_wire[358];							inform_L[363][3] = l_cell_wire[359];							inform_L[356][3] = l_cell_wire[360];							inform_L[364][3] = l_cell_wire[361];							inform_L[357][3] = l_cell_wire[362];							inform_L[365][3] = l_cell_wire[363];							inform_L[358][3] = l_cell_wire[364];							inform_L[366][3] = l_cell_wire[365];							inform_L[359][3] = l_cell_wire[366];							inform_L[367][3] = l_cell_wire[367];							inform_L[368][3] = l_cell_wire[368];							inform_L[376][3] = l_cell_wire[369];							inform_L[369][3] = l_cell_wire[370];							inform_L[377][3] = l_cell_wire[371];							inform_L[370][3] = l_cell_wire[372];							inform_L[378][3] = l_cell_wire[373];							inform_L[371][3] = l_cell_wire[374];							inform_L[379][3] = l_cell_wire[375];							inform_L[372][3] = l_cell_wire[376];							inform_L[380][3] = l_cell_wire[377];							inform_L[373][3] = l_cell_wire[378];							inform_L[381][3] = l_cell_wire[379];							inform_L[374][3] = l_cell_wire[380];							inform_L[382][3] = l_cell_wire[381];							inform_L[375][3] = l_cell_wire[382];							inform_L[383][3] = l_cell_wire[383];							inform_L[384][3] = l_cell_wire[384];							inform_L[392][3] = l_cell_wire[385];							inform_L[385][3] = l_cell_wire[386];							inform_L[393][3] = l_cell_wire[387];							inform_L[386][3] = l_cell_wire[388];							inform_L[394][3] = l_cell_wire[389];							inform_L[387][3] = l_cell_wire[390];							inform_L[395][3] = l_cell_wire[391];							inform_L[388][3] = l_cell_wire[392];							inform_L[396][3] = l_cell_wire[393];							inform_L[389][3] = l_cell_wire[394];							inform_L[397][3] = l_cell_wire[395];							inform_L[390][3] = l_cell_wire[396];							inform_L[398][3] = l_cell_wire[397];							inform_L[391][3] = l_cell_wire[398];							inform_L[399][3] = l_cell_wire[399];							inform_L[400][3] = l_cell_wire[400];							inform_L[408][3] = l_cell_wire[401];							inform_L[401][3] = l_cell_wire[402];							inform_L[409][3] = l_cell_wire[403];							inform_L[402][3] = l_cell_wire[404];							inform_L[410][3] = l_cell_wire[405];							inform_L[403][3] = l_cell_wire[406];							inform_L[411][3] = l_cell_wire[407];							inform_L[404][3] = l_cell_wire[408];							inform_L[412][3] = l_cell_wire[409];							inform_L[405][3] = l_cell_wire[410];							inform_L[413][3] = l_cell_wire[411];							inform_L[406][3] = l_cell_wire[412];							inform_L[414][3] = l_cell_wire[413];							inform_L[407][3] = l_cell_wire[414];							inform_L[415][3] = l_cell_wire[415];							inform_L[416][3] = l_cell_wire[416];							inform_L[424][3] = l_cell_wire[417];							inform_L[417][3] = l_cell_wire[418];							inform_L[425][3] = l_cell_wire[419];							inform_L[418][3] = l_cell_wire[420];							inform_L[426][3] = l_cell_wire[421];							inform_L[419][3] = l_cell_wire[422];							inform_L[427][3] = l_cell_wire[423];							inform_L[420][3] = l_cell_wire[424];							inform_L[428][3] = l_cell_wire[425];							inform_L[421][3] = l_cell_wire[426];							inform_L[429][3] = l_cell_wire[427];							inform_L[422][3] = l_cell_wire[428];							inform_L[430][3] = l_cell_wire[429];							inform_L[423][3] = l_cell_wire[430];							inform_L[431][3] = l_cell_wire[431];							inform_L[432][3] = l_cell_wire[432];							inform_L[440][3] = l_cell_wire[433];							inform_L[433][3] = l_cell_wire[434];							inform_L[441][3] = l_cell_wire[435];							inform_L[434][3] = l_cell_wire[436];							inform_L[442][3] = l_cell_wire[437];							inform_L[435][3] = l_cell_wire[438];							inform_L[443][3] = l_cell_wire[439];							inform_L[436][3] = l_cell_wire[440];							inform_L[444][3] = l_cell_wire[441];							inform_L[437][3] = l_cell_wire[442];							inform_L[445][3] = l_cell_wire[443];							inform_L[438][3] = l_cell_wire[444];							inform_L[446][3] = l_cell_wire[445];							inform_L[439][3] = l_cell_wire[446];							inform_L[447][3] = l_cell_wire[447];							inform_L[448][3] = l_cell_wire[448];							inform_L[456][3] = l_cell_wire[449];							inform_L[449][3] = l_cell_wire[450];							inform_L[457][3] = l_cell_wire[451];							inform_L[450][3] = l_cell_wire[452];							inform_L[458][3] = l_cell_wire[453];							inform_L[451][3] = l_cell_wire[454];							inform_L[459][3] = l_cell_wire[455];							inform_L[452][3] = l_cell_wire[456];							inform_L[460][3] = l_cell_wire[457];							inform_L[453][3] = l_cell_wire[458];							inform_L[461][3] = l_cell_wire[459];							inform_L[454][3] = l_cell_wire[460];							inform_L[462][3] = l_cell_wire[461];							inform_L[455][3] = l_cell_wire[462];							inform_L[463][3] = l_cell_wire[463];							inform_L[464][3] = l_cell_wire[464];							inform_L[472][3] = l_cell_wire[465];							inform_L[465][3] = l_cell_wire[466];							inform_L[473][3] = l_cell_wire[467];							inform_L[466][3] = l_cell_wire[468];							inform_L[474][3] = l_cell_wire[469];							inform_L[467][3] = l_cell_wire[470];							inform_L[475][3] = l_cell_wire[471];							inform_L[468][3] = l_cell_wire[472];							inform_L[476][3] = l_cell_wire[473];							inform_L[469][3] = l_cell_wire[474];							inform_L[477][3] = l_cell_wire[475];							inform_L[470][3] = l_cell_wire[476];							inform_L[478][3] = l_cell_wire[477];							inform_L[471][3] = l_cell_wire[478];							inform_L[479][3] = l_cell_wire[479];							inform_L[480][3] = l_cell_wire[480];							inform_L[488][3] = l_cell_wire[481];							inform_L[481][3] = l_cell_wire[482];							inform_L[489][3] = l_cell_wire[483];							inform_L[482][3] = l_cell_wire[484];							inform_L[490][3] = l_cell_wire[485];							inform_L[483][3] = l_cell_wire[486];							inform_L[491][3] = l_cell_wire[487];							inform_L[484][3] = l_cell_wire[488];							inform_L[492][3] = l_cell_wire[489];							inform_L[485][3] = l_cell_wire[490];							inform_L[493][3] = l_cell_wire[491];							inform_L[486][3] = l_cell_wire[492];							inform_L[494][3] = l_cell_wire[493];							inform_L[487][3] = l_cell_wire[494];							inform_L[495][3] = l_cell_wire[495];							inform_L[496][3] = l_cell_wire[496];							inform_L[504][3] = l_cell_wire[497];							inform_L[497][3] = l_cell_wire[498];							inform_L[505][3] = l_cell_wire[499];							inform_L[498][3] = l_cell_wire[500];							inform_L[506][3] = l_cell_wire[501];							inform_L[499][3] = l_cell_wire[502];							inform_L[507][3] = l_cell_wire[503];							inform_L[500][3] = l_cell_wire[504];							inform_L[508][3] = l_cell_wire[505];							inform_L[501][3] = l_cell_wire[506];							inform_L[509][3] = l_cell_wire[507];							inform_L[502][3] = l_cell_wire[508];							inform_L[510][3] = l_cell_wire[509];							inform_L[503][3] = l_cell_wire[510];							inform_L[511][3] = l_cell_wire[511];							inform_L[512][3] = l_cell_wire[512];							inform_L[520][3] = l_cell_wire[513];							inform_L[513][3] = l_cell_wire[514];							inform_L[521][3] = l_cell_wire[515];							inform_L[514][3] = l_cell_wire[516];							inform_L[522][3] = l_cell_wire[517];							inform_L[515][3] = l_cell_wire[518];							inform_L[523][3] = l_cell_wire[519];							inform_L[516][3] = l_cell_wire[520];							inform_L[524][3] = l_cell_wire[521];							inform_L[517][3] = l_cell_wire[522];							inform_L[525][3] = l_cell_wire[523];							inform_L[518][3] = l_cell_wire[524];							inform_L[526][3] = l_cell_wire[525];							inform_L[519][3] = l_cell_wire[526];							inform_L[527][3] = l_cell_wire[527];							inform_L[528][3] = l_cell_wire[528];							inform_L[536][3] = l_cell_wire[529];							inform_L[529][3] = l_cell_wire[530];							inform_L[537][3] = l_cell_wire[531];							inform_L[530][3] = l_cell_wire[532];							inform_L[538][3] = l_cell_wire[533];							inform_L[531][3] = l_cell_wire[534];							inform_L[539][3] = l_cell_wire[535];							inform_L[532][3] = l_cell_wire[536];							inform_L[540][3] = l_cell_wire[537];							inform_L[533][3] = l_cell_wire[538];							inform_L[541][3] = l_cell_wire[539];							inform_L[534][3] = l_cell_wire[540];							inform_L[542][3] = l_cell_wire[541];							inform_L[535][3] = l_cell_wire[542];							inform_L[543][3] = l_cell_wire[543];							inform_L[544][3] = l_cell_wire[544];							inform_L[552][3] = l_cell_wire[545];							inform_L[545][3] = l_cell_wire[546];							inform_L[553][3] = l_cell_wire[547];							inform_L[546][3] = l_cell_wire[548];							inform_L[554][3] = l_cell_wire[549];							inform_L[547][3] = l_cell_wire[550];							inform_L[555][3] = l_cell_wire[551];							inform_L[548][3] = l_cell_wire[552];							inform_L[556][3] = l_cell_wire[553];							inform_L[549][3] = l_cell_wire[554];							inform_L[557][3] = l_cell_wire[555];							inform_L[550][3] = l_cell_wire[556];							inform_L[558][3] = l_cell_wire[557];							inform_L[551][3] = l_cell_wire[558];							inform_L[559][3] = l_cell_wire[559];							inform_L[560][3] = l_cell_wire[560];							inform_L[568][3] = l_cell_wire[561];							inform_L[561][3] = l_cell_wire[562];							inform_L[569][3] = l_cell_wire[563];							inform_L[562][3] = l_cell_wire[564];							inform_L[570][3] = l_cell_wire[565];							inform_L[563][3] = l_cell_wire[566];							inform_L[571][3] = l_cell_wire[567];							inform_L[564][3] = l_cell_wire[568];							inform_L[572][3] = l_cell_wire[569];							inform_L[565][3] = l_cell_wire[570];							inform_L[573][3] = l_cell_wire[571];							inform_L[566][3] = l_cell_wire[572];							inform_L[574][3] = l_cell_wire[573];							inform_L[567][3] = l_cell_wire[574];							inform_L[575][3] = l_cell_wire[575];							inform_L[576][3] = l_cell_wire[576];							inform_L[584][3] = l_cell_wire[577];							inform_L[577][3] = l_cell_wire[578];							inform_L[585][3] = l_cell_wire[579];							inform_L[578][3] = l_cell_wire[580];							inform_L[586][3] = l_cell_wire[581];							inform_L[579][3] = l_cell_wire[582];							inform_L[587][3] = l_cell_wire[583];							inform_L[580][3] = l_cell_wire[584];							inform_L[588][3] = l_cell_wire[585];							inform_L[581][3] = l_cell_wire[586];							inform_L[589][3] = l_cell_wire[587];							inform_L[582][3] = l_cell_wire[588];							inform_L[590][3] = l_cell_wire[589];							inform_L[583][3] = l_cell_wire[590];							inform_L[591][3] = l_cell_wire[591];							inform_L[592][3] = l_cell_wire[592];							inform_L[600][3] = l_cell_wire[593];							inform_L[593][3] = l_cell_wire[594];							inform_L[601][3] = l_cell_wire[595];							inform_L[594][3] = l_cell_wire[596];							inform_L[602][3] = l_cell_wire[597];							inform_L[595][3] = l_cell_wire[598];							inform_L[603][3] = l_cell_wire[599];							inform_L[596][3] = l_cell_wire[600];							inform_L[604][3] = l_cell_wire[601];							inform_L[597][3] = l_cell_wire[602];							inform_L[605][3] = l_cell_wire[603];							inform_L[598][3] = l_cell_wire[604];							inform_L[606][3] = l_cell_wire[605];							inform_L[599][3] = l_cell_wire[606];							inform_L[607][3] = l_cell_wire[607];							inform_L[608][3] = l_cell_wire[608];							inform_L[616][3] = l_cell_wire[609];							inform_L[609][3] = l_cell_wire[610];							inform_L[617][3] = l_cell_wire[611];							inform_L[610][3] = l_cell_wire[612];							inform_L[618][3] = l_cell_wire[613];							inform_L[611][3] = l_cell_wire[614];							inform_L[619][3] = l_cell_wire[615];							inform_L[612][3] = l_cell_wire[616];							inform_L[620][3] = l_cell_wire[617];							inform_L[613][3] = l_cell_wire[618];							inform_L[621][3] = l_cell_wire[619];							inform_L[614][3] = l_cell_wire[620];							inform_L[622][3] = l_cell_wire[621];							inform_L[615][3] = l_cell_wire[622];							inform_L[623][3] = l_cell_wire[623];							inform_L[624][3] = l_cell_wire[624];							inform_L[632][3] = l_cell_wire[625];							inform_L[625][3] = l_cell_wire[626];							inform_L[633][3] = l_cell_wire[627];							inform_L[626][3] = l_cell_wire[628];							inform_L[634][3] = l_cell_wire[629];							inform_L[627][3] = l_cell_wire[630];							inform_L[635][3] = l_cell_wire[631];							inform_L[628][3] = l_cell_wire[632];							inform_L[636][3] = l_cell_wire[633];							inform_L[629][3] = l_cell_wire[634];							inform_L[637][3] = l_cell_wire[635];							inform_L[630][3] = l_cell_wire[636];							inform_L[638][3] = l_cell_wire[637];							inform_L[631][3] = l_cell_wire[638];							inform_L[639][3] = l_cell_wire[639];							inform_L[640][3] = l_cell_wire[640];							inform_L[648][3] = l_cell_wire[641];							inform_L[641][3] = l_cell_wire[642];							inform_L[649][3] = l_cell_wire[643];							inform_L[642][3] = l_cell_wire[644];							inform_L[650][3] = l_cell_wire[645];							inform_L[643][3] = l_cell_wire[646];							inform_L[651][3] = l_cell_wire[647];							inform_L[644][3] = l_cell_wire[648];							inform_L[652][3] = l_cell_wire[649];							inform_L[645][3] = l_cell_wire[650];							inform_L[653][3] = l_cell_wire[651];							inform_L[646][3] = l_cell_wire[652];							inform_L[654][3] = l_cell_wire[653];							inform_L[647][3] = l_cell_wire[654];							inform_L[655][3] = l_cell_wire[655];							inform_L[656][3] = l_cell_wire[656];							inform_L[664][3] = l_cell_wire[657];							inform_L[657][3] = l_cell_wire[658];							inform_L[665][3] = l_cell_wire[659];							inform_L[658][3] = l_cell_wire[660];							inform_L[666][3] = l_cell_wire[661];							inform_L[659][3] = l_cell_wire[662];							inform_L[667][3] = l_cell_wire[663];							inform_L[660][3] = l_cell_wire[664];							inform_L[668][3] = l_cell_wire[665];							inform_L[661][3] = l_cell_wire[666];							inform_L[669][3] = l_cell_wire[667];							inform_L[662][3] = l_cell_wire[668];							inform_L[670][3] = l_cell_wire[669];							inform_L[663][3] = l_cell_wire[670];							inform_L[671][3] = l_cell_wire[671];							inform_L[672][3] = l_cell_wire[672];							inform_L[680][3] = l_cell_wire[673];							inform_L[673][3] = l_cell_wire[674];							inform_L[681][3] = l_cell_wire[675];							inform_L[674][3] = l_cell_wire[676];							inform_L[682][3] = l_cell_wire[677];							inform_L[675][3] = l_cell_wire[678];							inform_L[683][3] = l_cell_wire[679];							inform_L[676][3] = l_cell_wire[680];							inform_L[684][3] = l_cell_wire[681];							inform_L[677][3] = l_cell_wire[682];							inform_L[685][3] = l_cell_wire[683];							inform_L[678][3] = l_cell_wire[684];							inform_L[686][3] = l_cell_wire[685];							inform_L[679][3] = l_cell_wire[686];							inform_L[687][3] = l_cell_wire[687];							inform_L[688][3] = l_cell_wire[688];							inform_L[696][3] = l_cell_wire[689];							inform_L[689][3] = l_cell_wire[690];							inform_L[697][3] = l_cell_wire[691];							inform_L[690][3] = l_cell_wire[692];							inform_L[698][3] = l_cell_wire[693];							inform_L[691][3] = l_cell_wire[694];							inform_L[699][3] = l_cell_wire[695];							inform_L[692][3] = l_cell_wire[696];							inform_L[700][3] = l_cell_wire[697];							inform_L[693][3] = l_cell_wire[698];							inform_L[701][3] = l_cell_wire[699];							inform_L[694][3] = l_cell_wire[700];							inform_L[702][3] = l_cell_wire[701];							inform_L[695][3] = l_cell_wire[702];							inform_L[703][3] = l_cell_wire[703];							inform_L[704][3] = l_cell_wire[704];							inform_L[712][3] = l_cell_wire[705];							inform_L[705][3] = l_cell_wire[706];							inform_L[713][3] = l_cell_wire[707];							inform_L[706][3] = l_cell_wire[708];							inform_L[714][3] = l_cell_wire[709];							inform_L[707][3] = l_cell_wire[710];							inform_L[715][3] = l_cell_wire[711];							inform_L[708][3] = l_cell_wire[712];							inform_L[716][3] = l_cell_wire[713];							inform_L[709][3] = l_cell_wire[714];							inform_L[717][3] = l_cell_wire[715];							inform_L[710][3] = l_cell_wire[716];							inform_L[718][3] = l_cell_wire[717];							inform_L[711][3] = l_cell_wire[718];							inform_L[719][3] = l_cell_wire[719];							inform_L[720][3] = l_cell_wire[720];							inform_L[728][3] = l_cell_wire[721];							inform_L[721][3] = l_cell_wire[722];							inform_L[729][3] = l_cell_wire[723];							inform_L[722][3] = l_cell_wire[724];							inform_L[730][3] = l_cell_wire[725];							inform_L[723][3] = l_cell_wire[726];							inform_L[731][3] = l_cell_wire[727];							inform_L[724][3] = l_cell_wire[728];							inform_L[732][3] = l_cell_wire[729];							inform_L[725][3] = l_cell_wire[730];							inform_L[733][3] = l_cell_wire[731];							inform_L[726][3] = l_cell_wire[732];							inform_L[734][3] = l_cell_wire[733];							inform_L[727][3] = l_cell_wire[734];							inform_L[735][3] = l_cell_wire[735];							inform_L[736][3] = l_cell_wire[736];							inform_L[744][3] = l_cell_wire[737];							inform_L[737][3] = l_cell_wire[738];							inform_L[745][3] = l_cell_wire[739];							inform_L[738][3] = l_cell_wire[740];							inform_L[746][3] = l_cell_wire[741];							inform_L[739][3] = l_cell_wire[742];							inform_L[747][3] = l_cell_wire[743];							inform_L[740][3] = l_cell_wire[744];							inform_L[748][3] = l_cell_wire[745];							inform_L[741][3] = l_cell_wire[746];							inform_L[749][3] = l_cell_wire[747];							inform_L[742][3] = l_cell_wire[748];							inform_L[750][3] = l_cell_wire[749];							inform_L[743][3] = l_cell_wire[750];							inform_L[751][3] = l_cell_wire[751];							inform_L[752][3] = l_cell_wire[752];							inform_L[760][3] = l_cell_wire[753];							inform_L[753][3] = l_cell_wire[754];							inform_L[761][3] = l_cell_wire[755];							inform_L[754][3] = l_cell_wire[756];							inform_L[762][3] = l_cell_wire[757];							inform_L[755][3] = l_cell_wire[758];							inform_L[763][3] = l_cell_wire[759];							inform_L[756][3] = l_cell_wire[760];							inform_L[764][3] = l_cell_wire[761];							inform_L[757][3] = l_cell_wire[762];							inform_L[765][3] = l_cell_wire[763];							inform_L[758][3] = l_cell_wire[764];							inform_L[766][3] = l_cell_wire[765];							inform_L[759][3] = l_cell_wire[766];							inform_L[767][3] = l_cell_wire[767];							inform_L[768][3] = l_cell_wire[768];							inform_L[776][3] = l_cell_wire[769];							inform_L[769][3] = l_cell_wire[770];							inform_L[777][3] = l_cell_wire[771];							inform_L[770][3] = l_cell_wire[772];							inform_L[778][3] = l_cell_wire[773];							inform_L[771][3] = l_cell_wire[774];							inform_L[779][3] = l_cell_wire[775];							inform_L[772][3] = l_cell_wire[776];							inform_L[780][3] = l_cell_wire[777];							inform_L[773][3] = l_cell_wire[778];							inform_L[781][3] = l_cell_wire[779];							inform_L[774][3] = l_cell_wire[780];							inform_L[782][3] = l_cell_wire[781];							inform_L[775][3] = l_cell_wire[782];							inform_L[783][3] = l_cell_wire[783];							inform_L[784][3] = l_cell_wire[784];							inform_L[792][3] = l_cell_wire[785];							inform_L[785][3] = l_cell_wire[786];							inform_L[793][3] = l_cell_wire[787];							inform_L[786][3] = l_cell_wire[788];							inform_L[794][3] = l_cell_wire[789];							inform_L[787][3] = l_cell_wire[790];							inform_L[795][3] = l_cell_wire[791];							inform_L[788][3] = l_cell_wire[792];							inform_L[796][3] = l_cell_wire[793];							inform_L[789][3] = l_cell_wire[794];							inform_L[797][3] = l_cell_wire[795];							inform_L[790][3] = l_cell_wire[796];							inform_L[798][3] = l_cell_wire[797];							inform_L[791][3] = l_cell_wire[798];							inform_L[799][3] = l_cell_wire[799];							inform_L[800][3] = l_cell_wire[800];							inform_L[808][3] = l_cell_wire[801];							inform_L[801][3] = l_cell_wire[802];							inform_L[809][3] = l_cell_wire[803];							inform_L[802][3] = l_cell_wire[804];							inform_L[810][3] = l_cell_wire[805];							inform_L[803][3] = l_cell_wire[806];							inform_L[811][3] = l_cell_wire[807];							inform_L[804][3] = l_cell_wire[808];							inform_L[812][3] = l_cell_wire[809];							inform_L[805][3] = l_cell_wire[810];							inform_L[813][3] = l_cell_wire[811];							inform_L[806][3] = l_cell_wire[812];							inform_L[814][3] = l_cell_wire[813];							inform_L[807][3] = l_cell_wire[814];							inform_L[815][3] = l_cell_wire[815];							inform_L[816][3] = l_cell_wire[816];							inform_L[824][3] = l_cell_wire[817];							inform_L[817][3] = l_cell_wire[818];							inform_L[825][3] = l_cell_wire[819];							inform_L[818][3] = l_cell_wire[820];							inform_L[826][3] = l_cell_wire[821];							inform_L[819][3] = l_cell_wire[822];							inform_L[827][3] = l_cell_wire[823];							inform_L[820][3] = l_cell_wire[824];							inform_L[828][3] = l_cell_wire[825];							inform_L[821][3] = l_cell_wire[826];							inform_L[829][3] = l_cell_wire[827];							inform_L[822][3] = l_cell_wire[828];							inform_L[830][3] = l_cell_wire[829];							inform_L[823][3] = l_cell_wire[830];							inform_L[831][3] = l_cell_wire[831];							inform_L[832][3] = l_cell_wire[832];							inform_L[840][3] = l_cell_wire[833];							inform_L[833][3] = l_cell_wire[834];							inform_L[841][3] = l_cell_wire[835];							inform_L[834][3] = l_cell_wire[836];							inform_L[842][3] = l_cell_wire[837];							inform_L[835][3] = l_cell_wire[838];							inform_L[843][3] = l_cell_wire[839];							inform_L[836][3] = l_cell_wire[840];							inform_L[844][3] = l_cell_wire[841];							inform_L[837][3] = l_cell_wire[842];							inform_L[845][3] = l_cell_wire[843];							inform_L[838][3] = l_cell_wire[844];							inform_L[846][3] = l_cell_wire[845];							inform_L[839][3] = l_cell_wire[846];							inform_L[847][3] = l_cell_wire[847];							inform_L[848][3] = l_cell_wire[848];							inform_L[856][3] = l_cell_wire[849];							inform_L[849][3] = l_cell_wire[850];							inform_L[857][3] = l_cell_wire[851];							inform_L[850][3] = l_cell_wire[852];							inform_L[858][3] = l_cell_wire[853];							inform_L[851][3] = l_cell_wire[854];							inform_L[859][3] = l_cell_wire[855];							inform_L[852][3] = l_cell_wire[856];							inform_L[860][3] = l_cell_wire[857];							inform_L[853][3] = l_cell_wire[858];							inform_L[861][3] = l_cell_wire[859];							inform_L[854][3] = l_cell_wire[860];							inform_L[862][3] = l_cell_wire[861];							inform_L[855][3] = l_cell_wire[862];							inform_L[863][3] = l_cell_wire[863];							inform_L[864][3] = l_cell_wire[864];							inform_L[872][3] = l_cell_wire[865];							inform_L[865][3] = l_cell_wire[866];							inform_L[873][3] = l_cell_wire[867];							inform_L[866][3] = l_cell_wire[868];							inform_L[874][3] = l_cell_wire[869];							inform_L[867][3] = l_cell_wire[870];							inform_L[875][3] = l_cell_wire[871];							inform_L[868][3] = l_cell_wire[872];							inform_L[876][3] = l_cell_wire[873];							inform_L[869][3] = l_cell_wire[874];							inform_L[877][3] = l_cell_wire[875];							inform_L[870][3] = l_cell_wire[876];							inform_L[878][3] = l_cell_wire[877];							inform_L[871][3] = l_cell_wire[878];							inform_L[879][3] = l_cell_wire[879];							inform_L[880][3] = l_cell_wire[880];							inform_L[888][3] = l_cell_wire[881];							inform_L[881][3] = l_cell_wire[882];							inform_L[889][3] = l_cell_wire[883];							inform_L[882][3] = l_cell_wire[884];							inform_L[890][3] = l_cell_wire[885];							inform_L[883][3] = l_cell_wire[886];							inform_L[891][3] = l_cell_wire[887];							inform_L[884][3] = l_cell_wire[888];							inform_L[892][3] = l_cell_wire[889];							inform_L[885][3] = l_cell_wire[890];							inform_L[893][3] = l_cell_wire[891];							inform_L[886][3] = l_cell_wire[892];							inform_L[894][3] = l_cell_wire[893];							inform_L[887][3] = l_cell_wire[894];							inform_L[895][3] = l_cell_wire[895];							inform_L[896][3] = l_cell_wire[896];							inform_L[904][3] = l_cell_wire[897];							inform_L[897][3] = l_cell_wire[898];							inform_L[905][3] = l_cell_wire[899];							inform_L[898][3] = l_cell_wire[900];							inform_L[906][3] = l_cell_wire[901];							inform_L[899][3] = l_cell_wire[902];							inform_L[907][3] = l_cell_wire[903];							inform_L[900][3] = l_cell_wire[904];							inform_L[908][3] = l_cell_wire[905];							inform_L[901][3] = l_cell_wire[906];							inform_L[909][3] = l_cell_wire[907];							inform_L[902][3] = l_cell_wire[908];							inform_L[910][3] = l_cell_wire[909];							inform_L[903][3] = l_cell_wire[910];							inform_L[911][3] = l_cell_wire[911];							inform_L[912][3] = l_cell_wire[912];							inform_L[920][3] = l_cell_wire[913];							inform_L[913][3] = l_cell_wire[914];							inform_L[921][3] = l_cell_wire[915];							inform_L[914][3] = l_cell_wire[916];							inform_L[922][3] = l_cell_wire[917];							inform_L[915][3] = l_cell_wire[918];							inform_L[923][3] = l_cell_wire[919];							inform_L[916][3] = l_cell_wire[920];							inform_L[924][3] = l_cell_wire[921];							inform_L[917][3] = l_cell_wire[922];							inform_L[925][3] = l_cell_wire[923];							inform_L[918][3] = l_cell_wire[924];							inform_L[926][3] = l_cell_wire[925];							inform_L[919][3] = l_cell_wire[926];							inform_L[927][3] = l_cell_wire[927];							inform_L[928][3] = l_cell_wire[928];							inform_L[936][3] = l_cell_wire[929];							inform_L[929][3] = l_cell_wire[930];							inform_L[937][3] = l_cell_wire[931];							inform_L[930][3] = l_cell_wire[932];							inform_L[938][3] = l_cell_wire[933];							inform_L[931][3] = l_cell_wire[934];							inform_L[939][3] = l_cell_wire[935];							inform_L[932][3] = l_cell_wire[936];							inform_L[940][3] = l_cell_wire[937];							inform_L[933][3] = l_cell_wire[938];							inform_L[941][3] = l_cell_wire[939];							inform_L[934][3] = l_cell_wire[940];							inform_L[942][3] = l_cell_wire[941];							inform_L[935][3] = l_cell_wire[942];							inform_L[943][3] = l_cell_wire[943];							inform_L[944][3] = l_cell_wire[944];							inform_L[952][3] = l_cell_wire[945];							inform_L[945][3] = l_cell_wire[946];							inform_L[953][3] = l_cell_wire[947];							inform_L[946][3] = l_cell_wire[948];							inform_L[954][3] = l_cell_wire[949];							inform_L[947][3] = l_cell_wire[950];							inform_L[955][3] = l_cell_wire[951];							inform_L[948][3] = l_cell_wire[952];							inform_L[956][3] = l_cell_wire[953];							inform_L[949][3] = l_cell_wire[954];							inform_L[957][3] = l_cell_wire[955];							inform_L[950][3] = l_cell_wire[956];							inform_L[958][3] = l_cell_wire[957];							inform_L[951][3] = l_cell_wire[958];							inform_L[959][3] = l_cell_wire[959];							inform_L[960][3] = l_cell_wire[960];							inform_L[968][3] = l_cell_wire[961];							inform_L[961][3] = l_cell_wire[962];							inform_L[969][3] = l_cell_wire[963];							inform_L[962][3] = l_cell_wire[964];							inform_L[970][3] = l_cell_wire[965];							inform_L[963][3] = l_cell_wire[966];							inform_L[971][3] = l_cell_wire[967];							inform_L[964][3] = l_cell_wire[968];							inform_L[972][3] = l_cell_wire[969];							inform_L[965][3] = l_cell_wire[970];							inform_L[973][3] = l_cell_wire[971];							inform_L[966][3] = l_cell_wire[972];							inform_L[974][3] = l_cell_wire[973];							inform_L[967][3] = l_cell_wire[974];							inform_L[975][3] = l_cell_wire[975];							inform_L[976][3] = l_cell_wire[976];							inform_L[984][3] = l_cell_wire[977];							inform_L[977][3] = l_cell_wire[978];							inform_L[985][3] = l_cell_wire[979];							inform_L[978][3] = l_cell_wire[980];							inform_L[986][3] = l_cell_wire[981];							inform_L[979][3] = l_cell_wire[982];							inform_L[987][3] = l_cell_wire[983];							inform_L[980][3] = l_cell_wire[984];							inform_L[988][3] = l_cell_wire[985];							inform_L[981][3] = l_cell_wire[986];							inform_L[989][3] = l_cell_wire[987];							inform_L[982][3] = l_cell_wire[988];							inform_L[990][3] = l_cell_wire[989];							inform_L[983][3] = l_cell_wire[990];							inform_L[991][3] = l_cell_wire[991];							inform_L[992][3] = l_cell_wire[992];							inform_L[1000][3] = l_cell_wire[993];							inform_L[993][3] = l_cell_wire[994];							inform_L[1001][3] = l_cell_wire[995];							inform_L[994][3] = l_cell_wire[996];							inform_L[1002][3] = l_cell_wire[997];							inform_L[995][3] = l_cell_wire[998];							inform_L[1003][3] = l_cell_wire[999];							inform_L[996][3] = l_cell_wire[1000];							inform_L[1004][3] = l_cell_wire[1001];							inform_L[997][3] = l_cell_wire[1002];							inform_L[1005][3] = l_cell_wire[1003];							inform_L[998][3] = l_cell_wire[1004];							inform_L[1006][3] = l_cell_wire[1005];							inform_L[999][3] = l_cell_wire[1006];							inform_L[1007][3] = l_cell_wire[1007];							inform_L[1008][3] = l_cell_wire[1008];							inform_L[1016][3] = l_cell_wire[1009];							inform_L[1009][3] = l_cell_wire[1010];							inform_L[1017][3] = l_cell_wire[1011];							inform_L[1010][3] = l_cell_wire[1012];							inform_L[1018][3] = l_cell_wire[1013];							inform_L[1011][3] = l_cell_wire[1014];							inform_L[1019][3] = l_cell_wire[1015];							inform_L[1012][3] = l_cell_wire[1016];							inform_L[1020][3] = l_cell_wire[1017];							inform_L[1013][3] = l_cell_wire[1018];							inform_L[1021][3] = l_cell_wire[1019];							inform_L[1014][3] = l_cell_wire[1020];							inform_L[1022][3] = l_cell_wire[1021];							inform_L[1015][3] = l_cell_wire[1022];							inform_L[1023][3] = l_cell_wire[1023];						end
						5:						begin							inform_R[0][5] = r_cell_wire[0];							inform_R[16][5] = r_cell_wire[1];							inform_R[1][5] = r_cell_wire[2];							inform_R[17][5] = r_cell_wire[3];							inform_R[2][5] = r_cell_wire[4];							inform_R[18][5] = r_cell_wire[5];							inform_R[3][5] = r_cell_wire[6];							inform_R[19][5] = r_cell_wire[7];							inform_R[4][5] = r_cell_wire[8];							inform_R[20][5] = r_cell_wire[9];							inform_R[5][5] = r_cell_wire[10];							inform_R[21][5] = r_cell_wire[11];							inform_R[6][5] = r_cell_wire[12];							inform_R[22][5] = r_cell_wire[13];							inform_R[7][5] = r_cell_wire[14];							inform_R[23][5] = r_cell_wire[15];							inform_R[8][5] = r_cell_wire[16];							inform_R[24][5] = r_cell_wire[17];							inform_R[9][5] = r_cell_wire[18];							inform_R[25][5] = r_cell_wire[19];							inform_R[10][5] = r_cell_wire[20];							inform_R[26][5] = r_cell_wire[21];							inform_R[11][5] = r_cell_wire[22];							inform_R[27][5] = r_cell_wire[23];							inform_R[12][5] = r_cell_wire[24];							inform_R[28][5] = r_cell_wire[25];							inform_R[13][5] = r_cell_wire[26];							inform_R[29][5] = r_cell_wire[27];							inform_R[14][5] = r_cell_wire[28];							inform_R[30][5] = r_cell_wire[29];							inform_R[15][5] = r_cell_wire[30];							inform_R[31][5] = r_cell_wire[31];							inform_R[32][5] = r_cell_wire[32];							inform_R[48][5] = r_cell_wire[33];							inform_R[33][5] = r_cell_wire[34];							inform_R[49][5] = r_cell_wire[35];							inform_R[34][5] = r_cell_wire[36];							inform_R[50][5] = r_cell_wire[37];							inform_R[35][5] = r_cell_wire[38];							inform_R[51][5] = r_cell_wire[39];							inform_R[36][5] = r_cell_wire[40];							inform_R[52][5] = r_cell_wire[41];							inform_R[37][5] = r_cell_wire[42];							inform_R[53][5] = r_cell_wire[43];							inform_R[38][5] = r_cell_wire[44];							inform_R[54][5] = r_cell_wire[45];							inform_R[39][5] = r_cell_wire[46];							inform_R[55][5] = r_cell_wire[47];							inform_R[40][5] = r_cell_wire[48];							inform_R[56][5] = r_cell_wire[49];							inform_R[41][5] = r_cell_wire[50];							inform_R[57][5] = r_cell_wire[51];							inform_R[42][5] = r_cell_wire[52];							inform_R[58][5] = r_cell_wire[53];							inform_R[43][5] = r_cell_wire[54];							inform_R[59][5] = r_cell_wire[55];							inform_R[44][5] = r_cell_wire[56];							inform_R[60][5] = r_cell_wire[57];							inform_R[45][5] = r_cell_wire[58];							inform_R[61][5] = r_cell_wire[59];							inform_R[46][5] = r_cell_wire[60];							inform_R[62][5] = r_cell_wire[61];							inform_R[47][5] = r_cell_wire[62];							inform_R[63][5] = r_cell_wire[63];							inform_R[64][5] = r_cell_wire[64];							inform_R[80][5] = r_cell_wire[65];							inform_R[65][5] = r_cell_wire[66];							inform_R[81][5] = r_cell_wire[67];							inform_R[66][5] = r_cell_wire[68];							inform_R[82][5] = r_cell_wire[69];							inform_R[67][5] = r_cell_wire[70];							inform_R[83][5] = r_cell_wire[71];							inform_R[68][5] = r_cell_wire[72];							inform_R[84][5] = r_cell_wire[73];							inform_R[69][5] = r_cell_wire[74];							inform_R[85][5] = r_cell_wire[75];							inform_R[70][5] = r_cell_wire[76];							inform_R[86][5] = r_cell_wire[77];							inform_R[71][5] = r_cell_wire[78];							inform_R[87][5] = r_cell_wire[79];							inform_R[72][5] = r_cell_wire[80];							inform_R[88][5] = r_cell_wire[81];							inform_R[73][5] = r_cell_wire[82];							inform_R[89][5] = r_cell_wire[83];							inform_R[74][5] = r_cell_wire[84];							inform_R[90][5] = r_cell_wire[85];							inform_R[75][5] = r_cell_wire[86];							inform_R[91][5] = r_cell_wire[87];							inform_R[76][5] = r_cell_wire[88];							inform_R[92][5] = r_cell_wire[89];							inform_R[77][5] = r_cell_wire[90];							inform_R[93][5] = r_cell_wire[91];							inform_R[78][5] = r_cell_wire[92];							inform_R[94][5] = r_cell_wire[93];							inform_R[79][5] = r_cell_wire[94];							inform_R[95][5] = r_cell_wire[95];							inform_R[96][5] = r_cell_wire[96];							inform_R[112][5] = r_cell_wire[97];							inform_R[97][5] = r_cell_wire[98];							inform_R[113][5] = r_cell_wire[99];							inform_R[98][5] = r_cell_wire[100];							inform_R[114][5] = r_cell_wire[101];							inform_R[99][5] = r_cell_wire[102];							inform_R[115][5] = r_cell_wire[103];							inform_R[100][5] = r_cell_wire[104];							inform_R[116][5] = r_cell_wire[105];							inform_R[101][5] = r_cell_wire[106];							inform_R[117][5] = r_cell_wire[107];							inform_R[102][5] = r_cell_wire[108];							inform_R[118][5] = r_cell_wire[109];							inform_R[103][5] = r_cell_wire[110];							inform_R[119][5] = r_cell_wire[111];							inform_R[104][5] = r_cell_wire[112];							inform_R[120][5] = r_cell_wire[113];							inform_R[105][5] = r_cell_wire[114];							inform_R[121][5] = r_cell_wire[115];							inform_R[106][5] = r_cell_wire[116];							inform_R[122][5] = r_cell_wire[117];							inform_R[107][5] = r_cell_wire[118];							inform_R[123][5] = r_cell_wire[119];							inform_R[108][5] = r_cell_wire[120];							inform_R[124][5] = r_cell_wire[121];							inform_R[109][5] = r_cell_wire[122];							inform_R[125][5] = r_cell_wire[123];							inform_R[110][5] = r_cell_wire[124];							inform_R[126][5] = r_cell_wire[125];							inform_R[111][5] = r_cell_wire[126];							inform_R[127][5] = r_cell_wire[127];							inform_R[128][5] = r_cell_wire[128];							inform_R[144][5] = r_cell_wire[129];							inform_R[129][5] = r_cell_wire[130];							inform_R[145][5] = r_cell_wire[131];							inform_R[130][5] = r_cell_wire[132];							inform_R[146][5] = r_cell_wire[133];							inform_R[131][5] = r_cell_wire[134];							inform_R[147][5] = r_cell_wire[135];							inform_R[132][5] = r_cell_wire[136];							inform_R[148][5] = r_cell_wire[137];							inform_R[133][5] = r_cell_wire[138];							inform_R[149][5] = r_cell_wire[139];							inform_R[134][5] = r_cell_wire[140];							inform_R[150][5] = r_cell_wire[141];							inform_R[135][5] = r_cell_wire[142];							inform_R[151][5] = r_cell_wire[143];							inform_R[136][5] = r_cell_wire[144];							inform_R[152][5] = r_cell_wire[145];							inform_R[137][5] = r_cell_wire[146];							inform_R[153][5] = r_cell_wire[147];							inform_R[138][5] = r_cell_wire[148];							inform_R[154][5] = r_cell_wire[149];							inform_R[139][5] = r_cell_wire[150];							inform_R[155][5] = r_cell_wire[151];							inform_R[140][5] = r_cell_wire[152];							inform_R[156][5] = r_cell_wire[153];							inform_R[141][5] = r_cell_wire[154];							inform_R[157][5] = r_cell_wire[155];							inform_R[142][5] = r_cell_wire[156];							inform_R[158][5] = r_cell_wire[157];							inform_R[143][5] = r_cell_wire[158];							inform_R[159][5] = r_cell_wire[159];							inform_R[160][5] = r_cell_wire[160];							inform_R[176][5] = r_cell_wire[161];							inform_R[161][5] = r_cell_wire[162];							inform_R[177][5] = r_cell_wire[163];							inform_R[162][5] = r_cell_wire[164];							inform_R[178][5] = r_cell_wire[165];							inform_R[163][5] = r_cell_wire[166];							inform_R[179][5] = r_cell_wire[167];							inform_R[164][5] = r_cell_wire[168];							inform_R[180][5] = r_cell_wire[169];							inform_R[165][5] = r_cell_wire[170];							inform_R[181][5] = r_cell_wire[171];							inform_R[166][5] = r_cell_wire[172];							inform_R[182][5] = r_cell_wire[173];							inform_R[167][5] = r_cell_wire[174];							inform_R[183][5] = r_cell_wire[175];							inform_R[168][5] = r_cell_wire[176];							inform_R[184][5] = r_cell_wire[177];							inform_R[169][5] = r_cell_wire[178];							inform_R[185][5] = r_cell_wire[179];							inform_R[170][5] = r_cell_wire[180];							inform_R[186][5] = r_cell_wire[181];							inform_R[171][5] = r_cell_wire[182];							inform_R[187][5] = r_cell_wire[183];							inform_R[172][5] = r_cell_wire[184];							inform_R[188][5] = r_cell_wire[185];							inform_R[173][5] = r_cell_wire[186];							inform_R[189][5] = r_cell_wire[187];							inform_R[174][5] = r_cell_wire[188];							inform_R[190][5] = r_cell_wire[189];							inform_R[175][5] = r_cell_wire[190];							inform_R[191][5] = r_cell_wire[191];							inform_R[192][5] = r_cell_wire[192];							inform_R[208][5] = r_cell_wire[193];							inform_R[193][5] = r_cell_wire[194];							inform_R[209][5] = r_cell_wire[195];							inform_R[194][5] = r_cell_wire[196];							inform_R[210][5] = r_cell_wire[197];							inform_R[195][5] = r_cell_wire[198];							inform_R[211][5] = r_cell_wire[199];							inform_R[196][5] = r_cell_wire[200];							inform_R[212][5] = r_cell_wire[201];							inform_R[197][5] = r_cell_wire[202];							inform_R[213][5] = r_cell_wire[203];							inform_R[198][5] = r_cell_wire[204];							inform_R[214][5] = r_cell_wire[205];							inform_R[199][5] = r_cell_wire[206];							inform_R[215][5] = r_cell_wire[207];							inform_R[200][5] = r_cell_wire[208];							inform_R[216][5] = r_cell_wire[209];							inform_R[201][5] = r_cell_wire[210];							inform_R[217][5] = r_cell_wire[211];							inform_R[202][5] = r_cell_wire[212];							inform_R[218][5] = r_cell_wire[213];							inform_R[203][5] = r_cell_wire[214];							inform_R[219][5] = r_cell_wire[215];							inform_R[204][5] = r_cell_wire[216];							inform_R[220][5] = r_cell_wire[217];							inform_R[205][5] = r_cell_wire[218];							inform_R[221][5] = r_cell_wire[219];							inform_R[206][5] = r_cell_wire[220];							inform_R[222][5] = r_cell_wire[221];							inform_R[207][5] = r_cell_wire[222];							inform_R[223][5] = r_cell_wire[223];							inform_R[224][5] = r_cell_wire[224];							inform_R[240][5] = r_cell_wire[225];							inform_R[225][5] = r_cell_wire[226];							inform_R[241][5] = r_cell_wire[227];							inform_R[226][5] = r_cell_wire[228];							inform_R[242][5] = r_cell_wire[229];							inform_R[227][5] = r_cell_wire[230];							inform_R[243][5] = r_cell_wire[231];							inform_R[228][5] = r_cell_wire[232];							inform_R[244][5] = r_cell_wire[233];							inform_R[229][5] = r_cell_wire[234];							inform_R[245][5] = r_cell_wire[235];							inform_R[230][5] = r_cell_wire[236];							inform_R[246][5] = r_cell_wire[237];							inform_R[231][5] = r_cell_wire[238];							inform_R[247][5] = r_cell_wire[239];							inform_R[232][5] = r_cell_wire[240];							inform_R[248][5] = r_cell_wire[241];							inform_R[233][5] = r_cell_wire[242];							inform_R[249][5] = r_cell_wire[243];							inform_R[234][5] = r_cell_wire[244];							inform_R[250][5] = r_cell_wire[245];							inform_R[235][5] = r_cell_wire[246];							inform_R[251][5] = r_cell_wire[247];							inform_R[236][5] = r_cell_wire[248];							inform_R[252][5] = r_cell_wire[249];							inform_R[237][5] = r_cell_wire[250];							inform_R[253][5] = r_cell_wire[251];							inform_R[238][5] = r_cell_wire[252];							inform_R[254][5] = r_cell_wire[253];							inform_R[239][5] = r_cell_wire[254];							inform_R[255][5] = r_cell_wire[255];							inform_R[256][5] = r_cell_wire[256];							inform_R[272][5] = r_cell_wire[257];							inform_R[257][5] = r_cell_wire[258];							inform_R[273][5] = r_cell_wire[259];							inform_R[258][5] = r_cell_wire[260];							inform_R[274][5] = r_cell_wire[261];							inform_R[259][5] = r_cell_wire[262];							inform_R[275][5] = r_cell_wire[263];							inform_R[260][5] = r_cell_wire[264];							inform_R[276][5] = r_cell_wire[265];							inform_R[261][5] = r_cell_wire[266];							inform_R[277][5] = r_cell_wire[267];							inform_R[262][5] = r_cell_wire[268];							inform_R[278][5] = r_cell_wire[269];							inform_R[263][5] = r_cell_wire[270];							inform_R[279][5] = r_cell_wire[271];							inform_R[264][5] = r_cell_wire[272];							inform_R[280][5] = r_cell_wire[273];							inform_R[265][5] = r_cell_wire[274];							inform_R[281][5] = r_cell_wire[275];							inform_R[266][5] = r_cell_wire[276];							inform_R[282][5] = r_cell_wire[277];							inform_R[267][5] = r_cell_wire[278];							inform_R[283][5] = r_cell_wire[279];							inform_R[268][5] = r_cell_wire[280];							inform_R[284][5] = r_cell_wire[281];							inform_R[269][5] = r_cell_wire[282];							inform_R[285][5] = r_cell_wire[283];							inform_R[270][5] = r_cell_wire[284];							inform_R[286][5] = r_cell_wire[285];							inform_R[271][5] = r_cell_wire[286];							inform_R[287][5] = r_cell_wire[287];							inform_R[288][5] = r_cell_wire[288];							inform_R[304][5] = r_cell_wire[289];							inform_R[289][5] = r_cell_wire[290];							inform_R[305][5] = r_cell_wire[291];							inform_R[290][5] = r_cell_wire[292];							inform_R[306][5] = r_cell_wire[293];							inform_R[291][5] = r_cell_wire[294];							inform_R[307][5] = r_cell_wire[295];							inform_R[292][5] = r_cell_wire[296];							inform_R[308][5] = r_cell_wire[297];							inform_R[293][5] = r_cell_wire[298];							inform_R[309][5] = r_cell_wire[299];							inform_R[294][5] = r_cell_wire[300];							inform_R[310][5] = r_cell_wire[301];							inform_R[295][5] = r_cell_wire[302];							inform_R[311][5] = r_cell_wire[303];							inform_R[296][5] = r_cell_wire[304];							inform_R[312][5] = r_cell_wire[305];							inform_R[297][5] = r_cell_wire[306];							inform_R[313][5] = r_cell_wire[307];							inform_R[298][5] = r_cell_wire[308];							inform_R[314][5] = r_cell_wire[309];							inform_R[299][5] = r_cell_wire[310];							inform_R[315][5] = r_cell_wire[311];							inform_R[300][5] = r_cell_wire[312];							inform_R[316][5] = r_cell_wire[313];							inform_R[301][5] = r_cell_wire[314];							inform_R[317][5] = r_cell_wire[315];							inform_R[302][5] = r_cell_wire[316];							inform_R[318][5] = r_cell_wire[317];							inform_R[303][5] = r_cell_wire[318];							inform_R[319][5] = r_cell_wire[319];							inform_R[320][5] = r_cell_wire[320];							inform_R[336][5] = r_cell_wire[321];							inform_R[321][5] = r_cell_wire[322];							inform_R[337][5] = r_cell_wire[323];							inform_R[322][5] = r_cell_wire[324];							inform_R[338][5] = r_cell_wire[325];							inform_R[323][5] = r_cell_wire[326];							inform_R[339][5] = r_cell_wire[327];							inform_R[324][5] = r_cell_wire[328];							inform_R[340][5] = r_cell_wire[329];							inform_R[325][5] = r_cell_wire[330];							inform_R[341][5] = r_cell_wire[331];							inform_R[326][5] = r_cell_wire[332];							inform_R[342][5] = r_cell_wire[333];							inform_R[327][5] = r_cell_wire[334];							inform_R[343][5] = r_cell_wire[335];							inform_R[328][5] = r_cell_wire[336];							inform_R[344][5] = r_cell_wire[337];							inform_R[329][5] = r_cell_wire[338];							inform_R[345][5] = r_cell_wire[339];							inform_R[330][5] = r_cell_wire[340];							inform_R[346][5] = r_cell_wire[341];							inform_R[331][5] = r_cell_wire[342];							inform_R[347][5] = r_cell_wire[343];							inform_R[332][5] = r_cell_wire[344];							inform_R[348][5] = r_cell_wire[345];							inform_R[333][5] = r_cell_wire[346];							inform_R[349][5] = r_cell_wire[347];							inform_R[334][5] = r_cell_wire[348];							inform_R[350][5] = r_cell_wire[349];							inform_R[335][5] = r_cell_wire[350];							inform_R[351][5] = r_cell_wire[351];							inform_R[352][5] = r_cell_wire[352];							inform_R[368][5] = r_cell_wire[353];							inform_R[353][5] = r_cell_wire[354];							inform_R[369][5] = r_cell_wire[355];							inform_R[354][5] = r_cell_wire[356];							inform_R[370][5] = r_cell_wire[357];							inform_R[355][5] = r_cell_wire[358];							inform_R[371][5] = r_cell_wire[359];							inform_R[356][5] = r_cell_wire[360];							inform_R[372][5] = r_cell_wire[361];							inform_R[357][5] = r_cell_wire[362];							inform_R[373][5] = r_cell_wire[363];							inform_R[358][5] = r_cell_wire[364];							inform_R[374][5] = r_cell_wire[365];							inform_R[359][5] = r_cell_wire[366];							inform_R[375][5] = r_cell_wire[367];							inform_R[360][5] = r_cell_wire[368];							inform_R[376][5] = r_cell_wire[369];							inform_R[361][5] = r_cell_wire[370];							inform_R[377][5] = r_cell_wire[371];							inform_R[362][5] = r_cell_wire[372];							inform_R[378][5] = r_cell_wire[373];							inform_R[363][5] = r_cell_wire[374];							inform_R[379][5] = r_cell_wire[375];							inform_R[364][5] = r_cell_wire[376];							inform_R[380][5] = r_cell_wire[377];							inform_R[365][5] = r_cell_wire[378];							inform_R[381][5] = r_cell_wire[379];							inform_R[366][5] = r_cell_wire[380];							inform_R[382][5] = r_cell_wire[381];							inform_R[367][5] = r_cell_wire[382];							inform_R[383][5] = r_cell_wire[383];							inform_R[384][5] = r_cell_wire[384];							inform_R[400][5] = r_cell_wire[385];							inform_R[385][5] = r_cell_wire[386];							inform_R[401][5] = r_cell_wire[387];							inform_R[386][5] = r_cell_wire[388];							inform_R[402][5] = r_cell_wire[389];							inform_R[387][5] = r_cell_wire[390];							inform_R[403][5] = r_cell_wire[391];							inform_R[388][5] = r_cell_wire[392];							inform_R[404][5] = r_cell_wire[393];							inform_R[389][5] = r_cell_wire[394];							inform_R[405][5] = r_cell_wire[395];							inform_R[390][5] = r_cell_wire[396];							inform_R[406][5] = r_cell_wire[397];							inform_R[391][5] = r_cell_wire[398];							inform_R[407][5] = r_cell_wire[399];							inform_R[392][5] = r_cell_wire[400];							inform_R[408][5] = r_cell_wire[401];							inform_R[393][5] = r_cell_wire[402];							inform_R[409][5] = r_cell_wire[403];							inform_R[394][5] = r_cell_wire[404];							inform_R[410][5] = r_cell_wire[405];							inform_R[395][5] = r_cell_wire[406];							inform_R[411][5] = r_cell_wire[407];							inform_R[396][5] = r_cell_wire[408];							inform_R[412][5] = r_cell_wire[409];							inform_R[397][5] = r_cell_wire[410];							inform_R[413][5] = r_cell_wire[411];							inform_R[398][5] = r_cell_wire[412];							inform_R[414][5] = r_cell_wire[413];							inform_R[399][5] = r_cell_wire[414];							inform_R[415][5] = r_cell_wire[415];							inform_R[416][5] = r_cell_wire[416];							inform_R[432][5] = r_cell_wire[417];							inform_R[417][5] = r_cell_wire[418];							inform_R[433][5] = r_cell_wire[419];							inform_R[418][5] = r_cell_wire[420];							inform_R[434][5] = r_cell_wire[421];							inform_R[419][5] = r_cell_wire[422];							inform_R[435][5] = r_cell_wire[423];							inform_R[420][5] = r_cell_wire[424];							inform_R[436][5] = r_cell_wire[425];							inform_R[421][5] = r_cell_wire[426];							inform_R[437][5] = r_cell_wire[427];							inform_R[422][5] = r_cell_wire[428];							inform_R[438][5] = r_cell_wire[429];							inform_R[423][5] = r_cell_wire[430];							inform_R[439][5] = r_cell_wire[431];							inform_R[424][5] = r_cell_wire[432];							inform_R[440][5] = r_cell_wire[433];							inform_R[425][5] = r_cell_wire[434];							inform_R[441][5] = r_cell_wire[435];							inform_R[426][5] = r_cell_wire[436];							inform_R[442][5] = r_cell_wire[437];							inform_R[427][5] = r_cell_wire[438];							inform_R[443][5] = r_cell_wire[439];							inform_R[428][5] = r_cell_wire[440];							inform_R[444][5] = r_cell_wire[441];							inform_R[429][5] = r_cell_wire[442];							inform_R[445][5] = r_cell_wire[443];							inform_R[430][5] = r_cell_wire[444];							inform_R[446][5] = r_cell_wire[445];							inform_R[431][5] = r_cell_wire[446];							inform_R[447][5] = r_cell_wire[447];							inform_R[448][5] = r_cell_wire[448];							inform_R[464][5] = r_cell_wire[449];							inform_R[449][5] = r_cell_wire[450];							inform_R[465][5] = r_cell_wire[451];							inform_R[450][5] = r_cell_wire[452];							inform_R[466][5] = r_cell_wire[453];							inform_R[451][5] = r_cell_wire[454];							inform_R[467][5] = r_cell_wire[455];							inform_R[452][5] = r_cell_wire[456];							inform_R[468][5] = r_cell_wire[457];							inform_R[453][5] = r_cell_wire[458];							inform_R[469][5] = r_cell_wire[459];							inform_R[454][5] = r_cell_wire[460];							inform_R[470][5] = r_cell_wire[461];							inform_R[455][5] = r_cell_wire[462];							inform_R[471][5] = r_cell_wire[463];							inform_R[456][5] = r_cell_wire[464];							inform_R[472][5] = r_cell_wire[465];							inform_R[457][5] = r_cell_wire[466];							inform_R[473][5] = r_cell_wire[467];							inform_R[458][5] = r_cell_wire[468];							inform_R[474][5] = r_cell_wire[469];							inform_R[459][5] = r_cell_wire[470];							inform_R[475][5] = r_cell_wire[471];							inform_R[460][5] = r_cell_wire[472];							inform_R[476][5] = r_cell_wire[473];							inform_R[461][5] = r_cell_wire[474];							inform_R[477][5] = r_cell_wire[475];							inform_R[462][5] = r_cell_wire[476];							inform_R[478][5] = r_cell_wire[477];							inform_R[463][5] = r_cell_wire[478];							inform_R[479][5] = r_cell_wire[479];							inform_R[480][5] = r_cell_wire[480];							inform_R[496][5] = r_cell_wire[481];							inform_R[481][5] = r_cell_wire[482];							inform_R[497][5] = r_cell_wire[483];							inform_R[482][5] = r_cell_wire[484];							inform_R[498][5] = r_cell_wire[485];							inform_R[483][5] = r_cell_wire[486];							inform_R[499][5] = r_cell_wire[487];							inform_R[484][5] = r_cell_wire[488];							inform_R[500][5] = r_cell_wire[489];							inform_R[485][5] = r_cell_wire[490];							inform_R[501][5] = r_cell_wire[491];							inform_R[486][5] = r_cell_wire[492];							inform_R[502][5] = r_cell_wire[493];							inform_R[487][5] = r_cell_wire[494];							inform_R[503][5] = r_cell_wire[495];							inform_R[488][5] = r_cell_wire[496];							inform_R[504][5] = r_cell_wire[497];							inform_R[489][5] = r_cell_wire[498];							inform_R[505][5] = r_cell_wire[499];							inform_R[490][5] = r_cell_wire[500];							inform_R[506][5] = r_cell_wire[501];							inform_R[491][5] = r_cell_wire[502];							inform_R[507][5] = r_cell_wire[503];							inform_R[492][5] = r_cell_wire[504];							inform_R[508][5] = r_cell_wire[505];							inform_R[493][5] = r_cell_wire[506];							inform_R[509][5] = r_cell_wire[507];							inform_R[494][5] = r_cell_wire[508];							inform_R[510][5] = r_cell_wire[509];							inform_R[495][5] = r_cell_wire[510];							inform_R[511][5] = r_cell_wire[511];							inform_R[512][5] = r_cell_wire[512];							inform_R[528][5] = r_cell_wire[513];							inform_R[513][5] = r_cell_wire[514];							inform_R[529][5] = r_cell_wire[515];							inform_R[514][5] = r_cell_wire[516];							inform_R[530][5] = r_cell_wire[517];							inform_R[515][5] = r_cell_wire[518];							inform_R[531][5] = r_cell_wire[519];							inform_R[516][5] = r_cell_wire[520];							inform_R[532][5] = r_cell_wire[521];							inform_R[517][5] = r_cell_wire[522];							inform_R[533][5] = r_cell_wire[523];							inform_R[518][5] = r_cell_wire[524];							inform_R[534][5] = r_cell_wire[525];							inform_R[519][5] = r_cell_wire[526];							inform_R[535][5] = r_cell_wire[527];							inform_R[520][5] = r_cell_wire[528];							inform_R[536][5] = r_cell_wire[529];							inform_R[521][5] = r_cell_wire[530];							inform_R[537][5] = r_cell_wire[531];							inform_R[522][5] = r_cell_wire[532];							inform_R[538][5] = r_cell_wire[533];							inform_R[523][5] = r_cell_wire[534];							inform_R[539][5] = r_cell_wire[535];							inform_R[524][5] = r_cell_wire[536];							inform_R[540][5] = r_cell_wire[537];							inform_R[525][5] = r_cell_wire[538];							inform_R[541][5] = r_cell_wire[539];							inform_R[526][5] = r_cell_wire[540];							inform_R[542][5] = r_cell_wire[541];							inform_R[527][5] = r_cell_wire[542];							inform_R[543][5] = r_cell_wire[543];							inform_R[544][5] = r_cell_wire[544];							inform_R[560][5] = r_cell_wire[545];							inform_R[545][5] = r_cell_wire[546];							inform_R[561][5] = r_cell_wire[547];							inform_R[546][5] = r_cell_wire[548];							inform_R[562][5] = r_cell_wire[549];							inform_R[547][5] = r_cell_wire[550];							inform_R[563][5] = r_cell_wire[551];							inform_R[548][5] = r_cell_wire[552];							inform_R[564][5] = r_cell_wire[553];							inform_R[549][5] = r_cell_wire[554];							inform_R[565][5] = r_cell_wire[555];							inform_R[550][5] = r_cell_wire[556];							inform_R[566][5] = r_cell_wire[557];							inform_R[551][5] = r_cell_wire[558];							inform_R[567][5] = r_cell_wire[559];							inform_R[552][5] = r_cell_wire[560];							inform_R[568][5] = r_cell_wire[561];							inform_R[553][5] = r_cell_wire[562];							inform_R[569][5] = r_cell_wire[563];							inform_R[554][5] = r_cell_wire[564];							inform_R[570][5] = r_cell_wire[565];							inform_R[555][5] = r_cell_wire[566];							inform_R[571][5] = r_cell_wire[567];							inform_R[556][5] = r_cell_wire[568];							inform_R[572][5] = r_cell_wire[569];							inform_R[557][5] = r_cell_wire[570];							inform_R[573][5] = r_cell_wire[571];							inform_R[558][5] = r_cell_wire[572];							inform_R[574][5] = r_cell_wire[573];							inform_R[559][5] = r_cell_wire[574];							inform_R[575][5] = r_cell_wire[575];							inform_R[576][5] = r_cell_wire[576];							inform_R[592][5] = r_cell_wire[577];							inform_R[577][5] = r_cell_wire[578];							inform_R[593][5] = r_cell_wire[579];							inform_R[578][5] = r_cell_wire[580];							inform_R[594][5] = r_cell_wire[581];							inform_R[579][5] = r_cell_wire[582];							inform_R[595][5] = r_cell_wire[583];							inform_R[580][5] = r_cell_wire[584];							inform_R[596][5] = r_cell_wire[585];							inform_R[581][5] = r_cell_wire[586];							inform_R[597][5] = r_cell_wire[587];							inform_R[582][5] = r_cell_wire[588];							inform_R[598][5] = r_cell_wire[589];							inform_R[583][5] = r_cell_wire[590];							inform_R[599][5] = r_cell_wire[591];							inform_R[584][5] = r_cell_wire[592];							inform_R[600][5] = r_cell_wire[593];							inform_R[585][5] = r_cell_wire[594];							inform_R[601][5] = r_cell_wire[595];							inform_R[586][5] = r_cell_wire[596];							inform_R[602][5] = r_cell_wire[597];							inform_R[587][5] = r_cell_wire[598];							inform_R[603][5] = r_cell_wire[599];							inform_R[588][5] = r_cell_wire[600];							inform_R[604][5] = r_cell_wire[601];							inform_R[589][5] = r_cell_wire[602];							inform_R[605][5] = r_cell_wire[603];							inform_R[590][5] = r_cell_wire[604];							inform_R[606][5] = r_cell_wire[605];							inform_R[591][5] = r_cell_wire[606];							inform_R[607][5] = r_cell_wire[607];							inform_R[608][5] = r_cell_wire[608];							inform_R[624][5] = r_cell_wire[609];							inform_R[609][5] = r_cell_wire[610];							inform_R[625][5] = r_cell_wire[611];							inform_R[610][5] = r_cell_wire[612];							inform_R[626][5] = r_cell_wire[613];							inform_R[611][5] = r_cell_wire[614];							inform_R[627][5] = r_cell_wire[615];							inform_R[612][5] = r_cell_wire[616];							inform_R[628][5] = r_cell_wire[617];							inform_R[613][5] = r_cell_wire[618];							inform_R[629][5] = r_cell_wire[619];							inform_R[614][5] = r_cell_wire[620];							inform_R[630][5] = r_cell_wire[621];							inform_R[615][5] = r_cell_wire[622];							inform_R[631][5] = r_cell_wire[623];							inform_R[616][5] = r_cell_wire[624];							inform_R[632][5] = r_cell_wire[625];							inform_R[617][5] = r_cell_wire[626];							inform_R[633][5] = r_cell_wire[627];							inform_R[618][5] = r_cell_wire[628];							inform_R[634][5] = r_cell_wire[629];							inform_R[619][5] = r_cell_wire[630];							inform_R[635][5] = r_cell_wire[631];							inform_R[620][5] = r_cell_wire[632];							inform_R[636][5] = r_cell_wire[633];							inform_R[621][5] = r_cell_wire[634];							inform_R[637][5] = r_cell_wire[635];							inform_R[622][5] = r_cell_wire[636];							inform_R[638][5] = r_cell_wire[637];							inform_R[623][5] = r_cell_wire[638];							inform_R[639][5] = r_cell_wire[639];							inform_R[640][5] = r_cell_wire[640];							inform_R[656][5] = r_cell_wire[641];							inform_R[641][5] = r_cell_wire[642];							inform_R[657][5] = r_cell_wire[643];							inform_R[642][5] = r_cell_wire[644];							inform_R[658][5] = r_cell_wire[645];							inform_R[643][5] = r_cell_wire[646];							inform_R[659][5] = r_cell_wire[647];							inform_R[644][5] = r_cell_wire[648];							inform_R[660][5] = r_cell_wire[649];							inform_R[645][5] = r_cell_wire[650];							inform_R[661][5] = r_cell_wire[651];							inform_R[646][5] = r_cell_wire[652];							inform_R[662][5] = r_cell_wire[653];							inform_R[647][5] = r_cell_wire[654];							inform_R[663][5] = r_cell_wire[655];							inform_R[648][5] = r_cell_wire[656];							inform_R[664][5] = r_cell_wire[657];							inform_R[649][5] = r_cell_wire[658];							inform_R[665][5] = r_cell_wire[659];							inform_R[650][5] = r_cell_wire[660];							inform_R[666][5] = r_cell_wire[661];							inform_R[651][5] = r_cell_wire[662];							inform_R[667][5] = r_cell_wire[663];							inform_R[652][5] = r_cell_wire[664];							inform_R[668][5] = r_cell_wire[665];							inform_R[653][5] = r_cell_wire[666];							inform_R[669][5] = r_cell_wire[667];							inform_R[654][5] = r_cell_wire[668];							inform_R[670][5] = r_cell_wire[669];							inform_R[655][5] = r_cell_wire[670];							inform_R[671][5] = r_cell_wire[671];							inform_R[672][5] = r_cell_wire[672];							inform_R[688][5] = r_cell_wire[673];							inform_R[673][5] = r_cell_wire[674];							inform_R[689][5] = r_cell_wire[675];							inform_R[674][5] = r_cell_wire[676];							inform_R[690][5] = r_cell_wire[677];							inform_R[675][5] = r_cell_wire[678];							inform_R[691][5] = r_cell_wire[679];							inform_R[676][5] = r_cell_wire[680];							inform_R[692][5] = r_cell_wire[681];							inform_R[677][5] = r_cell_wire[682];							inform_R[693][5] = r_cell_wire[683];							inform_R[678][5] = r_cell_wire[684];							inform_R[694][5] = r_cell_wire[685];							inform_R[679][5] = r_cell_wire[686];							inform_R[695][5] = r_cell_wire[687];							inform_R[680][5] = r_cell_wire[688];							inform_R[696][5] = r_cell_wire[689];							inform_R[681][5] = r_cell_wire[690];							inform_R[697][5] = r_cell_wire[691];							inform_R[682][5] = r_cell_wire[692];							inform_R[698][5] = r_cell_wire[693];							inform_R[683][5] = r_cell_wire[694];							inform_R[699][5] = r_cell_wire[695];							inform_R[684][5] = r_cell_wire[696];							inform_R[700][5] = r_cell_wire[697];							inform_R[685][5] = r_cell_wire[698];							inform_R[701][5] = r_cell_wire[699];							inform_R[686][5] = r_cell_wire[700];							inform_R[702][5] = r_cell_wire[701];							inform_R[687][5] = r_cell_wire[702];							inform_R[703][5] = r_cell_wire[703];							inform_R[704][5] = r_cell_wire[704];							inform_R[720][5] = r_cell_wire[705];							inform_R[705][5] = r_cell_wire[706];							inform_R[721][5] = r_cell_wire[707];							inform_R[706][5] = r_cell_wire[708];							inform_R[722][5] = r_cell_wire[709];							inform_R[707][5] = r_cell_wire[710];							inform_R[723][5] = r_cell_wire[711];							inform_R[708][5] = r_cell_wire[712];							inform_R[724][5] = r_cell_wire[713];							inform_R[709][5] = r_cell_wire[714];							inform_R[725][5] = r_cell_wire[715];							inform_R[710][5] = r_cell_wire[716];							inform_R[726][5] = r_cell_wire[717];							inform_R[711][5] = r_cell_wire[718];							inform_R[727][5] = r_cell_wire[719];							inform_R[712][5] = r_cell_wire[720];							inform_R[728][5] = r_cell_wire[721];							inform_R[713][5] = r_cell_wire[722];							inform_R[729][5] = r_cell_wire[723];							inform_R[714][5] = r_cell_wire[724];							inform_R[730][5] = r_cell_wire[725];							inform_R[715][5] = r_cell_wire[726];							inform_R[731][5] = r_cell_wire[727];							inform_R[716][5] = r_cell_wire[728];							inform_R[732][5] = r_cell_wire[729];							inform_R[717][5] = r_cell_wire[730];							inform_R[733][5] = r_cell_wire[731];							inform_R[718][5] = r_cell_wire[732];							inform_R[734][5] = r_cell_wire[733];							inform_R[719][5] = r_cell_wire[734];							inform_R[735][5] = r_cell_wire[735];							inform_R[736][5] = r_cell_wire[736];							inform_R[752][5] = r_cell_wire[737];							inform_R[737][5] = r_cell_wire[738];							inform_R[753][5] = r_cell_wire[739];							inform_R[738][5] = r_cell_wire[740];							inform_R[754][5] = r_cell_wire[741];							inform_R[739][5] = r_cell_wire[742];							inform_R[755][5] = r_cell_wire[743];							inform_R[740][5] = r_cell_wire[744];							inform_R[756][5] = r_cell_wire[745];							inform_R[741][5] = r_cell_wire[746];							inform_R[757][5] = r_cell_wire[747];							inform_R[742][5] = r_cell_wire[748];							inform_R[758][5] = r_cell_wire[749];							inform_R[743][5] = r_cell_wire[750];							inform_R[759][5] = r_cell_wire[751];							inform_R[744][5] = r_cell_wire[752];							inform_R[760][5] = r_cell_wire[753];							inform_R[745][5] = r_cell_wire[754];							inform_R[761][5] = r_cell_wire[755];							inform_R[746][5] = r_cell_wire[756];							inform_R[762][5] = r_cell_wire[757];							inform_R[747][5] = r_cell_wire[758];							inform_R[763][5] = r_cell_wire[759];							inform_R[748][5] = r_cell_wire[760];							inform_R[764][5] = r_cell_wire[761];							inform_R[749][5] = r_cell_wire[762];							inform_R[765][5] = r_cell_wire[763];							inform_R[750][5] = r_cell_wire[764];							inform_R[766][5] = r_cell_wire[765];							inform_R[751][5] = r_cell_wire[766];							inform_R[767][5] = r_cell_wire[767];							inform_R[768][5] = r_cell_wire[768];							inform_R[784][5] = r_cell_wire[769];							inform_R[769][5] = r_cell_wire[770];							inform_R[785][5] = r_cell_wire[771];							inform_R[770][5] = r_cell_wire[772];							inform_R[786][5] = r_cell_wire[773];							inform_R[771][5] = r_cell_wire[774];							inform_R[787][5] = r_cell_wire[775];							inform_R[772][5] = r_cell_wire[776];							inform_R[788][5] = r_cell_wire[777];							inform_R[773][5] = r_cell_wire[778];							inform_R[789][5] = r_cell_wire[779];							inform_R[774][5] = r_cell_wire[780];							inform_R[790][5] = r_cell_wire[781];							inform_R[775][5] = r_cell_wire[782];							inform_R[791][5] = r_cell_wire[783];							inform_R[776][5] = r_cell_wire[784];							inform_R[792][5] = r_cell_wire[785];							inform_R[777][5] = r_cell_wire[786];							inform_R[793][5] = r_cell_wire[787];							inform_R[778][5] = r_cell_wire[788];							inform_R[794][5] = r_cell_wire[789];							inform_R[779][5] = r_cell_wire[790];							inform_R[795][5] = r_cell_wire[791];							inform_R[780][5] = r_cell_wire[792];							inform_R[796][5] = r_cell_wire[793];							inform_R[781][5] = r_cell_wire[794];							inform_R[797][5] = r_cell_wire[795];							inform_R[782][5] = r_cell_wire[796];							inform_R[798][5] = r_cell_wire[797];							inform_R[783][5] = r_cell_wire[798];							inform_R[799][5] = r_cell_wire[799];							inform_R[800][5] = r_cell_wire[800];							inform_R[816][5] = r_cell_wire[801];							inform_R[801][5] = r_cell_wire[802];							inform_R[817][5] = r_cell_wire[803];							inform_R[802][5] = r_cell_wire[804];							inform_R[818][5] = r_cell_wire[805];							inform_R[803][5] = r_cell_wire[806];							inform_R[819][5] = r_cell_wire[807];							inform_R[804][5] = r_cell_wire[808];							inform_R[820][5] = r_cell_wire[809];							inform_R[805][5] = r_cell_wire[810];							inform_R[821][5] = r_cell_wire[811];							inform_R[806][5] = r_cell_wire[812];							inform_R[822][5] = r_cell_wire[813];							inform_R[807][5] = r_cell_wire[814];							inform_R[823][5] = r_cell_wire[815];							inform_R[808][5] = r_cell_wire[816];							inform_R[824][5] = r_cell_wire[817];							inform_R[809][5] = r_cell_wire[818];							inform_R[825][5] = r_cell_wire[819];							inform_R[810][5] = r_cell_wire[820];							inform_R[826][5] = r_cell_wire[821];							inform_R[811][5] = r_cell_wire[822];							inform_R[827][5] = r_cell_wire[823];							inform_R[812][5] = r_cell_wire[824];							inform_R[828][5] = r_cell_wire[825];							inform_R[813][5] = r_cell_wire[826];							inform_R[829][5] = r_cell_wire[827];							inform_R[814][5] = r_cell_wire[828];							inform_R[830][5] = r_cell_wire[829];							inform_R[815][5] = r_cell_wire[830];							inform_R[831][5] = r_cell_wire[831];							inform_R[832][5] = r_cell_wire[832];							inform_R[848][5] = r_cell_wire[833];							inform_R[833][5] = r_cell_wire[834];							inform_R[849][5] = r_cell_wire[835];							inform_R[834][5] = r_cell_wire[836];							inform_R[850][5] = r_cell_wire[837];							inform_R[835][5] = r_cell_wire[838];							inform_R[851][5] = r_cell_wire[839];							inform_R[836][5] = r_cell_wire[840];							inform_R[852][5] = r_cell_wire[841];							inform_R[837][5] = r_cell_wire[842];							inform_R[853][5] = r_cell_wire[843];							inform_R[838][5] = r_cell_wire[844];							inform_R[854][5] = r_cell_wire[845];							inform_R[839][5] = r_cell_wire[846];							inform_R[855][5] = r_cell_wire[847];							inform_R[840][5] = r_cell_wire[848];							inform_R[856][5] = r_cell_wire[849];							inform_R[841][5] = r_cell_wire[850];							inform_R[857][5] = r_cell_wire[851];							inform_R[842][5] = r_cell_wire[852];							inform_R[858][5] = r_cell_wire[853];							inform_R[843][5] = r_cell_wire[854];							inform_R[859][5] = r_cell_wire[855];							inform_R[844][5] = r_cell_wire[856];							inform_R[860][5] = r_cell_wire[857];							inform_R[845][5] = r_cell_wire[858];							inform_R[861][5] = r_cell_wire[859];							inform_R[846][5] = r_cell_wire[860];							inform_R[862][5] = r_cell_wire[861];							inform_R[847][5] = r_cell_wire[862];							inform_R[863][5] = r_cell_wire[863];							inform_R[864][5] = r_cell_wire[864];							inform_R[880][5] = r_cell_wire[865];							inform_R[865][5] = r_cell_wire[866];							inform_R[881][5] = r_cell_wire[867];							inform_R[866][5] = r_cell_wire[868];							inform_R[882][5] = r_cell_wire[869];							inform_R[867][5] = r_cell_wire[870];							inform_R[883][5] = r_cell_wire[871];							inform_R[868][5] = r_cell_wire[872];							inform_R[884][5] = r_cell_wire[873];							inform_R[869][5] = r_cell_wire[874];							inform_R[885][5] = r_cell_wire[875];							inform_R[870][5] = r_cell_wire[876];							inform_R[886][5] = r_cell_wire[877];							inform_R[871][5] = r_cell_wire[878];							inform_R[887][5] = r_cell_wire[879];							inform_R[872][5] = r_cell_wire[880];							inform_R[888][5] = r_cell_wire[881];							inform_R[873][5] = r_cell_wire[882];							inform_R[889][5] = r_cell_wire[883];							inform_R[874][5] = r_cell_wire[884];							inform_R[890][5] = r_cell_wire[885];							inform_R[875][5] = r_cell_wire[886];							inform_R[891][5] = r_cell_wire[887];							inform_R[876][5] = r_cell_wire[888];							inform_R[892][5] = r_cell_wire[889];							inform_R[877][5] = r_cell_wire[890];							inform_R[893][5] = r_cell_wire[891];							inform_R[878][5] = r_cell_wire[892];							inform_R[894][5] = r_cell_wire[893];							inform_R[879][5] = r_cell_wire[894];							inform_R[895][5] = r_cell_wire[895];							inform_R[896][5] = r_cell_wire[896];							inform_R[912][5] = r_cell_wire[897];							inform_R[897][5] = r_cell_wire[898];							inform_R[913][5] = r_cell_wire[899];							inform_R[898][5] = r_cell_wire[900];							inform_R[914][5] = r_cell_wire[901];							inform_R[899][5] = r_cell_wire[902];							inform_R[915][5] = r_cell_wire[903];							inform_R[900][5] = r_cell_wire[904];							inform_R[916][5] = r_cell_wire[905];							inform_R[901][5] = r_cell_wire[906];							inform_R[917][5] = r_cell_wire[907];							inform_R[902][5] = r_cell_wire[908];							inform_R[918][5] = r_cell_wire[909];							inform_R[903][5] = r_cell_wire[910];							inform_R[919][5] = r_cell_wire[911];							inform_R[904][5] = r_cell_wire[912];							inform_R[920][5] = r_cell_wire[913];							inform_R[905][5] = r_cell_wire[914];							inform_R[921][5] = r_cell_wire[915];							inform_R[906][5] = r_cell_wire[916];							inform_R[922][5] = r_cell_wire[917];							inform_R[907][5] = r_cell_wire[918];							inform_R[923][5] = r_cell_wire[919];							inform_R[908][5] = r_cell_wire[920];							inform_R[924][5] = r_cell_wire[921];							inform_R[909][5] = r_cell_wire[922];							inform_R[925][5] = r_cell_wire[923];							inform_R[910][5] = r_cell_wire[924];							inform_R[926][5] = r_cell_wire[925];							inform_R[911][5] = r_cell_wire[926];							inform_R[927][5] = r_cell_wire[927];							inform_R[928][5] = r_cell_wire[928];							inform_R[944][5] = r_cell_wire[929];							inform_R[929][5] = r_cell_wire[930];							inform_R[945][5] = r_cell_wire[931];							inform_R[930][5] = r_cell_wire[932];							inform_R[946][5] = r_cell_wire[933];							inform_R[931][5] = r_cell_wire[934];							inform_R[947][5] = r_cell_wire[935];							inform_R[932][5] = r_cell_wire[936];							inform_R[948][5] = r_cell_wire[937];							inform_R[933][5] = r_cell_wire[938];							inform_R[949][5] = r_cell_wire[939];							inform_R[934][5] = r_cell_wire[940];							inform_R[950][5] = r_cell_wire[941];							inform_R[935][5] = r_cell_wire[942];							inform_R[951][5] = r_cell_wire[943];							inform_R[936][5] = r_cell_wire[944];							inform_R[952][5] = r_cell_wire[945];							inform_R[937][5] = r_cell_wire[946];							inform_R[953][5] = r_cell_wire[947];							inform_R[938][5] = r_cell_wire[948];							inform_R[954][5] = r_cell_wire[949];							inform_R[939][5] = r_cell_wire[950];							inform_R[955][5] = r_cell_wire[951];							inform_R[940][5] = r_cell_wire[952];							inform_R[956][5] = r_cell_wire[953];							inform_R[941][5] = r_cell_wire[954];							inform_R[957][5] = r_cell_wire[955];							inform_R[942][5] = r_cell_wire[956];							inform_R[958][5] = r_cell_wire[957];							inform_R[943][5] = r_cell_wire[958];							inform_R[959][5] = r_cell_wire[959];							inform_R[960][5] = r_cell_wire[960];							inform_R[976][5] = r_cell_wire[961];							inform_R[961][5] = r_cell_wire[962];							inform_R[977][5] = r_cell_wire[963];							inform_R[962][5] = r_cell_wire[964];							inform_R[978][5] = r_cell_wire[965];							inform_R[963][5] = r_cell_wire[966];							inform_R[979][5] = r_cell_wire[967];							inform_R[964][5] = r_cell_wire[968];							inform_R[980][5] = r_cell_wire[969];							inform_R[965][5] = r_cell_wire[970];							inform_R[981][5] = r_cell_wire[971];							inform_R[966][5] = r_cell_wire[972];							inform_R[982][5] = r_cell_wire[973];							inform_R[967][5] = r_cell_wire[974];							inform_R[983][5] = r_cell_wire[975];							inform_R[968][5] = r_cell_wire[976];							inform_R[984][5] = r_cell_wire[977];							inform_R[969][5] = r_cell_wire[978];							inform_R[985][5] = r_cell_wire[979];							inform_R[970][5] = r_cell_wire[980];							inform_R[986][5] = r_cell_wire[981];							inform_R[971][5] = r_cell_wire[982];							inform_R[987][5] = r_cell_wire[983];							inform_R[972][5] = r_cell_wire[984];							inform_R[988][5] = r_cell_wire[985];							inform_R[973][5] = r_cell_wire[986];							inform_R[989][5] = r_cell_wire[987];							inform_R[974][5] = r_cell_wire[988];							inform_R[990][5] = r_cell_wire[989];							inform_R[975][5] = r_cell_wire[990];							inform_R[991][5] = r_cell_wire[991];							inform_R[992][5] = r_cell_wire[992];							inform_R[1008][5] = r_cell_wire[993];							inform_R[993][5] = r_cell_wire[994];							inform_R[1009][5] = r_cell_wire[995];							inform_R[994][5] = r_cell_wire[996];							inform_R[1010][5] = r_cell_wire[997];							inform_R[995][5] = r_cell_wire[998];							inform_R[1011][5] = r_cell_wire[999];							inform_R[996][5] = r_cell_wire[1000];							inform_R[1012][5] = r_cell_wire[1001];							inform_R[997][5] = r_cell_wire[1002];							inform_R[1013][5] = r_cell_wire[1003];							inform_R[998][5] = r_cell_wire[1004];							inform_R[1014][5] = r_cell_wire[1005];							inform_R[999][5] = r_cell_wire[1006];							inform_R[1015][5] = r_cell_wire[1007];							inform_R[1000][5] = r_cell_wire[1008];							inform_R[1016][5] = r_cell_wire[1009];							inform_R[1001][5] = r_cell_wire[1010];							inform_R[1017][5] = r_cell_wire[1011];							inform_R[1002][5] = r_cell_wire[1012];							inform_R[1018][5] = r_cell_wire[1013];							inform_R[1003][5] = r_cell_wire[1014];							inform_R[1019][5] = r_cell_wire[1015];							inform_R[1004][5] = r_cell_wire[1016];							inform_R[1020][5] = r_cell_wire[1017];							inform_R[1005][5] = r_cell_wire[1018];							inform_R[1021][5] = r_cell_wire[1019];							inform_R[1006][5] = r_cell_wire[1020];							inform_R[1022][5] = r_cell_wire[1021];							inform_R[1007][5] = r_cell_wire[1022];							inform_R[1023][5] = r_cell_wire[1023];							inform_L[0][4] = l_cell_wire[0];							inform_L[16][4] = l_cell_wire[1];							inform_L[1][4] = l_cell_wire[2];							inform_L[17][4] = l_cell_wire[3];							inform_L[2][4] = l_cell_wire[4];							inform_L[18][4] = l_cell_wire[5];							inform_L[3][4] = l_cell_wire[6];							inform_L[19][4] = l_cell_wire[7];							inform_L[4][4] = l_cell_wire[8];							inform_L[20][4] = l_cell_wire[9];							inform_L[5][4] = l_cell_wire[10];							inform_L[21][4] = l_cell_wire[11];							inform_L[6][4] = l_cell_wire[12];							inform_L[22][4] = l_cell_wire[13];							inform_L[7][4] = l_cell_wire[14];							inform_L[23][4] = l_cell_wire[15];							inform_L[8][4] = l_cell_wire[16];							inform_L[24][4] = l_cell_wire[17];							inform_L[9][4] = l_cell_wire[18];							inform_L[25][4] = l_cell_wire[19];							inform_L[10][4] = l_cell_wire[20];							inform_L[26][4] = l_cell_wire[21];							inform_L[11][4] = l_cell_wire[22];							inform_L[27][4] = l_cell_wire[23];							inform_L[12][4] = l_cell_wire[24];							inform_L[28][4] = l_cell_wire[25];							inform_L[13][4] = l_cell_wire[26];							inform_L[29][4] = l_cell_wire[27];							inform_L[14][4] = l_cell_wire[28];							inform_L[30][4] = l_cell_wire[29];							inform_L[15][4] = l_cell_wire[30];							inform_L[31][4] = l_cell_wire[31];							inform_L[32][4] = l_cell_wire[32];							inform_L[48][4] = l_cell_wire[33];							inform_L[33][4] = l_cell_wire[34];							inform_L[49][4] = l_cell_wire[35];							inform_L[34][4] = l_cell_wire[36];							inform_L[50][4] = l_cell_wire[37];							inform_L[35][4] = l_cell_wire[38];							inform_L[51][4] = l_cell_wire[39];							inform_L[36][4] = l_cell_wire[40];							inform_L[52][4] = l_cell_wire[41];							inform_L[37][4] = l_cell_wire[42];							inform_L[53][4] = l_cell_wire[43];							inform_L[38][4] = l_cell_wire[44];							inform_L[54][4] = l_cell_wire[45];							inform_L[39][4] = l_cell_wire[46];							inform_L[55][4] = l_cell_wire[47];							inform_L[40][4] = l_cell_wire[48];							inform_L[56][4] = l_cell_wire[49];							inform_L[41][4] = l_cell_wire[50];							inform_L[57][4] = l_cell_wire[51];							inform_L[42][4] = l_cell_wire[52];							inform_L[58][4] = l_cell_wire[53];							inform_L[43][4] = l_cell_wire[54];							inform_L[59][4] = l_cell_wire[55];							inform_L[44][4] = l_cell_wire[56];							inform_L[60][4] = l_cell_wire[57];							inform_L[45][4] = l_cell_wire[58];							inform_L[61][4] = l_cell_wire[59];							inform_L[46][4] = l_cell_wire[60];							inform_L[62][4] = l_cell_wire[61];							inform_L[47][4] = l_cell_wire[62];							inform_L[63][4] = l_cell_wire[63];							inform_L[64][4] = l_cell_wire[64];							inform_L[80][4] = l_cell_wire[65];							inform_L[65][4] = l_cell_wire[66];							inform_L[81][4] = l_cell_wire[67];							inform_L[66][4] = l_cell_wire[68];							inform_L[82][4] = l_cell_wire[69];							inform_L[67][4] = l_cell_wire[70];							inform_L[83][4] = l_cell_wire[71];							inform_L[68][4] = l_cell_wire[72];							inform_L[84][4] = l_cell_wire[73];							inform_L[69][4] = l_cell_wire[74];							inform_L[85][4] = l_cell_wire[75];							inform_L[70][4] = l_cell_wire[76];							inform_L[86][4] = l_cell_wire[77];							inform_L[71][4] = l_cell_wire[78];							inform_L[87][4] = l_cell_wire[79];							inform_L[72][4] = l_cell_wire[80];							inform_L[88][4] = l_cell_wire[81];							inform_L[73][4] = l_cell_wire[82];							inform_L[89][4] = l_cell_wire[83];							inform_L[74][4] = l_cell_wire[84];							inform_L[90][4] = l_cell_wire[85];							inform_L[75][4] = l_cell_wire[86];							inform_L[91][4] = l_cell_wire[87];							inform_L[76][4] = l_cell_wire[88];							inform_L[92][4] = l_cell_wire[89];							inform_L[77][4] = l_cell_wire[90];							inform_L[93][4] = l_cell_wire[91];							inform_L[78][4] = l_cell_wire[92];							inform_L[94][4] = l_cell_wire[93];							inform_L[79][4] = l_cell_wire[94];							inform_L[95][4] = l_cell_wire[95];							inform_L[96][4] = l_cell_wire[96];							inform_L[112][4] = l_cell_wire[97];							inform_L[97][4] = l_cell_wire[98];							inform_L[113][4] = l_cell_wire[99];							inform_L[98][4] = l_cell_wire[100];							inform_L[114][4] = l_cell_wire[101];							inform_L[99][4] = l_cell_wire[102];							inform_L[115][4] = l_cell_wire[103];							inform_L[100][4] = l_cell_wire[104];							inform_L[116][4] = l_cell_wire[105];							inform_L[101][4] = l_cell_wire[106];							inform_L[117][4] = l_cell_wire[107];							inform_L[102][4] = l_cell_wire[108];							inform_L[118][4] = l_cell_wire[109];							inform_L[103][4] = l_cell_wire[110];							inform_L[119][4] = l_cell_wire[111];							inform_L[104][4] = l_cell_wire[112];							inform_L[120][4] = l_cell_wire[113];							inform_L[105][4] = l_cell_wire[114];							inform_L[121][4] = l_cell_wire[115];							inform_L[106][4] = l_cell_wire[116];							inform_L[122][4] = l_cell_wire[117];							inform_L[107][4] = l_cell_wire[118];							inform_L[123][4] = l_cell_wire[119];							inform_L[108][4] = l_cell_wire[120];							inform_L[124][4] = l_cell_wire[121];							inform_L[109][4] = l_cell_wire[122];							inform_L[125][4] = l_cell_wire[123];							inform_L[110][4] = l_cell_wire[124];							inform_L[126][4] = l_cell_wire[125];							inform_L[111][4] = l_cell_wire[126];							inform_L[127][4] = l_cell_wire[127];							inform_L[128][4] = l_cell_wire[128];							inform_L[144][4] = l_cell_wire[129];							inform_L[129][4] = l_cell_wire[130];							inform_L[145][4] = l_cell_wire[131];							inform_L[130][4] = l_cell_wire[132];							inform_L[146][4] = l_cell_wire[133];							inform_L[131][4] = l_cell_wire[134];							inform_L[147][4] = l_cell_wire[135];							inform_L[132][4] = l_cell_wire[136];							inform_L[148][4] = l_cell_wire[137];							inform_L[133][4] = l_cell_wire[138];							inform_L[149][4] = l_cell_wire[139];							inform_L[134][4] = l_cell_wire[140];							inform_L[150][4] = l_cell_wire[141];							inform_L[135][4] = l_cell_wire[142];							inform_L[151][4] = l_cell_wire[143];							inform_L[136][4] = l_cell_wire[144];							inform_L[152][4] = l_cell_wire[145];							inform_L[137][4] = l_cell_wire[146];							inform_L[153][4] = l_cell_wire[147];							inform_L[138][4] = l_cell_wire[148];							inform_L[154][4] = l_cell_wire[149];							inform_L[139][4] = l_cell_wire[150];							inform_L[155][4] = l_cell_wire[151];							inform_L[140][4] = l_cell_wire[152];							inform_L[156][4] = l_cell_wire[153];							inform_L[141][4] = l_cell_wire[154];							inform_L[157][4] = l_cell_wire[155];							inform_L[142][4] = l_cell_wire[156];							inform_L[158][4] = l_cell_wire[157];							inform_L[143][4] = l_cell_wire[158];							inform_L[159][4] = l_cell_wire[159];							inform_L[160][4] = l_cell_wire[160];							inform_L[176][4] = l_cell_wire[161];							inform_L[161][4] = l_cell_wire[162];							inform_L[177][4] = l_cell_wire[163];							inform_L[162][4] = l_cell_wire[164];							inform_L[178][4] = l_cell_wire[165];							inform_L[163][4] = l_cell_wire[166];							inform_L[179][4] = l_cell_wire[167];							inform_L[164][4] = l_cell_wire[168];							inform_L[180][4] = l_cell_wire[169];							inform_L[165][4] = l_cell_wire[170];							inform_L[181][4] = l_cell_wire[171];							inform_L[166][4] = l_cell_wire[172];							inform_L[182][4] = l_cell_wire[173];							inform_L[167][4] = l_cell_wire[174];							inform_L[183][4] = l_cell_wire[175];							inform_L[168][4] = l_cell_wire[176];							inform_L[184][4] = l_cell_wire[177];							inform_L[169][4] = l_cell_wire[178];							inform_L[185][4] = l_cell_wire[179];							inform_L[170][4] = l_cell_wire[180];							inform_L[186][4] = l_cell_wire[181];							inform_L[171][4] = l_cell_wire[182];							inform_L[187][4] = l_cell_wire[183];							inform_L[172][4] = l_cell_wire[184];							inform_L[188][4] = l_cell_wire[185];							inform_L[173][4] = l_cell_wire[186];							inform_L[189][4] = l_cell_wire[187];							inform_L[174][4] = l_cell_wire[188];							inform_L[190][4] = l_cell_wire[189];							inform_L[175][4] = l_cell_wire[190];							inform_L[191][4] = l_cell_wire[191];							inform_L[192][4] = l_cell_wire[192];							inform_L[208][4] = l_cell_wire[193];							inform_L[193][4] = l_cell_wire[194];							inform_L[209][4] = l_cell_wire[195];							inform_L[194][4] = l_cell_wire[196];							inform_L[210][4] = l_cell_wire[197];							inform_L[195][4] = l_cell_wire[198];							inform_L[211][4] = l_cell_wire[199];							inform_L[196][4] = l_cell_wire[200];							inform_L[212][4] = l_cell_wire[201];							inform_L[197][4] = l_cell_wire[202];							inform_L[213][4] = l_cell_wire[203];							inform_L[198][4] = l_cell_wire[204];							inform_L[214][4] = l_cell_wire[205];							inform_L[199][4] = l_cell_wire[206];							inform_L[215][4] = l_cell_wire[207];							inform_L[200][4] = l_cell_wire[208];							inform_L[216][4] = l_cell_wire[209];							inform_L[201][4] = l_cell_wire[210];							inform_L[217][4] = l_cell_wire[211];							inform_L[202][4] = l_cell_wire[212];							inform_L[218][4] = l_cell_wire[213];							inform_L[203][4] = l_cell_wire[214];							inform_L[219][4] = l_cell_wire[215];							inform_L[204][4] = l_cell_wire[216];							inform_L[220][4] = l_cell_wire[217];							inform_L[205][4] = l_cell_wire[218];							inform_L[221][4] = l_cell_wire[219];							inform_L[206][4] = l_cell_wire[220];							inform_L[222][4] = l_cell_wire[221];							inform_L[207][4] = l_cell_wire[222];							inform_L[223][4] = l_cell_wire[223];							inform_L[224][4] = l_cell_wire[224];							inform_L[240][4] = l_cell_wire[225];							inform_L[225][4] = l_cell_wire[226];							inform_L[241][4] = l_cell_wire[227];							inform_L[226][4] = l_cell_wire[228];							inform_L[242][4] = l_cell_wire[229];							inform_L[227][4] = l_cell_wire[230];							inform_L[243][4] = l_cell_wire[231];							inform_L[228][4] = l_cell_wire[232];							inform_L[244][4] = l_cell_wire[233];							inform_L[229][4] = l_cell_wire[234];							inform_L[245][4] = l_cell_wire[235];							inform_L[230][4] = l_cell_wire[236];							inform_L[246][4] = l_cell_wire[237];							inform_L[231][4] = l_cell_wire[238];							inform_L[247][4] = l_cell_wire[239];							inform_L[232][4] = l_cell_wire[240];							inform_L[248][4] = l_cell_wire[241];							inform_L[233][4] = l_cell_wire[242];							inform_L[249][4] = l_cell_wire[243];							inform_L[234][4] = l_cell_wire[244];							inform_L[250][4] = l_cell_wire[245];							inform_L[235][4] = l_cell_wire[246];							inform_L[251][4] = l_cell_wire[247];							inform_L[236][4] = l_cell_wire[248];							inform_L[252][4] = l_cell_wire[249];							inform_L[237][4] = l_cell_wire[250];							inform_L[253][4] = l_cell_wire[251];							inform_L[238][4] = l_cell_wire[252];							inform_L[254][4] = l_cell_wire[253];							inform_L[239][4] = l_cell_wire[254];							inform_L[255][4] = l_cell_wire[255];							inform_L[256][4] = l_cell_wire[256];							inform_L[272][4] = l_cell_wire[257];							inform_L[257][4] = l_cell_wire[258];							inform_L[273][4] = l_cell_wire[259];							inform_L[258][4] = l_cell_wire[260];							inform_L[274][4] = l_cell_wire[261];							inform_L[259][4] = l_cell_wire[262];							inform_L[275][4] = l_cell_wire[263];							inform_L[260][4] = l_cell_wire[264];							inform_L[276][4] = l_cell_wire[265];							inform_L[261][4] = l_cell_wire[266];							inform_L[277][4] = l_cell_wire[267];							inform_L[262][4] = l_cell_wire[268];							inform_L[278][4] = l_cell_wire[269];							inform_L[263][4] = l_cell_wire[270];							inform_L[279][4] = l_cell_wire[271];							inform_L[264][4] = l_cell_wire[272];							inform_L[280][4] = l_cell_wire[273];							inform_L[265][4] = l_cell_wire[274];							inform_L[281][4] = l_cell_wire[275];							inform_L[266][4] = l_cell_wire[276];							inform_L[282][4] = l_cell_wire[277];							inform_L[267][4] = l_cell_wire[278];							inform_L[283][4] = l_cell_wire[279];							inform_L[268][4] = l_cell_wire[280];							inform_L[284][4] = l_cell_wire[281];							inform_L[269][4] = l_cell_wire[282];							inform_L[285][4] = l_cell_wire[283];							inform_L[270][4] = l_cell_wire[284];							inform_L[286][4] = l_cell_wire[285];							inform_L[271][4] = l_cell_wire[286];							inform_L[287][4] = l_cell_wire[287];							inform_L[288][4] = l_cell_wire[288];							inform_L[304][4] = l_cell_wire[289];							inform_L[289][4] = l_cell_wire[290];							inform_L[305][4] = l_cell_wire[291];							inform_L[290][4] = l_cell_wire[292];							inform_L[306][4] = l_cell_wire[293];							inform_L[291][4] = l_cell_wire[294];							inform_L[307][4] = l_cell_wire[295];							inform_L[292][4] = l_cell_wire[296];							inform_L[308][4] = l_cell_wire[297];							inform_L[293][4] = l_cell_wire[298];							inform_L[309][4] = l_cell_wire[299];							inform_L[294][4] = l_cell_wire[300];							inform_L[310][4] = l_cell_wire[301];							inform_L[295][4] = l_cell_wire[302];							inform_L[311][4] = l_cell_wire[303];							inform_L[296][4] = l_cell_wire[304];							inform_L[312][4] = l_cell_wire[305];							inform_L[297][4] = l_cell_wire[306];							inform_L[313][4] = l_cell_wire[307];							inform_L[298][4] = l_cell_wire[308];							inform_L[314][4] = l_cell_wire[309];							inform_L[299][4] = l_cell_wire[310];							inform_L[315][4] = l_cell_wire[311];							inform_L[300][4] = l_cell_wire[312];							inform_L[316][4] = l_cell_wire[313];							inform_L[301][4] = l_cell_wire[314];							inform_L[317][4] = l_cell_wire[315];							inform_L[302][4] = l_cell_wire[316];							inform_L[318][4] = l_cell_wire[317];							inform_L[303][4] = l_cell_wire[318];							inform_L[319][4] = l_cell_wire[319];							inform_L[320][4] = l_cell_wire[320];							inform_L[336][4] = l_cell_wire[321];							inform_L[321][4] = l_cell_wire[322];							inform_L[337][4] = l_cell_wire[323];							inform_L[322][4] = l_cell_wire[324];							inform_L[338][4] = l_cell_wire[325];							inform_L[323][4] = l_cell_wire[326];							inform_L[339][4] = l_cell_wire[327];							inform_L[324][4] = l_cell_wire[328];							inform_L[340][4] = l_cell_wire[329];							inform_L[325][4] = l_cell_wire[330];							inform_L[341][4] = l_cell_wire[331];							inform_L[326][4] = l_cell_wire[332];							inform_L[342][4] = l_cell_wire[333];							inform_L[327][4] = l_cell_wire[334];							inform_L[343][4] = l_cell_wire[335];							inform_L[328][4] = l_cell_wire[336];							inform_L[344][4] = l_cell_wire[337];							inform_L[329][4] = l_cell_wire[338];							inform_L[345][4] = l_cell_wire[339];							inform_L[330][4] = l_cell_wire[340];							inform_L[346][4] = l_cell_wire[341];							inform_L[331][4] = l_cell_wire[342];							inform_L[347][4] = l_cell_wire[343];							inform_L[332][4] = l_cell_wire[344];							inform_L[348][4] = l_cell_wire[345];							inform_L[333][4] = l_cell_wire[346];							inform_L[349][4] = l_cell_wire[347];							inform_L[334][4] = l_cell_wire[348];							inform_L[350][4] = l_cell_wire[349];							inform_L[335][4] = l_cell_wire[350];							inform_L[351][4] = l_cell_wire[351];							inform_L[352][4] = l_cell_wire[352];							inform_L[368][4] = l_cell_wire[353];							inform_L[353][4] = l_cell_wire[354];							inform_L[369][4] = l_cell_wire[355];							inform_L[354][4] = l_cell_wire[356];							inform_L[370][4] = l_cell_wire[357];							inform_L[355][4] = l_cell_wire[358];							inform_L[371][4] = l_cell_wire[359];							inform_L[356][4] = l_cell_wire[360];							inform_L[372][4] = l_cell_wire[361];							inform_L[357][4] = l_cell_wire[362];							inform_L[373][4] = l_cell_wire[363];							inform_L[358][4] = l_cell_wire[364];							inform_L[374][4] = l_cell_wire[365];							inform_L[359][4] = l_cell_wire[366];							inform_L[375][4] = l_cell_wire[367];							inform_L[360][4] = l_cell_wire[368];							inform_L[376][4] = l_cell_wire[369];							inform_L[361][4] = l_cell_wire[370];							inform_L[377][4] = l_cell_wire[371];							inform_L[362][4] = l_cell_wire[372];							inform_L[378][4] = l_cell_wire[373];							inform_L[363][4] = l_cell_wire[374];							inform_L[379][4] = l_cell_wire[375];							inform_L[364][4] = l_cell_wire[376];							inform_L[380][4] = l_cell_wire[377];							inform_L[365][4] = l_cell_wire[378];							inform_L[381][4] = l_cell_wire[379];							inform_L[366][4] = l_cell_wire[380];							inform_L[382][4] = l_cell_wire[381];							inform_L[367][4] = l_cell_wire[382];							inform_L[383][4] = l_cell_wire[383];							inform_L[384][4] = l_cell_wire[384];							inform_L[400][4] = l_cell_wire[385];							inform_L[385][4] = l_cell_wire[386];							inform_L[401][4] = l_cell_wire[387];							inform_L[386][4] = l_cell_wire[388];							inform_L[402][4] = l_cell_wire[389];							inform_L[387][4] = l_cell_wire[390];							inform_L[403][4] = l_cell_wire[391];							inform_L[388][4] = l_cell_wire[392];							inform_L[404][4] = l_cell_wire[393];							inform_L[389][4] = l_cell_wire[394];							inform_L[405][4] = l_cell_wire[395];							inform_L[390][4] = l_cell_wire[396];							inform_L[406][4] = l_cell_wire[397];							inform_L[391][4] = l_cell_wire[398];							inform_L[407][4] = l_cell_wire[399];							inform_L[392][4] = l_cell_wire[400];							inform_L[408][4] = l_cell_wire[401];							inform_L[393][4] = l_cell_wire[402];							inform_L[409][4] = l_cell_wire[403];							inform_L[394][4] = l_cell_wire[404];							inform_L[410][4] = l_cell_wire[405];							inform_L[395][4] = l_cell_wire[406];							inform_L[411][4] = l_cell_wire[407];							inform_L[396][4] = l_cell_wire[408];							inform_L[412][4] = l_cell_wire[409];							inform_L[397][4] = l_cell_wire[410];							inform_L[413][4] = l_cell_wire[411];							inform_L[398][4] = l_cell_wire[412];							inform_L[414][4] = l_cell_wire[413];							inform_L[399][4] = l_cell_wire[414];							inform_L[415][4] = l_cell_wire[415];							inform_L[416][4] = l_cell_wire[416];							inform_L[432][4] = l_cell_wire[417];							inform_L[417][4] = l_cell_wire[418];							inform_L[433][4] = l_cell_wire[419];							inform_L[418][4] = l_cell_wire[420];							inform_L[434][4] = l_cell_wire[421];							inform_L[419][4] = l_cell_wire[422];							inform_L[435][4] = l_cell_wire[423];							inform_L[420][4] = l_cell_wire[424];							inform_L[436][4] = l_cell_wire[425];							inform_L[421][4] = l_cell_wire[426];							inform_L[437][4] = l_cell_wire[427];							inform_L[422][4] = l_cell_wire[428];							inform_L[438][4] = l_cell_wire[429];							inform_L[423][4] = l_cell_wire[430];							inform_L[439][4] = l_cell_wire[431];							inform_L[424][4] = l_cell_wire[432];							inform_L[440][4] = l_cell_wire[433];							inform_L[425][4] = l_cell_wire[434];							inform_L[441][4] = l_cell_wire[435];							inform_L[426][4] = l_cell_wire[436];							inform_L[442][4] = l_cell_wire[437];							inform_L[427][4] = l_cell_wire[438];							inform_L[443][4] = l_cell_wire[439];							inform_L[428][4] = l_cell_wire[440];							inform_L[444][4] = l_cell_wire[441];							inform_L[429][4] = l_cell_wire[442];							inform_L[445][4] = l_cell_wire[443];							inform_L[430][4] = l_cell_wire[444];							inform_L[446][4] = l_cell_wire[445];							inform_L[431][4] = l_cell_wire[446];							inform_L[447][4] = l_cell_wire[447];							inform_L[448][4] = l_cell_wire[448];							inform_L[464][4] = l_cell_wire[449];							inform_L[449][4] = l_cell_wire[450];							inform_L[465][4] = l_cell_wire[451];							inform_L[450][4] = l_cell_wire[452];							inform_L[466][4] = l_cell_wire[453];							inform_L[451][4] = l_cell_wire[454];							inform_L[467][4] = l_cell_wire[455];							inform_L[452][4] = l_cell_wire[456];							inform_L[468][4] = l_cell_wire[457];							inform_L[453][4] = l_cell_wire[458];							inform_L[469][4] = l_cell_wire[459];							inform_L[454][4] = l_cell_wire[460];							inform_L[470][4] = l_cell_wire[461];							inform_L[455][4] = l_cell_wire[462];							inform_L[471][4] = l_cell_wire[463];							inform_L[456][4] = l_cell_wire[464];							inform_L[472][4] = l_cell_wire[465];							inform_L[457][4] = l_cell_wire[466];							inform_L[473][4] = l_cell_wire[467];							inform_L[458][4] = l_cell_wire[468];							inform_L[474][4] = l_cell_wire[469];							inform_L[459][4] = l_cell_wire[470];							inform_L[475][4] = l_cell_wire[471];							inform_L[460][4] = l_cell_wire[472];							inform_L[476][4] = l_cell_wire[473];							inform_L[461][4] = l_cell_wire[474];							inform_L[477][4] = l_cell_wire[475];							inform_L[462][4] = l_cell_wire[476];							inform_L[478][4] = l_cell_wire[477];							inform_L[463][4] = l_cell_wire[478];							inform_L[479][4] = l_cell_wire[479];							inform_L[480][4] = l_cell_wire[480];							inform_L[496][4] = l_cell_wire[481];							inform_L[481][4] = l_cell_wire[482];							inform_L[497][4] = l_cell_wire[483];							inform_L[482][4] = l_cell_wire[484];							inform_L[498][4] = l_cell_wire[485];							inform_L[483][4] = l_cell_wire[486];							inform_L[499][4] = l_cell_wire[487];							inform_L[484][4] = l_cell_wire[488];							inform_L[500][4] = l_cell_wire[489];							inform_L[485][4] = l_cell_wire[490];							inform_L[501][4] = l_cell_wire[491];							inform_L[486][4] = l_cell_wire[492];							inform_L[502][4] = l_cell_wire[493];							inform_L[487][4] = l_cell_wire[494];							inform_L[503][4] = l_cell_wire[495];							inform_L[488][4] = l_cell_wire[496];							inform_L[504][4] = l_cell_wire[497];							inform_L[489][4] = l_cell_wire[498];							inform_L[505][4] = l_cell_wire[499];							inform_L[490][4] = l_cell_wire[500];							inform_L[506][4] = l_cell_wire[501];							inform_L[491][4] = l_cell_wire[502];							inform_L[507][4] = l_cell_wire[503];							inform_L[492][4] = l_cell_wire[504];							inform_L[508][4] = l_cell_wire[505];							inform_L[493][4] = l_cell_wire[506];							inform_L[509][4] = l_cell_wire[507];							inform_L[494][4] = l_cell_wire[508];							inform_L[510][4] = l_cell_wire[509];							inform_L[495][4] = l_cell_wire[510];							inform_L[511][4] = l_cell_wire[511];							inform_L[512][4] = l_cell_wire[512];							inform_L[528][4] = l_cell_wire[513];							inform_L[513][4] = l_cell_wire[514];							inform_L[529][4] = l_cell_wire[515];							inform_L[514][4] = l_cell_wire[516];							inform_L[530][4] = l_cell_wire[517];							inform_L[515][4] = l_cell_wire[518];							inform_L[531][4] = l_cell_wire[519];							inform_L[516][4] = l_cell_wire[520];							inform_L[532][4] = l_cell_wire[521];							inform_L[517][4] = l_cell_wire[522];							inform_L[533][4] = l_cell_wire[523];							inform_L[518][4] = l_cell_wire[524];							inform_L[534][4] = l_cell_wire[525];							inform_L[519][4] = l_cell_wire[526];							inform_L[535][4] = l_cell_wire[527];							inform_L[520][4] = l_cell_wire[528];							inform_L[536][4] = l_cell_wire[529];							inform_L[521][4] = l_cell_wire[530];							inform_L[537][4] = l_cell_wire[531];							inform_L[522][4] = l_cell_wire[532];							inform_L[538][4] = l_cell_wire[533];							inform_L[523][4] = l_cell_wire[534];							inform_L[539][4] = l_cell_wire[535];							inform_L[524][4] = l_cell_wire[536];							inform_L[540][4] = l_cell_wire[537];							inform_L[525][4] = l_cell_wire[538];							inform_L[541][4] = l_cell_wire[539];							inform_L[526][4] = l_cell_wire[540];							inform_L[542][4] = l_cell_wire[541];							inform_L[527][4] = l_cell_wire[542];							inform_L[543][4] = l_cell_wire[543];							inform_L[544][4] = l_cell_wire[544];							inform_L[560][4] = l_cell_wire[545];							inform_L[545][4] = l_cell_wire[546];							inform_L[561][4] = l_cell_wire[547];							inform_L[546][4] = l_cell_wire[548];							inform_L[562][4] = l_cell_wire[549];							inform_L[547][4] = l_cell_wire[550];							inform_L[563][4] = l_cell_wire[551];							inform_L[548][4] = l_cell_wire[552];							inform_L[564][4] = l_cell_wire[553];							inform_L[549][4] = l_cell_wire[554];							inform_L[565][4] = l_cell_wire[555];							inform_L[550][4] = l_cell_wire[556];							inform_L[566][4] = l_cell_wire[557];							inform_L[551][4] = l_cell_wire[558];							inform_L[567][4] = l_cell_wire[559];							inform_L[552][4] = l_cell_wire[560];							inform_L[568][4] = l_cell_wire[561];							inform_L[553][4] = l_cell_wire[562];							inform_L[569][4] = l_cell_wire[563];							inform_L[554][4] = l_cell_wire[564];							inform_L[570][4] = l_cell_wire[565];							inform_L[555][4] = l_cell_wire[566];							inform_L[571][4] = l_cell_wire[567];							inform_L[556][4] = l_cell_wire[568];							inform_L[572][4] = l_cell_wire[569];							inform_L[557][4] = l_cell_wire[570];							inform_L[573][4] = l_cell_wire[571];							inform_L[558][4] = l_cell_wire[572];							inform_L[574][4] = l_cell_wire[573];							inform_L[559][4] = l_cell_wire[574];							inform_L[575][4] = l_cell_wire[575];							inform_L[576][4] = l_cell_wire[576];							inform_L[592][4] = l_cell_wire[577];							inform_L[577][4] = l_cell_wire[578];							inform_L[593][4] = l_cell_wire[579];							inform_L[578][4] = l_cell_wire[580];							inform_L[594][4] = l_cell_wire[581];							inform_L[579][4] = l_cell_wire[582];							inform_L[595][4] = l_cell_wire[583];							inform_L[580][4] = l_cell_wire[584];							inform_L[596][4] = l_cell_wire[585];							inform_L[581][4] = l_cell_wire[586];							inform_L[597][4] = l_cell_wire[587];							inform_L[582][4] = l_cell_wire[588];							inform_L[598][4] = l_cell_wire[589];							inform_L[583][4] = l_cell_wire[590];							inform_L[599][4] = l_cell_wire[591];							inform_L[584][4] = l_cell_wire[592];							inform_L[600][4] = l_cell_wire[593];							inform_L[585][4] = l_cell_wire[594];							inform_L[601][4] = l_cell_wire[595];							inform_L[586][4] = l_cell_wire[596];							inform_L[602][4] = l_cell_wire[597];							inform_L[587][4] = l_cell_wire[598];							inform_L[603][4] = l_cell_wire[599];							inform_L[588][4] = l_cell_wire[600];							inform_L[604][4] = l_cell_wire[601];							inform_L[589][4] = l_cell_wire[602];							inform_L[605][4] = l_cell_wire[603];							inform_L[590][4] = l_cell_wire[604];							inform_L[606][4] = l_cell_wire[605];							inform_L[591][4] = l_cell_wire[606];							inform_L[607][4] = l_cell_wire[607];							inform_L[608][4] = l_cell_wire[608];							inform_L[624][4] = l_cell_wire[609];							inform_L[609][4] = l_cell_wire[610];							inform_L[625][4] = l_cell_wire[611];							inform_L[610][4] = l_cell_wire[612];							inform_L[626][4] = l_cell_wire[613];							inform_L[611][4] = l_cell_wire[614];							inform_L[627][4] = l_cell_wire[615];							inform_L[612][4] = l_cell_wire[616];							inform_L[628][4] = l_cell_wire[617];							inform_L[613][4] = l_cell_wire[618];							inform_L[629][4] = l_cell_wire[619];							inform_L[614][4] = l_cell_wire[620];							inform_L[630][4] = l_cell_wire[621];							inform_L[615][4] = l_cell_wire[622];							inform_L[631][4] = l_cell_wire[623];							inform_L[616][4] = l_cell_wire[624];							inform_L[632][4] = l_cell_wire[625];							inform_L[617][4] = l_cell_wire[626];							inform_L[633][4] = l_cell_wire[627];							inform_L[618][4] = l_cell_wire[628];							inform_L[634][4] = l_cell_wire[629];							inform_L[619][4] = l_cell_wire[630];							inform_L[635][4] = l_cell_wire[631];							inform_L[620][4] = l_cell_wire[632];							inform_L[636][4] = l_cell_wire[633];							inform_L[621][4] = l_cell_wire[634];							inform_L[637][4] = l_cell_wire[635];							inform_L[622][4] = l_cell_wire[636];							inform_L[638][4] = l_cell_wire[637];							inform_L[623][4] = l_cell_wire[638];							inform_L[639][4] = l_cell_wire[639];							inform_L[640][4] = l_cell_wire[640];							inform_L[656][4] = l_cell_wire[641];							inform_L[641][4] = l_cell_wire[642];							inform_L[657][4] = l_cell_wire[643];							inform_L[642][4] = l_cell_wire[644];							inform_L[658][4] = l_cell_wire[645];							inform_L[643][4] = l_cell_wire[646];							inform_L[659][4] = l_cell_wire[647];							inform_L[644][4] = l_cell_wire[648];							inform_L[660][4] = l_cell_wire[649];							inform_L[645][4] = l_cell_wire[650];							inform_L[661][4] = l_cell_wire[651];							inform_L[646][4] = l_cell_wire[652];							inform_L[662][4] = l_cell_wire[653];							inform_L[647][4] = l_cell_wire[654];							inform_L[663][4] = l_cell_wire[655];							inform_L[648][4] = l_cell_wire[656];							inform_L[664][4] = l_cell_wire[657];							inform_L[649][4] = l_cell_wire[658];							inform_L[665][4] = l_cell_wire[659];							inform_L[650][4] = l_cell_wire[660];							inform_L[666][4] = l_cell_wire[661];							inform_L[651][4] = l_cell_wire[662];							inform_L[667][4] = l_cell_wire[663];							inform_L[652][4] = l_cell_wire[664];							inform_L[668][4] = l_cell_wire[665];							inform_L[653][4] = l_cell_wire[666];							inform_L[669][4] = l_cell_wire[667];							inform_L[654][4] = l_cell_wire[668];							inform_L[670][4] = l_cell_wire[669];							inform_L[655][4] = l_cell_wire[670];							inform_L[671][4] = l_cell_wire[671];							inform_L[672][4] = l_cell_wire[672];							inform_L[688][4] = l_cell_wire[673];							inform_L[673][4] = l_cell_wire[674];							inform_L[689][4] = l_cell_wire[675];							inform_L[674][4] = l_cell_wire[676];							inform_L[690][4] = l_cell_wire[677];							inform_L[675][4] = l_cell_wire[678];							inform_L[691][4] = l_cell_wire[679];							inform_L[676][4] = l_cell_wire[680];							inform_L[692][4] = l_cell_wire[681];							inform_L[677][4] = l_cell_wire[682];							inform_L[693][4] = l_cell_wire[683];							inform_L[678][4] = l_cell_wire[684];							inform_L[694][4] = l_cell_wire[685];							inform_L[679][4] = l_cell_wire[686];							inform_L[695][4] = l_cell_wire[687];							inform_L[680][4] = l_cell_wire[688];							inform_L[696][4] = l_cell_wire[689];							inform_L[681][4] = l_cell_wire[690];							inform_L[697][4] = l_cell_wire[691];							inform_L[682][4] = l_cell_wire[692];							inform_L[698][4] = l_cell_wire[693];							inform_L[683][4] = l_cell_wire[694];							inform_L[699][4] = l_cell_wire[695];							inform_L[684][4] = l_cell_wire[696];							inform_L[700][4] = l_cell_wire[697];							inform_L[685][4] = l_cell_wire[698];							inform_L[701][4] = l_cell_wire[699];							inform_L[686][4] = l_cell_wire[700];							inform_L[702][4] = l_cell_wire[701];							inform_L[687][4] = l_cell_wire[702];							inform_L[703][4] = l_cell_wire[703];							inform_L[704][4] = l_cell_wire[704];							inform_L[720][4] = l_cell_wire[705];							inform_L[705][4] = l_cell_wire[706];							inform_L[721][4] = l_cell_wire[707];							inform_L[706][4] = l_cell_wire[708];							inform_L[722][4] = l_cell_wire[709];							inform_L[707][4] = l_cell_wire[710];							inform_L[723][4] = l_cell_wire[711];							inform_L[708][4] = l_cell_wire[712];							inform_L[724][4] = l_cell_wire[713];							inform_L[709][4] = l_cell_wire[714];							inform_L[725][4] = l_cell_wire[715];							inform_L[710][4] = l_cell_wire[716];							inform_L[726][4] = l_cell_wire[717];							inform_L[711][4] = l_cell_wire[718];							inform_L[727][4] = l_cell_wire[719];							inform_L[712][4] = l_cell_wire[720];							inform_L[728][4] = l_cell_wire[721];							inform_L[713][4] = l_cell_wire[722];							inform_L[729][4] = l_cell_wire[723];							inform_L[714][4] = l_cell_wire[724];							inform_L[730][4] = l_cell_wire[725];							inform_L[715][4] = l_cell_wire[726];							inform_L[731][4] = l_cell_wire[727];							inform_L[716][4] = l_cell_wire[728];							inform_L[732][4] = l_cell_wire[729];							inform_L[717][4] = l_cell_wire[730];							inform_L[733][4] = l_cell_wire[731];							inform_L[718][4] = l_cell_wire[732];							inform_L[734][4] = l_cell_wire[733];							inform_L[719][4] = l_cell_wire[734];							inform_L[735][4] = l_cell_wire[735];							inform_L[736][4] = l_cell_wire[736];							inform_L[752][4] = l_cell_wire[737];							inform_L[737][4] = l_cell_wire[738];							inform_L[753][4] = l_cell_wire[739];							inform_L[738][4] = l_cell_wire[740];							inform_L[754][4] = l_cell_wire[741];							inform_L[739][4] = l_cell_wire[742];							inform_L[755][4] = l_cell_wire[743];							inform_L[740][4] = l_cell_wire[744];							inform_L[756][4] = l_cell_wire[745];							inform_L[741][4] = l_cell_wire[746];							inform_L[757][4] = l_cell_wire[747];							inform_L[742][4] = l_cell_wire[748];							inform_L[758][4] = l_cell_wire[749];							inform_L[743][4] = l_cell_wire[750];							inform_L[759][4] = l_cell_wire[751];							inform_L[744][4] = l_cell_wire[752];							inform_L[760][4] = l_cell_wire[753];							inform_L[745][4] = l_cell_wire[754];							inform_L[761][4] = l_cell_wire[755];							inform_L[746][4] = l_cell_wire[756];							inform_L[762][4] = l_cell_wire[757];							inform_L[747][4] = l_cell_wire[758];							inform_L[763][4] = l_cell_wire[759];							inform_L[748][4] = l_cell_wire[760];							inform_L[764][4] = l_cell_wire[761];							inform_L[749][4] = l_cell_wire[762];							inform_L[765][4] = l_cell_wire[763];							inform_L[750][4] = l_cell_wire[764];							inform_L[766][4] = l_cell_wire[765];							inform_L[751][4] = l_cell_wire[766];							inform_L[767][4] = l_cell_wire[767];							inform_L[768][4] = l_cell_wire[768];							inform_L[784][4] = l_cell_wire[769];							inform_L[769][4] = l_cell_wire[770];							inform_L[785][4] = l_cell_wire[771];							inform_L[770][4] = l_cell_wire[772];							inform_L[786][4] = l_cell_wire[773];							inform_L[771][4] = l_cell_wire[774];							inform_L[787][4] = l_cell_wire[775];							inform_L[772][4] = l_cell_wire[776];							inform_L[788][4] = l_cell_wire[777];							inform_L[773][4] = l_cell_wire[778];							inform_L[789][4] = l_cell_wire[779];							inform_L[774][4] = l_cell_wire[780];							inform_L[790][4] = l_cell_wire[781];							inform_L[775][4] = l_cell_wire[782];							inform_L[791][4] = l_cell_wire[783];							inform_L[776][4] = l_cell_wire[784];							inform_L[792][4] = l_cell_wire[785];							inform_L[777][4] = l_cell_wire[786];							inform_L[793][4] = l_cell_wire[787];							inform_L[778][4] = l_cell_wire[788];							inform_L[794][4] = l_cell_wire[789];							inform_L[779][4] = l_cell_wire[790];							inform_L[795][4] = l_cell_wire[791];							inform_L[780][4] = l_cell_wire[792];							inform_L[796][4] = l_cell_wire[793];							inform_L[781][4] = l_cell_wire[794];							inform_L[797][4] = l_cell_wire[795];							inform_L[782][4] = l_cell_wire[796];							inform_L[798][4] = l_cell_wire[797];							inform_L[783][4] = l_cell_wire[798];							inform_L[799][4] = l_cell_wire[799];							inform_L[800][4] = l_cell_wire[800];							inform_L[816][4] = l_cell_wire[801];							inform_L[801][4] = l_cell_wire[802];							inform_L[817][4] = l_cell_wire[803];							inform_L[802][4] = l_cell_wire[804];							inform_L[818][4] = l_cell_wire[805];							inform_L[803][4] = l_cell_wire[806];							inform_L[819][4] = l_cell_wire[807];							inform_L[804][4] = l_cell_wire[808];							inform_L[820][4] = l_cell_wire[809];							inform_L[805][4] = l_cell_wire[810];							inform_L[821][4] = l_cell_wire[811];							inform_L[806][4] = l_cell_wire[812];							inform_L[822][4] = l_cell_wire[813];							inform_L[807][4] = l_cell_wire[814];							inform_L[823][4] = l_cell_wire[815];							inform_L[808][4] = l_cell_wire[816];							inform_L[824][4] = l_cell_wire[817];							inform_L[809][4] = l_cell_wire[818];							inform_L[825][4] = l_cell_wire[819];							inform_L[810][4] = l_cell_wire[820];							inform_L[826][4] = l_cell_wire[821];							inform_L[811][4] = l_cell_wire[822];							inform_L[827][4] = l_cell_wire[823];							inform_L[812][4] = l_cell_wire[824];							inform_L[828][4] = l_cell_wire[825];							inform_L[813][4] = l_cell_wire[826];							inform_L[829][4] = l_cell_wire[827];							inform_L[814][4] = l_cell_wire[828];							inform_L[830][4] = l_cell_wire[829];							inform_L[815][4] = l_cell_wire[830];							inform_L[831][4] = l_cell_wire[831];							inform_L[832][4] = l_cell_wire[832];							inform_L[848][4] = l_cell_wire[833];							inform_L[833][4] = l_cell_wire[834];							inform_L[849][4] = l_cell_wire[835];							inform_L[834][4] = l_cell_wire[836];							inform_L[850][4] = l_cell_wire[837];							inform_L[835][4] = l_cell_wire[838];							inform_L[851][4] = l_cell_wire[839];							inform_L[836][4] = l_cell_wire[840];							inform_L[852][4] = l_cell_wire[841];							inform_L[837][4] = l_cell_wire[842];							inform_L[853][4] = l_cell_wire[843];							inform_L[838][4] = l_cell_wire[844];							inform_L[854][4] = l_cell_wire[845];							inform_L[839][4] = l_cell_wire[846];							inform_L[855][4] = l_cell_wire[847];							inform_L[840][4] = l_cell_wire[848];							inform_L[856][4] = l_cell_wire[849];							inform_L[841][4] = l_cell_wire[850];							inform_L[857][4] = l_cell_wire[851];							inform_L[842][4] = l_cell_wire[852];							inform_L[858][4] = l_cell_wire[853];							inform_L[843][4] = l_cell_wire[854];							inform_L[859][4] = l_cell_wire[855];							inform_L[844][4] = l_cell_wire[856];							inform_L[860][4] = l_cell_wire[857];							inform_L[845][4] = l_cell_wire[858];							inform_L[861][4] = l_cell_wire[859];							inform_L[846][4] = l_cell_wire[860];							inform_L[862][4] = l_cell_wire[861];							inform_L[847][4] = l_cell_wire[862];							inform_L[863][4] = l_cell_wire[863];							inform_L[864][4] = l_cell_wire[864];							inform_L[880][4] = l_cell_wire[865];							inform_L[865][4] = l_cell_wire[866];							inform_L[881][4] = l_cell_wire[867];							inform_L[866][4] = l_cell_wire[868];							inform_L[882][4] = l_cell_wire[869];							inform_L[867][4] = l_cell_wire[870];							inform_L[883][4] = l_cell_wire[871];							inform_L[868][4] = l_cell_wire[872];							inform_L[884][4] = l_cell_wire[873];							inform_L[869][4] = l_cell_wire[874];							inform_L[885][4] = l_cell_wire[875];							inform_L[870][4] = l_cell_wire[876];							inform_L[886][4] = l_cell_wire[877];							inform_L[871][4] = l_cell_wire[878];							inform_L[887][4] = l_cell_wire[879];							inform_L[872][4] = l_cell_wire[880];							inform_L[888][4] = l_cell_wire[881];							inform_L[873][4] = l_cell_wire[882];							inform_L[889][4] = l_cell_wire[883];							inform_L[874][4] = l_cell_wire[884];							inform_L[890][4] = l_cell_wire[885];							inform_L[875][4] = l_cell_wire[886];							inform_L[891][4] = l_cell_wire[887];							inform_L[876][4] = l_cell_wire[888];							inform_L[892][4] = l_cell_wire[889];							inform_L[877][4] = l_cell_wire[890];							inform_L[893][4] = l_cell_wire[891];							inform_L[878][4] = l_cell_wire[892];							inform_L[894][4] = l_cell_wire[893];							inform_L[879][4] = l_cell_wire[894];							inform_L[895][4] = l_cell_wire[895];							inform_L[896][4] = l_cell_wire[896];							inform_L[912][4] = l_cell_wire[897];							inform_L[897][4] = l_cell_wire[898];							inform_L[913][4] = l_cell_wire[899];							inform_L[898][4] = l_cell_wire[900];							inform_L[914][4] = l_cell_wire[901];							inform_L[899][4] = l_cell_wire[902];							inform_L[915][4] = l_cell_wire[903];							inform_L[900][4] = l_cell_wire[904];							inform_L[916][4] = l_cell_wire[905];							inform_L[901][4] = l_cell_wire[906];							inform_L[917][4] = l_cell_wire[907];							inform_L[902][4] = l_cell_wire[908];							inform_L[918][4] = l_cell_wire[909];							inform_L[903][4] = l_cell_wire[910];							inform_L[919][4] = l_cell_wire[911];							inform_L[904][4] = l_cell_wire[912];							inform_L[920][4] = l_cell_wire[913];							inform_L[905][4] = l_cell_wire[914];							inform_L[921][4] = l_cell_wire[915];							inform_L[906][4] = l_cell_wire[916];							inform_L[922][4] = l_cell_wire[917];							inform_L[907][4] = l_cell_wire[918];							inform_L[923][4] = l_cell_wire[919];							inform_L[908][4] = l_cell_wire[920];							inform_L[924][4] = l_cell_wire[921];							inform_L[909][4] = l_cell_wire[922];							inform_L[925][4] = l_cell_wire[923];							inform_L[910][4] = l_cell_wire[924];							inform_L[926][4] = l_cell_wire[925];							inform_L[911][4] = l_cell_wire[926];							inform_L[927][4] = l_cell_wire[927];							inform_L[928][4] = l_cell_wire[928];							inform_L[944][4] = l_cell_wire[929];							inform_L[929][4] = l_cell_wire[930];							inform_L[945][4] = l_cell_wire[931];							inform_L[930][4] = l_cell_wire[932];							inform_L[946][4] = l_cell_wire[933];							inform_L[931][4] = l_cell_wire[934];							inform_L[947][4] = l_cell_wire[935];							inform_L[932][4] = l_cell_wire[936];							inform_L[948][4] = l_cell_wire[937];							inform_L[933][4] = l_cell_wire[938];							inform_L[949][4] = l_cell_wire[939];							inform_L[934][4] = l_cell_wire[940];							inform_L[950][4] = l_cell_wire[941];							inform_L[935][4] = l_cell_wire[942];							inform_L[951][4] = l_cell_wire[943];							inform_L[936][4] = l_cell_wire[944];							inform_L[952][4] = l_cell_wire[945];							inform_L[937][4] = l_cell_wire[946];							inform_L[953][4] = l_cell_wire[947];							inform_L[938][4] = l_cell_wire[948];							inform_L[954][4] = l_cell_wire[949];							inform_L[939][4] = l_cell_wire[950];							inform_L[955][4] = l_cell_wire[951];							inform_L[940][4] = l_cell_wire[952];							inform_L[956][4] = l_cell_wire[953];							inform_L[941][4] = l_cell_wire[954];							inform_L[957][4] = l_cell_wire[955];							inform_L[942][4] = l_cell_wire[956];							inform_L[958][4] = l_cell_wire[957];							inform_L[943][4] = l_cell_wire[958];							inform_L[959][4] = l_cell_wire[959];							inform_L[960][4] = l_cell_wire[960];							inform_L[976][4] = l_cell_wire[961];							inform_L[961][4] = l_cell_wire[962];							inform_L[977][4] = l_cell_wire[963];							inform_L[962][4] = l_cell_wire[964];							inform_L[978][4] = l_cell_wire[965];							inform_L[963][4] = l_cell_wire[966];							inform_L[979][4] = l_cell_wire[967];							inform_L[964][4] = l_cell_wire[968];							inform_L[980][4] = l_cell_wire[969];							inform_L[965][4] = l_cell_wire[970];							inform_L[981][4] = l_cell_wire[971];							inform_L[966][4] = l_cell_wire[972];							inform_L[982][4] = l_cell_wire[973];							inform_L[967][4] = l_cell_wire[974];							inform_L[983][4] = l_cell_wire[975];							inform_L[968][4] = l_cell_wire[976];							inform_L[984][4] = l_cell_wire[977];							inform_L[969][4] = l_cell_wire[978];							inform_L[985][4] = l_cell_wire[979];							inform_L[970][4] = l_cell_wire[980];							inform_L[986][4] = l_cell_wire[981];							inform_L[971][4] = l_cell_wire[982];							inform_L[987][4] = l_cell_wire[983];							inform_L[972][4] = l_cell_wire[984];							inform_L[988][4] = l_cell_wire[985];							inform_L[973][4] = l_cell_wire[986];							inform_L[989][4] = l_cell_wire[987];							inform_L[974][4] = l_cell_wire[988];							inform_L[990][4] = l_cell_wire[989];							inform_L[975][4] = l_cell_wire[990];							inform_L[991][4] = l_cell_wire[991];							inform_L[992][4] = l_cell_wire[992];							inform_L[1008][4] = l_cell_wire[993];							inform_L[993][4] = l_cell_wire[994];							inform_L[1009][4] = l_cell_wire[995];							inform_L[994][4] = l_cell_wire[996];							inform_L[1010][4] = l_cell_wire[997];							inform_L[995][4] = l_cell_wire[998];							inform_L[1011][4] = l_cell_wire[999];							inform_L[996][4] = l_cell_wire[1000];							inform_L[1012][4] = l_cell_wire[1001];							inform_L[997][4] = l_cell_wire[1002];							inform_L[1013][4] = l_cell_wire[1003];							inform_L[998][4] = l_cell_wire[1004];							inform_L[1014][4] = l_cell_wire[1005];							inform_L[999][4] = l_cell_wire[1006];							inform_L[1015][4] = l_cell_wire[1007];							inform_L[1000][4] = l_cell_wire[1008];							inform_L[1016][4] = l_cell_wire[1009];							inform_L[1001][4] = l_cell_wire[1010];							inform_L[1017][4] = l_cell_wire[1011];							inform_L[1002][4] = l_cell_wire[1012];							inform_L[1018][4] = l_cell_wire[1013];							inform_L[1003][4] = l_cell_wire[1014];							inform_L[1019][4] = l_cell_wire[1015];							inform_L[1004][4] = l_cell_wire[1016];							inform_L[1020][4] = l_cell_wire[1017];							inform_L[1005][4] = l_cell_wire[1018];							inform_L[1021][4] = l_cell_wire[1019];							inform_L[1006][4] = l_cell_wire[1020];							inform_L[1022][4] = l_cell_wire[1021];							inform_L[1007][4] = l_cell_wire[1022];							inform_L[1023][4] = l_cell_wire[1023];						end
						6:						begin							inform_R[0][6] = r_cell_wire[0];							inform_R[32][6] = r_cell_wire[1];							inform_R[1][6] = r_cell_wire[2];							inform_R[33][6] = r_cell_wire[3];							inform_R[2][6] = r_cell_wire[4];							inform_R[34][6] = r_cell_wire[5];							inform_R[3][6] = r_cell_wire[6];							inform_R[35][6] = r_cell_wire[7];							inform_R[4][6] = r_cell_wire[8];							inform_R[36][6] = r_cell_wire[9];							inform_R[5][6] = r_cell_wire[10];							inform_R[37][6] = r_cell_wire[11];							inform_R[6][6] = r_cell_wire[12];							inform_R[38][6] = r_cell_wire[13];							inform_R[7][6] = r_cell_wire[14];							inform_R[39][6] = r_cell_wire[15];							inform_R[8][6] = r_cell_wire[16];							inform_R[40][6] = r_cell_wire[17];							inform_R[9][6] = r_cell_wire[18];							inform_R[41][6] = r_cell_wire[19];							inform_R[10][6] = r_cell_wire[20];							inform_R[42][6] = r_cell_wire[21];							inform_R[11][6] = r_cell_wire[22];							inform_R[43][6] = r_cell_wire[23];							inform_R[12][6] = r_cell_wire[24];							inform_R[44][6] = r_cell_wire[25];							inform_R[13][6] = r_cell_wire[26];							inform_R[45][6] = r_cell_wire[27];							inform_R[14][6] = r_cell_wire[28];							inform_R[46][6] = r_cell_wire[29];							inform_R[15][6] = r_cell_wire[30];							inform_R[47][6] = r_cell_wire[31];							inform_R[16][6] = r_cell_wire[32];							inform_R[48][6] = r_cell_wire[33];							inform_R[17][6] = r_cell_wire[34];							inform_R[49][6] = r_cell_wire[35];							inform_R[18][6] = r_cell_wire[36];							inform_R[50][6] = r_cell_wire[37];							inform_R[19][6] = r_cell_wire[38];							inform_R[51][6] = r_cell_wire[39];							inform_R[20][6] = r_cell_wire[40];							inform_R[52][6] = r_cell_wire[41];							inform_R[21][6] = r_cell_wire[42];							inform_R[53][6] = r_cell_wire[43];							inform_R[22][6] = r_cell_wire[44];							inform_R[54][6] = r_cell_wire[45];							inform_R[23][6] = r_cell_wire[46];							inform_R[55][6] = r_cell_wire[47];							inform_R[24][6] = r_cell_wire[48];							inform_R[56][6] = r_cell_wire[49];							inform_R[25][6] = r_cell_wire[50];							inform_R[57][6] = r_cell_wire[51];							inform_R[26][6] = r_cell_wire[52];							inform_R[58][6] = r_cell_wire[53];							inform_R[27][6] = r_cell_wire[54];							inform_R[59][6] = r_cell_wire[55];							inform_R[28][6] = r_cell_wire[56];							inform_R[60][6] = r_cell_wire[57];							inform_R[29][6] = r_cell_wire[58];							inform_R[61][6] = r_cell_wire[59];							inform_R[30][6] = r_cell_wire[60];							inform_R[62][6] = r_cell_wire[61];							inform_R[31][6] = r_cell_wire[62];							inform_R[63][6] = r_cell_wire[63];							inform_R[64][6] = r_cell_wire[64];							inform_R[96][6] = r_cell_wire[65];							inform_R[65][6] = r_cell_wire[66];							inform_R[97][6] = r_cell_wire[67];							inform_R[66][6] = r_cell_wire[68];							inform_R[98][6] = r_cell_wire[69];							inform_R[67][6] = r_cell_wire[70];							inform_R[99][6] = r_cell_wire[71];							inform_R[68][6] = r_cell_wire[72];							inform_R[100][6] = r_cell_wire[73];							inform_R[69][6] = r_cell_wire[74];							inform_R[101][6] = r_cell_wire[75];							inform_R[70][6] = r_cell_wire[76];							inform_R[102][6] = r_cell_wire[77];							inform_R[71][6] = r_cell_wire[78];							inform_R[103][6] = r_cell_wire[79];							inform_R[72][6] = r_cell_wire[80];							inform_R[104][6] = r_cell_wire[81];							inform_R[73][6] = r_cell_wire[82];							inform_R[105][6] = r_cell_wire[83];							inform_R[74][6] = r_cell_wire[84];							inform_R[106][6] = r_cell_wire[85];							inform_R[75][6] = r_cell_wire[86];							inform_R[107][6] = r_cell_wire[87];							inform_R[76][6] = r_cell_wire[88];							inform_R[108][6] = r_cell_wire[89];							inform_R[77][6] = r_cell_wire[90];							inform_R[109][6] = r_cell_wire[91];							inform_R[78][6] = r_cell_wire[92];							inform_R[110][6] = r_cell_wire[93];							inform_R[79][6] = r_cell_wire[94];							inform_R[111][6] = r_cell_wire[95];							inform_R[80][6] = r_cell_wire[96];							inform_R[112][6] = r_cell_wire[97];							inform_R[81][6] = r_cell_wire[98];							inform_R[113][6] = r_cell_wire[99];							inform_R[82][6] = r_cell_wire[100];							inform_R[114][6] = r_cell_wire[101];							inform_R[83][6] = r_cell_wire[102];							inform_R[115][6] = r_cell_wire[103];							inform_R[84][6] = r_cell_wire[104];							inform_R[116][6] = r_cell_wire[105];							inform_R[85][6] = r_cell_wire[106];							inform_R[117][6] = r_cell_wire[107];							inform_R[86][6] = r_cell_wire[108];							inform_R[118][6] = r_cell_wire[109];							inform_R[87][6] = r_cell_wire[110];							inform_R[119][6] = r_cell_wire[111];							inform_R[88][6] = r_cell_wire[112];							inform_R[120][6] = r_cell_wire[113];							inform_R[89][6] = r_cell_wire[114];							inform_R[121][6] = r_cell_wire[115];							inform_R[90][6] = r_cell_wire[116];							inform_R[122][6] = r_cell_wire[117];							inform_R[91][6] = r_cell_wire[118];							inform_R[123][6] = r_cell_wire[119];							inform_R[92][6] = r_cell_wire[120];							inform_R[124][6] = r_cell_wire[121];							inform_R[93][6] = r_cell_wire[122];							inform_R[125][6] = r_cell_wire[123];							inform_R[94][6] = r_cell_wire[124];							inform_R[126][6] = r_cell_wire[125];							inform_R[95][6] = r_cell_wire[126];							inform_R[127][6] = r_cell_wire[127];							inform_R[128][6] = r_cell_wire[128];							inform_R[160][6] = r_cell_wire[129];							inform_R[129][6] = r_cell_wire[130];							inform_R[161][6] = r_cell_wire[131];							inform_R[130][6] = r_cell_wire[132];							inform_R[162][6] = r_cell_wire[133];							inform_R[131][6] = r_cell_wire[134];							inform_R[163][6] = r_cell_wire[135];							inform_R[132][6] = r_cell_wire[136];							inform_R[164][6] = r_cell_wire[137];							inform_R[133][6] = r_cell_wire[138];							inform_R[165][6] = r_cell_wire[139];							inform_R[134][6] = r_cell_wire[140];							inform_R[166][6] = r_cell_wire[141];							inform_R[135][6] = r_cell_wire[142];							inform_R[167][6] = r_cell_wire[143];							inform_R[136][6] = r_cell_wire[144];							inform_R[168][6] = r_cell_wire[145];							inform_R[137][6] = r_cell_wire[146];							inform_R[169][6] = r_cell_wire[147];							inform_R[138][6] = r_cell_wire[148];							inform_R[170][6] = r_cell_wire[149];							inform_R[139][6] = r_cell_wire[150];							inform_R[171][6] = r_cell_wire[151];							inform_R[140][6] = r_cell_wire[152];							inform_R[172][6] = r_cell_wire[153];							inform_R[141][6] = r_cell_wire[154];							inform_R[173][6] = r_cell_wire[155];							inform_R[142][6] = r_cell_wire[156];							inform_R[174][6] = r_cell_wire[157];							inform_R[143][6] = r_cell_wire[158];							inform_R[175][6] = r_cell_wire[159];							inform_R[144][6] = r_cell_wire[160];							inform_R[176][6] = r_cell_wire[161];							inform_R[145][6] = r_cell_wire[162];							inform_R[177][6] = r_cell_wire[163];							inform_R[146][6] = r_cell_wire[164];							inform_R[178][6] = r_cell_wire[165];							inform_R[147][6] = r_cell_wire[166];							inform_R[179][6] = r_cell_wire[167];							inform_R[148][6] = r_cell_wire[168];							inform_R[180][6] = r_cell_wire[169];							inform_R[149][6] = r_cell_wire[170];							inform_R[181][6] = r_cell_wire[171];							inform_R[150][6] = r_cell_wire[172];							inform_R[182][6] = r_cell_wire[173];							inform_R[151][6] = r_cell_wire[174];							inform_R[183][6] = r_cell_wire[175];							inform_R[152][6] = r_cell_wire[176];							inform_R[184][6] = r_cell_wire[177];							inform_R[153][6] = r_cell_wire[178];							inform_R[185][6] = r_cell_wire[179];							inform_R[154][6] = r_cell_wire[180];							inform_R[186][6] = r_cell_wire[181];							inform_R[155][6] = r_cell_wire[182];							inform_R[187][6] = r_cell_wire[183];							inform_R[156][6] = r_cell_wire[184];							inform_R[188][6] = r_cell_wire[185];							inform_R[157][6] = r_cell_wire[186];							inform_R[189][6] = r_cell_wire[187];							inform_R[158][6] = r_cell_wire[188];							inform_R[190][6] = r_cell_wire[189];							inform_R[159][6] = r_cell_wire[190];							inform_R[191][6] = r_cell_wire[191];							inform_R[192][6] = r_cell_wire[192];							inform_R[224][6] = r_cell_wire[193];							inform_R[193][6] = r_cell_wire[194];							inform_R[225][6] = r_cell_wire[195];							inform_R[194][6] = r_cell_wire[196];							inform_R[226][6] = r_cell_wire[197];							inform_R[195][6] = r_cell_wire[198];							inform_R[227][6] = r_cell_wire[199];							inform_R[196][6] = r_cell_wire[200];							inform_R[228][6] = r_cell_wire[201];							inform_R[197][6] = r_cell_wire[202];							inform_R[229][6] = r_cell_wire[203];							inform_R[198][6] = r_cell_wire[204];							inform_R[230][6] = r_cell_wire[205];							inform_R[199][6] = r_cell_wire[206];							inform_R[231][6] = r_cell_wire[207];							inform_R[200][6] = r_cell_wire[208];							inform_R[232][6] = r_cell_wire[209];							inform_R[201][6] = r_cell_wire[210];							inform_R[233][6] = r_cell_wire[211];							inform_R[202][6] = r_cell_wire[212];							inform_R[234][6] = r_cell_wire[213];							inform_R[203][6] = r_cell_wire[214];							inform_R[235][6] = r_cell_wire[215];							inform_R[204][6] = r_cell_wire[216];							inform_R[236][6] = r_cell_wire[217];							inform_R[205][6] = r_cell_wire[218];							inform_R[237][6] = r_cell_wire[219];							inform_R[206][6] = r_cell_wire[220];							inform_R[238][6] = r_cell_wire[221];							inform_R[207][6] = r_cell_wire[222];							inform_R[239][6] = r_cell_wire[223];							inform_R[208][6] = r_cell_wire[224];							inform_R[240][6] = r_cell_wire[225];							inform_R[209][6] = r_cell_wire[226];							inform_R[241][6] = r_cell_wire[227];							inform_R[210][6] = r_cell_wire[228];							inform_R[242][6] = r_cell_wire[229];							inform_R[211][6] = r_cell_wire[230];							inform_R[243][6] = r_cell_wire[231];							inform_R[212][6] = r_cell_wire[232];							inform_R[244][6] = r_cell_wire[233];							inform_R[213][6] = r_cell_wire[234];							inform_R[245][6] = r_cell_wire[235];							inform_R[214][6] = r_cell_wire[236];							inform_R[246][6] = r_cell_wire[237];							inform_R[215][6] = r_cell_wire[238];							inform_R[247][6] = r_cell_wire[239];							inform_R[216][6] = r_cell_wire[240];							inform_R[248][6] = r_cell_wire[241];							inform_R[217][6] = r_cell_wire[242];							inform_R[249][6] = r_cell_wire[243];							inform_R[218][6] = r_cell_wire[244];							inform_R[250][6] = r_cell_wire[245];							inform_R[219][6] = r_cell_wire[246];							inform_R[251][6] = r_cell_wire[247];							inform_R[220][6] = r_cell_wire[248];							inform_R[252][6] = r_cell_wire[249];							inform_R[221][6] = r_cell_wire[250];							inform_R[253][6] = r_cell_wire[251];							inform_R[222][6] = r_cell_wire[252];							inform_R[254][6] = r_cell_wire[253];							inform_R[223][6] = r_cell_wire[254];							inform_R[255][6] = r_cell_wire[255];							inform_R[256][6] = r_cell_wire[256];							inform_R[288][6] = r_cell_wire[257];							inform_R[257][6] = r_cell_wire[258];							inform_R[289][6] = r_cell_wire[259];							inform_R[258][6] = r_cell_wire[260];							inform_R[290][6] = r_cell_wire[261];							inform_R[259][6] = r_cell_wire[262];							inform_R[291][6] = r_cell_wire[263];							inform_R[260][6] = r_cell_wire[264];							inform_R[292][6] = r_cell_wire[265];							inform_R[261][6] = r_cell_wire[266];							inform_R[293][6] = r_cell_wire[267];							inform_R[262][6] = r_cell_wire[268];							inform_R[294][6] = r_cell_wire[269];							inform_R[263][6] = r_cell_wire[270];							inform_R[295][6] = r_cell_wire[271];							inform_R[264][6] = r_cell_wire[272];							inform_R[296][6] = r_cell_wire[273];							inform_R[265][6] = r_cell_wire[274];							inform_R[297][6] = r_cell_wire[275];							inform_R[266][6] = r_cell_wire[276];							inform_R[298][6] = r_cell_wire[277];							inform_R[267][6] = r_cell_wire[278];							inform_R[299][6] = r_cell_wire[279];							inform_R[268][6] = r_cell_wire[280];							inform_R[300][6] = r_cell_wire[281];							inform_R[269][6] = r_cell_wire[282];							inform_R[301][6] = r_cell_wire[283];							inform_R[270][6] = r_cell_wire[284];							inform_R[302][6] = r_cell_wire[285];							inform_R[271][6] = r_cell_wire[286];							inform_R[303][6] = r_cell_wire[287];							inform_R[272][6] = r_cell_wire[288];							inform_R[304][6] = r_cell_wire[289];							inform_R[273][6] = r_cell_wire[290];							inform_R[305][6] = r_cell_wire[291];							inform_R[274][6] = r_cell_wire[292];							inform_R[306][6] = r_cell_wire[293];							inform_R[275][6] = r_cell_wire[294];							inform_R[307][6] = r_cell_wire[295];							inform_R[276][6] = r_cell_wire[296];							inform_R[308][6] = r_cell_wire[297];							inform_R[277][6] = r_cell_wire[298];							inform_R[309][6] = r_cell_wire[299];							inform_R[278][6] = r_cell_wire[300];							inform_R[310][6] = r_cell_wire[301];							inform_R[279][6] = r_cell_wire[302];							inform_R[311][6] = r_cell_wire[303];							inform_R[280][6] = r_cell_wire[304];							inform_R[312][6] = r_cell_wire[305];							inform_R[281][6] = r_cell_wire[306];							inform_R[313][6] = r_cell_wire[307];							inform_R[282][6] = r_cell_wire[308];							inform_R[314][6] = r_cell_wire[309];							inform_R[283][6] = r_cell_wire[310];							inform_R[315][6] = r_cell_wire[311];							inform_R[284][6] = r_cell_wire[312];							inform_R[316][6] = r_cell_wire[313];							inform_R[285][6] = r_cell_wire[314];							inform_R[317][6] = r_cell_wire[315];							inform_R[286][6] = r_cell_wire[316];							inform_R[318][6] = r_cell_wire[317];							inform_R[287][6] = r_cell_wire[318];							inform_R[319][6] = r_cell_wire[319];							inform_R[320][6] = r_cell_wire[320];							inform_R[352][6] = r_cell_wire[321];							inform_R[321][6] = r_cell_wire[322];							inform_R[353][6] = r_cell_wire[323];							inform_R[322][6] = r_cell_wire[324];							inform_R[354][6] = r_cell_wire[325];							inform_R[323][6] = r_cell_wire[326];							inform_R[355][6] = r_cell_wire[327];							inform_R[324][6] = r_cell_wire[328];							inform_R[356][6] = r_cell_wire[329];							inform_R[325][6] = r_cell_wire[330];							inform_R[357][6] = r_cell_wire[331];							inform_R[326][6] = r_cell_wire[332];							inform_R[358][6] = r_cell_wire[333];							inform_R[327][6] = r_cell_wire[334];							inform_R[359][6] = r_cell_wire[335];							inform_R[328][6] = r_cell_wire[336];							inform_R[360][6] = r_cell_wire[337];							inform_R[329][6] = r_cell_wire[338];							inform_R[361][6] = r_cell_wire[339];							inform_R[330][6] = r_cell_wire[340];							inform_R[362][6] = r_cell_wire[341];							inform_R[331][6] = r_cell_wire[342];							inform_R[363][6] = r_cell_wire[343];							inform_R[332][6] = r_cell_wire[344];							inform_R[364][6] = r_cell_wire[345];							inform_R[333][6] = r_cell_wire[346];							inform_R[365][6] = r_cell_wire[347];							inform_R[334][6] = r_cell_wire[348];							inform_R[366][6] = r_cell_wire[349];							inform_R[335][6] = r_cell_wire[350];							inform_R[367][6] = r_cell_wire[351];							inform_R[336][6] = r_cell_wire[352];							inform_R[368][6] = r_cell_wire[353];							inform_R[337][6] = r_cell_wire[354];							inform_R[369][6] = r_cell_wire[355];							inform_R[338][6] = r_cell_wire[356];							inform_R[370][6] = r_cell_wire[357];							inform_R[339][6] = r_cell_wire[358];							inform_R[371][6] = r_cell_wire[359];							inform_R[340][6] = r_cell_wire[360];							inform_R[372][6] = r_cell_wire[361];							inform_R[341][6] = r_cell_wire[362];							inform_R[373][6] = r_cell_wire[363];							inform_R[342][6] = r_cell_wire[364];							inform_R[374][6] = r_cell_wire[365];							inform_R[343][6] = r_cell_wire[366];							inform_R[375][6] = r_cell_wire[367];							inform_R[344][6] = r_cell_wire[368];							inform_R[376][6] = r_cell_wire[369];							inform_R[345][6] = r_cell_wire[370];							inform_R[377][6] = r_cell_wire[371];							inform_R[346][6] = r_cell_wire[372];							inform_R[378][6] = r_cell_wire[373];							inform_R[347][6] = r_cell_wire[374];							inform_R[379][6] = r_cell_wire[375];							inform_R[348][6] = r_cell_wire[376];							inform_R[380][6] = r_cell_wire[377];							inform_R[349][6] = r_cell_wire[378];							inform_R[381][6] = r_cell_wire[379];							inform_R[350][6] = r_cell_wire[380];							inform_R[382][6] = r_cell_wire[381];							inform_R[351][6] = r_cell_wire[382];							inform_R[383][6] = r_cell_wire[383];							inform_R[384][6] = r_cell_wire[384];							inform_R[416][6] = r_cell_wire[385];							inform_R[385][6] = r_cell_wire[386];							inform_R[417][6] = r_cell_wire[387];							inform_R[386][6] = r_cell_wire[388];							inform_R[418][6] = r_cell_wire[389];							inform_R[387][6] = r_cell_wire[390];							inform_R[419][6] = r_cell_wire[391];							inform_R[388][6] = r_cell_wire[392];							inform_R[420][6] = r_cell_wire[393];							inform_R[389][6] = r_cell_wire[394];							inform_R[421][6] = r_cell_wire[395];							inform_R[390][6] = r_cell_wire[396];							inform_R[422][6] = r_cell_wire[397];							inform_R[391][6] = r_cell_wire[398];							inform_R[423][6] = r_cell_wire[399];							inform_R[392][6] = r_cell_wire[400];							inform_R[424][6] = r_cell_wire[401];							inform_R[393][6] = r_cell_wire[402];							inform_R[425][6] = r_cell_wire[403];							inform_R[394][6] = r_cell_wire[404];							inform_R[426][6] = r_cell_wire[405];							inform_R[395][6] = r_cell_wire[406];							inform_R[427][6] = r_cell_wire[407];							inform_R[396][6] = r_cell_wire[408];							inform_R[428][6] = r_cell_wire[409];							inform_R[397][6] = r_cell_wire[410];							inform_R[429][6] = r_cell_wire[411];							inform_R[398][6] = r_cell_wire[412];							inform_R[430][6] = r_cell_wire[413];							inform_R[399][6] = r_cell_wire[414];							inform_R[431][6] = r_cell_wire[415];							inform_R[400][6] = r_cell_wire[416];							inform_R[432][6] = r_cell_wire[417];							inform_R[401][6] = r_cell_wire[418];							inform_R[433][6] = r_cell_wire[419];							inform_R[402][6] = r_cell_wire[420];							inform_R[434][6] = r_cell_wire[421];							inform_R[403][6] = r_cell_wire[422];							inform_R[435][6] = r_cell_wire[423];							inform_R[404][6] = r_cell_wire[424];							inform_R[436][6] = r_cell_wire[425];							inform_R[405][6] = r_cell_wire[426];							inform_R[437][6] = r_cell_wire[427];							inform_R[406][6] = r_cell_wire[428];							inform_R[438][6] = r_cell_wire[429];							inform_R[407][6] = r_cell_wire[430];							inform_R[439][6] = r_cell_wire[431];							inform_R[408][6] = r_cell_wire[432];							inform_R[440][6] = r_cell_wire[433];							inform_R[409][6] = r_cell_wire[434];							inform_R[441][6] = r_cell_wire[435];							inform_R[410][6] = r_cell_wire[436];							inform_R[442][6] = r_cell_wire[437];							inform_R[411][6] = r_cell_wire[438];							inform_R[443][6] = r_cell_wire[439];							inform_R[412][6] = r_cell_wire[440];							inform_R[444][6] = r_cell_wire[441];							inform_R[413][6] = r_cell_wire[442];							inform_R[445][6] = r_cell_wire[443];							inform_R[414][6] = r_cell_wire[444];							inform_R[446][6] = r_cell_wire[445];							inform_R[415][6] = r_cell_wire[446];							inform_R[447][6] = r_cell_wire[447];							inform_R[448][6] = r_cell_wire[448];							inform_R[480][6] = r_cell_wire[449];							inform_R[449][6] = r_cell_wire[450];							inform_R[481][6] = r_cell_wire[451];							inform_R[450][6] = r_cell_wire[452];							inform_R[482][6] = r_cell_wire[453];							inform_R[451][6] = r_cell_wire[454];							inform_R[483][6] = r_cell_wire[455];							inform_R[452][6] = r_cell_wire[456];							inform_R[484][6] = r_cell_wire[457];							inform_R[453][6] = r_cell_wire[458];							inform_R[485][6] = r_cell_wire[459];							inform_R[454][6] = r_cell_wire[460];							inform_R[486][6] = r_cell_wire[461];							inform_R[455][6] = r_cell_wire[462];							inform_R[487][6] = r_cell_wire[463];							inform_R[456][6] = r_cell_wire[464];							inform_R[488][6] = r_cell_wire[465];							inform_R[457][6] = r_cell_wire[466];							inform_R[489][6] = r_cell_wire[467];							inform_R[458][6] = r_cell_wire[468];							inform_R[490][6] = r_cell_wire[469];							inform_R[459][6] = r_cell_wire[470];							inform_R[491][6] = r_cell_wire[471];							inform_R[460][6] = r_cell_wire[472];							inform_R[492][6] = r_cell_wire[473];							inform_R[461][6] = r_cell_wire[474];							inform_R[493][6] = r_cell_wire[475];							inform_R[462][6] = r_cell_wire[476];							inform_R[494][6] = r_cell_wire[477];							inform_R[463][6] = r_cell_wire[478];							inform_R[495][6] = r_cell_wire[479];							inform_R[464][6] = r_cell_wire[480];							inform_R[496][6] = r_cell_wire[481];							inform_R[465][6] = r_cell_wire[482];							inform_R[497][6] = r_cell_wire[483];							inform_R[466][6] = r_cell_wire[484];							inform_R[498][6] = r_cell_wire[485];							inform_R[467][6] = r_cell_wire[486];							inform_R[499][6] = r_cell_wire[487];							inform_R[468][6] = r_cell_wire[488];							inform_R[500][6] = r_cell_wire[489];							inform_R[469][6] = r_cell_wire[490];							inform_R[501][6] = r_cell_wire[491];							inform_R[470][6] = r_cell_wire[492];							inform_R[502][6] = r_cell_wire[493];							inform_R[471][6] = r_cell_wire[494];							inform_R[503][6] = r_cell_wire[495];							inform_R[472][6] = r_cell_wire[496];							inform_R[504][6] = r_cell_wire[497];							inform_R[473][6] = r_cell_wire[498];							inform_R[505][6] = r_cell_wire[499];							inform_R[474][6] = r_cell_wire[500];							inform_R[506][6] = r_cell_wire[501];							inform_R[475][6] = r_cell_wire[502];							inform_R[507][6] = r_cell_wire[503];							inform_R[476][6] = r_cell_wire[504];							inform_R[508][6] = r_cell_wire[505];							inform_R[477][6] = r_cell_wire[506];							inform_R[509][6] = r_cell_wire[507];							inform_R[478][6] = r_cell_wire[508];							inform_R[510][6] = r_cell_wire[509];							inform_R[479][6] = r_cell_wire[510];							inform_R[511][6] = r_cell_wire[511];							inform_R[512][6] = r_cell_wire[512];							inform_R[544][6] = r_cell_wire[513];							inform_R[513][6] = r_cell_wire[514];							inform_R[545][6] = r_cell_wire[515];							inform_R[514][6] = r_cell_wire[516];							inform_R[546][6] = r_cell_wire[517];							inform_R[515][6] = r_cell_wire[518];							inform_R[547][6] = r_cell_wire[519];							inform_R[516][6] = r_cell_wire[520];							inform_R[548][6] = r_cell_wire[521];							inform_R[517][6] = r_cell_wire[522];							inform_R[549][6] = r_cell_wire[523];							inform_R[518][6] = r_cell_wire[524];							inform_R[550][6] = r_cell_wire[525];							inform_R[519][6] = r_cell_wire[526];							inform_R[551][6] = r_cell_wire[527];							inform_R[520][6] = r_cell_wire[528];							inform_R[552][6] = r_cell_wire[529];							inform_R[521][6] = r_cell_wire[530];							inform_R[553][6] = r_cell_wire[531];							inform_R[522][6] = r_cell_wire[532];							inform_R[554][6] = r_cell_wire[533];							inform_R[523][6] = r_cell_wire[534];							inform_R[555][6] = r_cell_wire[535];							inform_R[524][6] = r_cell_wire[536];							inform_R[556][6] = r_cell_wire[537];							inform_R[525][6] = r_cell_wire[538];							inform_R[557][6] = r_cell_wire[539];							inform_R[526][6] = r_cell_wire[540];							inform_R[558][6] = r_cell_wire[541];							inform_R[527][6] = r_cell_wire[542];							inform_R[559][6] = r_cell_wire[543];							inform_R[528][6] = r_cell_wire[544];							inform_R[560][6] = r_cell_wire[545];							inform_R[529][6] = r_cell_wire[546];							inform_R[561][6] = r_cell_wire[547];							inform_R[530][6] = r_cell_wire[548];							inform_R[562][6] = r_cell_wire[549];							inform_R[531][6] = r_cell_wire[550];							inform_R[563][6] = r_cell_wire[551];							inform_R[532][6] = r_cell_wire[552];							inform_R[564][6] = r_cell_wire[553];							inform_R[533][6] = r_cell_wire[554];							inform_R[565][6] = r_cell_wire[555];							inform_R[534][6] = r_cell_wire[556];							inform_R[566][6] = r_cell_wire[557];							inform_R[535][6] = r_cell_wire[558];							inform_R[567][6] = r_cell_wire[559];							inform_R[536][6] = r_cell_wire[560];							inform_R[568][6] = r_cell_wire[561];							inform_R[537][6] = r_cell_wire[562];							inform_R[569][6] = r_cell_wire[563];							inform_R[538][6] = r_cell_wire[564];							inform_R[570][6] = r_cell_wire[565];							inform_R[539][6] = r_cell_wire[566];							inform_R[571][6] = r_cell_wire[567];							inform_R[540][6] = r_cell_wire[568];							inform_R[572][6] = r_cell_wire[569];							inform_R[541][6] = r_cell_wire[570];							inform_R[573][6] = r_cell_wire[571];							inform_R[542][6] = r_cell_wire[572];							inform_R[574][6] = r_cell_wire[573];							inform_R[543][6] = r_cell_wire[574];							inform_R[575][6] = r_cell_wire[575];							inform_R[576][6] = r_cell_wire[576];							inform_R[608][6] = r_cell_wire[577];							inform_R[577][6] = r_cell_wire[578];							inform_R[609][6] = r_cell_wire[579];							inform_R[578][6] = r_cell_wire[580];							inform_R[610][6] = r_cell_wire[581];							inform_R[579][6] = r_cell_wire[582];							inform_R[611][6] = r_cell_wire[583];							inform_R[580][6] = r_cell_wire[584];							inform_R[612][6] = r_cell_wire[585];							inform_R[581][6] = r_cell_wire[586];							inform_R[613][6] = r_cell_wire[587];							inform_R[582][6] = r_cell_wire[588];							inform_R[614][6] = r_cell_wire[589];							inform_R[583][6] = r_cell_wire[590];							inform_R[615][6] = r_cell_wire[591];							inform_R[584][6] = r_cell_wire[592];							inform_R[616][6] = r_cell_wire[593];							inform_R[585][6] = r_cell_wire[594];							inform_R[617][6] = r_cell_wire[595];							inform_R[586][6] = r_cell_wire[596];							inform_R[618][6] = r_cell_wire[597];							inform_R[587][6] = r_cell_wire[598];							inform_R[619][6] = r_cell_wire[599];							inform_R[588][6] = r_cell_wire[600];							inform_R[620][6] = r_cell_wire[601];							inform_R[589][6] = r_cell_wire[602];							inform_R[621][6] = r_cell_wire[603];							inform_R[590][6] = r_cell_wire[604];							inform_R[622][6] = r_cell_wire[605];							inform_R[591][6] = r_cell_wire[606];							inform_R[623][6] = r_cell_wire[607];							inform_R[592][6] = r_cell_wire[608];							inform_R[624][6] = r_cell_wire[609];							inform_R[593][6] = r_cell_wire[610];							inform_R[625][6] = r_cell_wire[611];							inform_R[594][6] = r_cell_wire[612];							inform_R[626][6] = r_cell_wire[613];							inform_R[595][6] = r_cell_wire[614];							inform_R[627][6] = r_cell_wire[615];							inform_R[596][6] = r_cell_wire[616];							inform_R[628][6] = r_cell_wire[617];							inform_R[597][6] = r_cell_wire[618];							inform_R[629][6] = r_cell_wire[619];							inform_R[598][6] = r_cell_wire[620];							inform_R[630][6] = r_cell_wire[621];							inform_R[599][6] = r_cell_wire[622];							inform_R[631][6] = r_cell_wire[623];							inform_R[600][6] = r_cell_wire[624];							inform_R[632][6] = r_cell_wire[625];							inform_R[601][6] = r_cell_wire[626];							inform_R[633][6] = r_cell_wire[627];							inform_R[602][6] = r_cell_wire[628];							inform_R[634][6] = r_cell_wire[629];							inform_R[603][6] = r_cell_wire[630];							inform_R[635][6] = r_cell_wire[631];							inform_R[604][6] = r_cell_wire[632];							inform_R[636][6] = r_cell_wire[633];							inform_R[605][6] = r_cell_wire[634];							inform_R[637][6] = r_cell_wire[635];							inform_R[606][6] = r_cell_wire[636];							inform_R[638][6] = r_cell_wire[637];							inform_R[607][6] = r_cell_wire[638];							inform_R[639][6] = r_cell_wire[639];							inform_R[640][6] = r_cell_wire[640];							inform_R[672][6] = r_cell_wire[641];							inform_R[641][6] = r_cell_wire[642];							inform_R[673][6] = r_cell_wire[643];							inform_R[642][6] = r_cell_wire[644];							inform_R[674][6] = r_cell_wire[645];							inform_R[643][6] = r_cell_wire[646];							inform_R[675][6] = r_cell_wire[647];							inform_R[644][6] = r_cell_wire[648];							inform_R[676][6] = r_cell_wire[649];							inform_R[645][6] = r_cell_wire[650];							inform_R[677][6] = r_cell_wire[651];							inform_R[646][6] = r_cell_wire[652];							inform_R[678][6] = r_cell_wire[653];							inform_R[647][6] = r_cell_wire[654];							inform_R[679][6] = r_cell_wire[655];							inform_R[648][6] = r_cell_wire[656];							inform_R[680][6] = r_cell_wire[657];							inform_R[649][6] = r_cell_wire[658];							inform_R[681][6] = r_cell_wire[659];							inform_R[650][6] = r_cell_wire[660];							inform_R[682][6] = r_cell_wire[661];							inform_R[651][6] = r_cell_wire[662];							inform_R[683][6] = r_cell_wire[663];							inform_R[652][6] = r_cell_wire[664];							inform_R[684][6] = r_cell_wire[665];							inform_R[653][6] = r_cell_wire[666];							inform_R[685][6] = r_cell_wire[667];							inform_R[654][6] = r_cell_wire[668];							inform_R[686][6] = r_cell_wire[669];							inform_R[655][6] = r_cell_wire[670];							inform_R[687][6] = r_cell_wire[671];							inform_R[656][6] = r_cell_wire[672];							inform_R[688][6] = r_cell_wire[673];							inform_R[657][6] = r_cell_wire[674];							inform_R[689][6] = r_cell_wire[675];							inform_R[658][6] = r_cell_wire[676];							inform_R[690][6] = r_cell_wire[677];							inform_R[659][6] = r_cell_wire[678];							inform_R[691][6] = r_cell_wire[679];							inform_R[660][6] = r_cell_wire[680];							inform_R[692][6] = r_cell_wire[681];							inform_R[661][6] = r_cell_wire[682];							inform_R[693][6] = r_cell_wire[683];							inform_R[662][6] = r_cell_wire[684];							inform_R[694][6] = r_cell_wire[685];							inform_R[663][6] = r_cell_wire[686];							inform_R[695][6] = r_cell_wire[687];							inform_R[664][6] = r_cell_wire[688];							inform_R[696][6] = r_cell_wire[689];							inform_R[665][6] = r_cell_wire[690];							inform_R[697][6] = r_cell_wire[691];							inform_R[666][6] = r_cell_wire[692];							inform_R[698][6] = r_cell_wire[693];							inform_R[667][6] = r_cell_wire[694];							inform_R[699][6] = r_cell_wire[695];							inform_R[668][6] = r_cell_wire[696];							inform_R[700][6] = r_cell_wire[697];							inform_R[669][6] = r_cell_wire[698];							inform_R[701][6] = r_cell_wire[699];							inform_R[670][6] = r_cell_wire[700];							inform_R[702][6] = r_cell_wire[701];							inform_R[671][6] = r_cell_wire[702];							inform_R[703][6] = r_cell_wire[703];							inform_R[704][6] = r_cell_wire[704];							inform_R[736][6] = r_cell_wire[705];							inform_R[705][6] = r_cell_wire[706];							inform_R[737][6] = r_cell_wire[707];							inform_R[706][6] = r_cell_wire[708];							inform_R[738][6] = r_cell_wire[709];							inform_R[707][6] = r_cell_wire[710];							inform_R[739][6] = r_cell_wire[711];							inform_R[708][6] = r_cell_wire[712];							inform_R[740][6] = r_cell_wire[713];							inform_R[709][6] = r_cell_wire[714];							inform_R[741][6] = r_cell_wire[715];							inform_R[710][6] = r_cell_wire[716];							inform_R[742][6] = r_cell_wire[717];							inform_R[711][6] = r_cell_wire[718];							inform_R[743][6] = r_cell_wire[719];							inform_R[712][6] = r_cell_wire[720];							inform_R[744][6] = r_cell_wire[721];							inform_R[713][6] = r_cell_wire[722];							inform_R[745][6] = r_cell_wire[723];							inform_R[714][6] = r_cell_wire[724];							inform_R[746][6] = r_cell_wire[725];							inform_R[715][6] = r_cell_wire[726];							inform_R[747][6] = r_cell_wire[727];							inform_R[716][6] = r_cell_wire[728];							inform_R[748][6] = r_cell_wire[729];							inform_R[717][6] = r_cell_wire[730];							inform_R[749][6] = r_cell_wire[731];							inform_R[718][6] = r_cell_wire[732];							inform_R[750][6] = r_cell_wire[733];							inform_R[719][6] = r_cell_wire[734];							inform_R[751][6] = r_cell_wire[735];							inform_R[720][6] = r_cell_wire[736];							inform_R[752][6] = r_cell_wire[737];							inform_R[721][6] = r_cell_wire[738];							inform_R[753][6] = r_cell_wire[739];							inform_R[722][6] = r_cell_wire[740];							inform_R[754][6] = r_cell_wire[741];							inform_R[723][6] = r_cell_wire[742];							inform_R[755][6] = r_cell_wire[743];							inform_R[724][6] = r_cell_wire[744];							inform_R[756][6] = r_cell_wire[745];							inform_R[725][6] = r_cell_wire[746];							inform_R[757][6] = r_cell_wire[747];							inform_R[726][6] = r_cell_wire[748];							inform_R[758][6] = r_cell_wire[749];							inform_R[727][6] = r_cell_wire[750];							inform_R[759][6] = r_cell_wire[751];							inform_R[728][6] = r_cell_wire[752];							inform_R[760][6] = r_cell_wire[753];							inform_R[729][6] = r_cell_wire[754];							inform_R[761][6] = r_cell_wire[755];							inform_R[730][6] = r_cell_wire[756];							inform_R[762][6] = r_cell_wire[757];							inform_R[731][6] = r_cell_wire[758];							inform_R[763][6] = r_cell_wire[759];							inform_R[732][6] = r_cell_wire[760];							inform_R[764][6] = r_cell_wire[761];							inform_R[733][6] = r_cell_wire[762];							inform_R[765][6] = r_cell_wire[763];							inform_R[734][6] = r_cell_wire[764];							inform_R[766][6] = r_cell_wire[765];							inform_R[735][6] = r_cell_wire[766];							inform_R[767][6] = r_cell_wire[767];							inform_R[768][6] = r_cell_wire[768];							inform_R[800][6] = r_cell_wire[769];							inform_R[769][6] = r_cell_wire[770];							inform_R[801][6] = r_cell_wire[771];							inform_R[770][6] = r_cell_wire[772];							inform_R[802][6] = r_cell_wire[773];							inform_R[771][6] = r_cell_wire[774];							inform_R[803][6] = r_cell_wire[775];							inform_R[772][6] = r_cell_wire[776];							inform_R[804][6] = r_cell_wire[777];							inform_R[773][6] = r_cell_wire[778];							inform_R[805][6] = r_cell_wire[779];							inform_R[774][6] = r_cell_wire[780];							inform_R[806][6] = r_cell_wire[781];							inform_R[775][6] = r_cell_wire[782];							inform_R[807][6] = r_cell_wire[783];							inform_R[776][6] = r_cell_wire[784];							inform_R[808][6] = r_cell_wire[785];							inform_R[777][6] = r_cell_wire[786];							inform_R[809][6] = r_cell_wire[787];							inform_R[778][6] = r_cell_wire[788];							inform_R[810][6] = r_cell_wire[789];							inform_R[779][6] = r_cell_wire[790];							inform_R[811][6] = r_cell_wire[791];							inform_R[780][6] = r_cell_wire[792];							inform_R[812][6] = r_cell_wire[793];							inform_R[781][6] = r_cell_wire[794];							inform_R[813][6] = r_cell_wire[795];							inform_R[782][6] = r_cell_wire[796];							inform_R[814][6] = r_cell_wire[797];							inform_R[783][6] = r_cell_wire[798];							inform_R[815][6] = r_cell_wire[799];							inform_R[784][6] = r_cell_wire[800];							inform_R[816][6] = r_cell_wire[801];							inform_R[785][6] = r_cell_wire[802];							inform_R[817][6] = r_cell_wire[803];							inform_R[786][6] = r_cell_wire[804];							inform_R[818][6] = r_cell_wire[805];							inform_R[787][6] = r_cell_wire[806];							inform_R[819][6] = r_cell_wire[807];							inform_R[788][6] = r_cell_wire[808];							inform_R[820][6] = r_cell_wire[809];							inform_R[789][6] = r_cell_wire[810];							inform_R[821][6] = r_cell_wire[811];							inform_R[790][6] = r_cell_wire[812];							inform_R[822][6] = r_cell_wire[813];							inform_R[791][6] = r_cell_wire[814];							inform_R[823][6] = r_cell_wire[815];							inform_R[792][6] = r_cell_wire[816];							inform_R[824][6] = r_cell_wire[817];							inform_R[793][6] = r_cell_wire[818];							inform_R[825][6] = r_cell_wire[819];							inform_R[794][6] = r_cell_wire[820];							inform_R[826][6] = r_cell_wire[821];							inform_R[795][6] = r_cell_wire[822];							inform_R[827][6] = r_cell_wire[823];							inform_R[796][6] = r_cell_wire[824];							inform_R[828][6] = r_cell_wire[825];							inform_R[797][6] = r_cell_wire[826];							inform_R[829][6] = r_cell_wire[827];							inform_R[798][6] = r_cell_wire[828];							inform_R[830][6] = r_cell_wire[829];							inform_R[799][6] = r_cell_wire[830];							inform_R[831][6] = r_cell_wire[831];							inform_R[832][6] = r_cell_wire[832];							inform_R[864][6] = r_cell_wire[833];							inform_R[833][6] = r_cell_wire[834];							inform_R[865][6] = r_cell_wire[835];							inform_R[834][6] = r_cell_wire[836];							inform_R[866][6] = r_cell_wire[837];							inform_R[835][6] = r_cell_wire[838];							inform_R[867][6] = r_cell_wire[839];							inform_R[836][6] = r_cell_wire[840];							inform_R[868][6] = r_cell_wire[841];							inform_R[837][6] = r_cell_wire[842];							inform_R[869][6] = r_cell_wire[843];							inform_R[838][6] = r_cell_wire[844];							inform_R[870][6] = r_cell_wire[845];							inform_R[839][6] = r_cell_wire[846];							inform_R[871][6] = r_cell_wire[847];							inform_R[840][6] = r_cell_wire[848];							inform_R[872][6] = r_cell_wire[849];							inform_R[841][6] = r_cell_wire[850];							inform_R[873][6] = r_cell_wire[851];							inform_R[842][6] = r_cell_wire[852];							inform_R[874][6] = r_cell_wire[853];							inform_R[843][6] = r_cell_wire[854];							inform_R[875][6] = r_cell_wire[855];							inform_R[844][6] = r_cell_wire[856];							inform_R[876][6] = r_cell_wire[857];							inform_R[845][6] = r_cell_wire[858];							inform_R[877][6] = r_cell_wire[859];							inform_R[846][6] = r_cell_wire[860];							inform_R[878][6] = r_cell_wire[861];							inform_R[847][6] = r_cell_wire[862];							inform_R[879][6] = r_cell_wire[863];							inform_R[848][6] = r_cell_wire[864];							inform_R[880][6] = r_cell_wire[865];							inform_R[849][6] = r_cell_wire[866];							inform_R[881][6] = r_cell_wire[867];							inform_R[850][6] = r_cell_wire[868];							inform_R[882][6] = r_cell_wire[869];							inform_R[851][6] = r_cell_wire[870];							inform_R[883][6] = r_cell_wire[871];							inform_R[852][6] = r_cell_wire[872];							inform_R[884][6] = r_cell_wire[873];							inform_R[853][6] = r_cell_wire[874];							inform_R[885][6] = r_cell_wire[875];							inform_R[854][6] = r_cell_wire[876];							inform_R[886][6] = r_cell_wire[877];							inform_R[855][6] = r_cell_wire[878];							inform_R[887][6] = r_cell_wire[879];							inform_R[856][6] = r_cell_wire[880];							inform_R[888][6] = r_cell_wire[881];							inform_R[857][6] = r_cell_wire[882];							inform_R[889][6] = r_cell_wire[883];							inform_R[858][6] = r_cell_wire[884];							inform_R[890][6] = r_cell_wire[885];							inform_R[859][6] = r_cell_wire[886];							inform_R[891][6] = r_cell_wire[887];							inform_R[860][6] = r_cell_wire[888];							inform_R[892][6] = r_cell_wire[889];							inform_R[861][6] = r_cell_wire[890];							inform_R[893][6] = r_cell_wire[891];							inform_R[862][6] = r_cell_wire[892];							inform_R[894][6] = r_cell_wire[893];							inform_R[863][6] = r_cell_wire[894];							inform_R[895][6] = r_cell_wire[895];							inform_R[896][6] = r_cell_wire[896];							inform_R[928][6] = r_cell_wire[897];							inform_R[897][6] = r_cell_wire[898];							inform_R[929][6] = r_cell_wire[899];							inform_R[898][6] = r_cell_wire[900];							inform_R[930][6] = r_cell_wire[901];							inform_R[899][6] = r_cell_wire[902];							inform_R[931][6] = r_cell_wire[903];							inform_R[900][6] = r_cell_wire[904];							inform_R[932][6] = r_cell_wire[905];							inform_R[901][6] = r_cell_wire[906];							inform_R[933][6] = r_cell_wire[907];							inform_R[902][6] = r_cell_wire[908];							inform_R[934][6] = r_cell_wire[909];							inform_R[903][6] = r_cell_wire[910];							inform_R[935][6] = r_cell_wire[911];							inform_R[904][6] = r_cell_wire[912];							inform_R[936][6] = r_cell_wire[913];							inform_R[905][6] = r_cell_wire[914];							inform_R[937][6] = r_cell_wire[915];							inform_R[906][6] = r_cell_wire[916];							inform_R[938][6] = r_cell_wire[917];							inform_R[907][6] = r_cell_wire[918];							inform_R[939][6] = r_cell_wire[919];							inform_R[908][6] = r_cell_wire[920];							inform_R[940][6] = r_cell_wire[921];							inform_R[909][6] = r_cell_wire[922];							inform_R[941][6] = r_cell_wire[923];							inform_R[910][6] = r_cell_wire[924];							inform_R[942][6] = r_cell_wire[925];							inform_R[911][6] = r_cell_wire[926];							inform_R[943][6] = r_cell_wire[927];							inform_R[912][6] = r_cell_wire[928];							inform_R[944][6] = r_cell_wire[929];							inform_R[913][6] = r_cell_wire[930];							inform_R[945][6] = r_cell_wire[931];							inform_R[914][6] = r_cell_wire[932];							inform_R[946][6] = r_cell_wire[933];							inform_R[915][6] = r_cell_wire[934];							inform_R[947][6] = r_cell_wire[935];							inform_R[916][6] = r_cell_wire[936];							inform_R[948][6] = r_cell_wire[937];							inform_R[917][6] = r_cell_wire[938];							inform_R[949][6] = r_cell_wire[939];							inform_R[918][6] = r_cell_wire[940];							inform_R[950][6] = r_cell_wire[941];							inform_R[919][6] = r_cell_wire[942];							inform_R[951][6] = r_cell_wire[943];							inform_R[920][6] = r_cell_wire[944];							inform_R[952][6] = r_cell_wire[945];							inform_R[921][6] = r_cell_wire[946];							inform_R[953][6] = r_cell_wire[947];							inform_R[922][6] = r_cell_wire[948];							inform_R[954][6] = r_cell_wire[949];							inform_R[923][6] = r_cell_wire[950];							inform_R[955][6] = r_cell_wire[951];							inform_R[924][6] = r_cell_wire[952];							inform_R[956][6] = r_cell_wire[953];							inform_R[925][6] = r_cell_wire[954];							inform_R[957][6] = r_cell_wire[955];							inform_R[926][6] = r_cell_wire[956];							inform_R[958][6] = r_cell_wire[957];							inform_R[927][6] = r_cell_wire[958];							inform_R[959][6] = r_cell_wire[959];							inform_R[960][6] = r_cell_wire[960];							inform_R[992][6] = r_cell_wire[961];							inform_R[961][6] = r_cell_wire[962];							inform_R[993][6] = r_cell_wire[963];							inform_R[962][6] = r_cell_wire[964];							inform_R[994][6] = r_cell_wire[965];							inform_R[963][6] = r_cell_wire[966];							inform_R[995][6] = r_cell_wire[967];							inform_R[964][6] = r_cell_wire[968];							inform_R[996][6] = r_cell_wire[969];							inform_R[965][6] = r_cell_wire[970];							inform_R[997][6] = r_cell_wire[971];							inform_R[966][6] = r_cell_wire[972];							inform_R[998][6] = r_cell_wire[973];							inform_R[967][6] = r_cell_wire[974];							inform_R[999][6] = r_cell_wire[975];							inform_R[968][6] = r_cell_wire[976];							inform_R[1000][6] = r_cell_wire[977];							inform_R[969][6] = r_cell_wire[978];							inform_R[1001][6] = r_cell_wire[979];							inform_R[970][6] = r_cell_wire[980];							inform_R[1002][6] = r_cell_wire[981];							inform_R[971][6] = r_cell_wire[982];							inform_R[1003][6] = r_cell_wire[983];							inform_R[972][6] = r_cell_wire[984];							inform_R[1004][6] = r_cell_wire[985];							inform_R[973][6] = r_cell_wire[986];							inform_R[1005][6] = r_cell_wire[987];							inform_R[974][6] = r_cell_wire[988];							inform_R[1006][6] = r_cell_wire[989];							inform_R[975][6] = r_cell_wire[990];							inform_R[1007][6] = r_cell_wire[991];							inform_R[976][6] = r_cell_wire[992];							inform_R[1008][6] = r_cell_wire[993];							inform_R[977][6] = r_cell_wire[994];							inform_R[1009][6] = r_cell_wire[995];							inform_R[978][6] = r_cell_wire[996];							inform_R[1010][6] = r_cell_wire[997];							inform_R[979][6] = r_cell_wire[998];							inform_R[1011][6] = r_cell_wire[999];							inform_R[980][6] = r_cell_wire[1000];							inform_R[1012][6] = r_cell_wire[1001];							inform_R[981][6] = r_cell_wire[1002];							inform_R[1013][6] = r_cell_wire[1003];							inform_R[982][6] = r_cell_wire[1004];							inform_R[1014][6] = r_cell_wire[1005];							inform_R[983][6] = r_cell_wire[1006];							inform_R[1015][6] = r_cell_wire[1007];							inform_R[984][6] = r_cell_wire[1008];							inform_R[1016][6] = r_cell_wire[1009];							inform_R[985][6] = r_cell_wire[1010];							inform_R[1017][6] = r_cell_wire[1011];							inform_R[986][6] = r_cell_wire[1012];							inform_R[1018][6] = r_cell_wire[1013];							inform_R[987][6] = r_cell_wire[1014];							inform_R[1019][6] = r_cell_wire[1015];							inform_R[988][6] = r_cell_wire[1016];							inform_R[1020][6] = r_cell_wire[1017];							inform_R[989][6] = r_cell_wire[1018];							inform_R[1021][6] = r_cell_wire[1019];							inform_R[990][6] = r_cell_wire[1020];							inform_R[1022][6] = r_cell_wire[1021];							inform_R[991][6] = r_cell_wire[1022];							inform_R[1023][6] = r_cell_wire[1023];							inform_L[0][5] = l_cell_wire[0];							inform_L[32][5] = l_cell_wire[1];							inform_L[1][5] = l_cell_wire[2];							inform_L[33][5] = l_cell_wire[3];							inform_L[2][5] = l_cell_wire[4];							inform_L[34][5] = l_cell_wire[5];							inform_L[3][5] = l_cell_wire[6];							inform_L[35][5] = l_cell_wire[7];							inform_L[4][5] = l_cell_wire[8];							inform_L[36][5] = l_cell_wire[9];							inform_L[5][5] = l_cell_wire[10];							inform_L[37][5] = l_cell_wire[11];							inform_L[6][5] = l_cell_wire[12];							inform_L[38][5] = l_cell_wire[13];							inform_L[7][5] = l_cell_wire[14];							inform_L[39][5] = l_cell_wire[15];							inform_L[8][5] = l_cell_wire[16];							inform_L[40][5] = l_cell_wire[17];							inform_L[9][5] = l_cell_wire[18];							inform_L[41][5] = l_cell_wire[19];							inform_L[10][5] = l_cell_wire[20];							inform_L[42][5] = l_cell_wire[21];							inform_L[11][5] = l_cell_wire[22];							inform_L[43][5] = l_cell_wire[23];							inform_L[12][5] = l_cell_wire[24];							inform_L[44][5] = l_cell_wire[25];							inform_L[13][5] = l_cell_wire[26];							inform_L[45][5] = l_cell_wire[27];							inform_L[14][5] = l_cell_wire[28];							inform_L[46][5] = l_cell_wire[29];							inform_L[15][5] = l_cell_wire[30];							inform_L[47][5] = l_cell_wire[31];							inform_L[16][5] = l_cell_wire[32];							inform_L[48][5] = l_cell_wire[33];							inform_L[17][5] = l_cell_wire[34];							inform_L[49][5] = l_cell_wire[35];							inform_L[18][5] = l_cell_wire[36];							inform_L[50][5] = l_cell_wire[37];							inform_L[19][5] = l_cell_wire[38];							inform_L[51][5] = l_cell_wire[39];							inform_L[20][5] = l_cell_wire[40];							inform_L[52][5] = l_cell_wire[41];							inform_L[21][5] = l_cell_wire[42];							inform_L[53][5] = l_cell_wire[43];							inform_L[22][5] = l_cell_wire[44];							inform_L[54][5] = l_cell_wire[45];							inform_L[23][5] = l_cell_wire[46];							inform_L[55][5] = l_cell_wire[47];							inform_L[24][5] = l_cell_wire[48];							inform_L[56][5] = l_cell_wire[49];							inform_L[25][5] = l_cell_wire[50];							inform_L[57][5] = l_cell_wire[51];							inform_L[26][5] = l_cell_wire[52];							inform_L[58][5] = l_cell_wire[53];							inform_L[27][5] = l_cell_wire[54];							inform_L[59][5] = l_cell_wire[55];							inform_L[28][5] = l_cell_wire[56];							inform_L[60][5] = l_cell_wire[57];							inform_L[29][5] = l_cell_wire[58];							inform_L[61][5] = l_cell_wire[59];							inform_L[30][5] = l_cell_wire[60];							inform_L[62][5] = l_cell_wire[61];							inform_L[31][5] = l_cell_wire[62];							inform_L[63][5] = l_cell_wire[63];							inform_L[64][5] = l_cell_wire[64];							inform_L[96][5] = l_cell_wire[65];							inform_L[65][5] = l_cell_wire[66];							inform_L[97][5] = l_cell_wire[67];							inform_L[66][5] = l_cell_wire[68];							inform_L[98][5] = l_cell_wire[69];							inform_L[67][5] = l_cell_wire[70];							inform_L[99][5] = l_cell_wire[71];							inform_L[68][5] = l_cell_wire[72];							inform_L[100][5] = l_cell_wire[73];							inform_L[69][5] = l_cell_wire[74];							inform_L[101][5] = l_cell_wire[75];							inform_L[70][5] = l_cell_wire[76];							inform_L[102][5] = l_cell_wire[77];							inform_L[71][5] = l_cell_wire[78];							inform_L[103][5] = l_cell_wire[79];							inform_L[72][5] = l_cell_wire[80];							inform_L[104][5] = l_cell_wire[81];							inform_L[73][5] = l_cell_wire[82];							inform_L[105][5] = l_cell_wire[83];							inform_L[74][5] = l_cell_wire[84];							inform_L[106][5] = l_cell_wire[85];							inform_L[75][5] = l_cell_wire[86];							inform_L[107][5] = l_cell_wire[87];							inform_L[76][5] = l_cell_wire[88];							inform_L[108][5] = l_cell_wire[89];							inform_L[77][5] = l_cell_wire[90];							inform_L[109][5] = l_cell_wire[91];							inform_L[78][5] = l_cell_wire[92];							inform_L[110][5] = l_cell_wire[93];							inform_L[79][5] = l_cell_wire[94];							inform_L[111][5] = l_cell_wire[95];							inform_L[80][5] = l_cell_wire[96];							inform_L[112][5] = l_cell_wire[97];							inform_L[81][5] = l_cell_wire[98];							inform_L[113][5] = l_cell_wire[99];							inform_L[82][5] = l_cell_wire[100];							inform_L[114][5] = l_cell_wire[101];							inform_L[83][5] = l_cell_wire[102];							inform_L[115][5] = l_cell_wire[103];							inform_L[84][5] = l_cell_wire[104];							inform_L[116][5] = l_cell_wire[105];							inform_L[85][5] = l_cell_wire[106];							inform_L[117][5] = l_cell_wire[107];							inform_L[86][5] = l_cell_wire[108];							inform_L[118][5] = l_cell_wire[109];							inform_L[87][5] = l_cell_wire[110];							inform_L[119][5] = l_cell_wire[111];							inform_L[88][5] = l_cell_wire[112];							inform_L[120][5] = l_cell_wire[113];							inform_L[89][5] = l_cell_wire[114];							inform_L[121][5] = l_cell_wire[115];							inform_L[90][5] = l_cell_wire[116];							inform_L[122][5] = l_cell_wire[117];							inform_L[91][5] = l_cell_wire[118];							inform_L[123][5] = l_cell_wire[119];							inform_L[92][5] = l_cell_wire[120];							inform_L[124][5] = l_cell_wire[121];							inform_L[93][5] = l_cell_wire[122];							inform_L[125][5] = l_cell_wire[123];							inform_L[94][5] = l_cell_wire[124];							inform_L[126][5] = l_cell_wire[125];							inform_L[95][5] = l_cell_wire[126];							inform_L[127][5] = l_cell_wire[127];							inform_L[128][5] = l_cell_wire[128];							inform_L[160][5] = l_cell_wire[129];							inform_L[129][5] = l_cell_wire[130];							inform_L[161][5] = l_cell_wire[131];							inform_L[130][5] = l_cell_wire[132];							inform_L[162][5] = l_cell_wire[133];							inform_L[131][5] = l_cell_wire[134];							inform_L[163][5] = l_cell_wire[135];							inform_L[132][5] = l_cell_wire[136];							inform_L[164][5] = l_cell_wire[137];							inform_L[133][5] = l_cell_wire[138];							inform_L[165][5] = l_cell_wire[139];							inform_L[134][5] = l_cell_wire[140];							inform_L[166][5] = l_cell_wire[141];							inform_L[135][5] = l_cell_wire[142];							inform_L[167][5] = l_cell_wire[143];							inform_L[136][5] = l_cell_wire[144];							inform_L[168][5] = l_cell_wire[145];							inform_L[137][5] = l_cell_wire[146];							inform_L[169][5] = l_cell_wire[147];							inform_L[138][5] = l_cell_wire[148];							inform_L[170][5] = l_cell_wire[149];							inform_L[139][5] = l_cell_wire[150];							inform_L[171][5] = l_cell_wire[151];							inform_L[140][5] = l_cell_wire[152];							inform_L[172][5] = l_cell_wire[153];							inform_L[141][5] = l_cell_wire[154];							inform_L[173][5] = l_cell_wire[155];							inform_L[142][5] = l_cell_wire[156];							inform_L[174][5] = l_cell_wire[157];							inform_L[143][5] = l_cell_wire[158];							inform_L[175][5] = l_cell_wire[159];							inform_L[144][5] = l_cell_wire[160];							inform_L[176][5] = l_cell_wire[161];							inform_L[145][5] = l_cell_wire[162];							inform_L[177][5] = l_cell_wire[163];							inform_L[146][5] = l_cell_wire[164];							inform_L[178][5] = l_cell_wire[165];							inform_L[147][5] = l_cell_wire[166];							inform_L[179][5] = l_cell_wire[167];							inform_L[148][5] = l_cell_wire[168];							inform_L[180][5] = l_cell_wire[169];							inform_L[149][5] = l_cell_wire[170];							inform_L[181][5] = l_cell_wire[171];							inform_L[150][5] = l_cell_wire[172];							inform_L[182][5] = l_cell_wire[173];							inform_L[151][5] = l_cell_wire[174];							inform_L[183][5] = l_cell_wire[175];							inform_L[152][5] = l_cell_wire[176];							inform_L[184][5] = l_cell_wire[177];							inform_L[153][5] = l_cell_wire[178];							inform_L[185][5] = l_cell_wire[179];							inform_L[154][5] = l_cell_wire[180];							inform_L[186][5] = l_cell_wire[181];							inform_L[155][5] = l_cell_wire[182];							inform_L[187][5] = l_cell_wire[183];							inform_L[156][5] = l_cell_wire[184];							inform_L[188][5] = l_cell_wire[185];							inform_L[157][5] = l_cell_wire[186];							inform_L[189][5] = l_cell_wire[187];							inform_L[158][5] = l_cell_wire[188];							inform_L[190][5] = l_cell_wire[189];							inform_L[159][5] = l_cell_wire[190];							inform_L[191][5] = l_cell_wire[191];							inform_L[192][5] = l_cell_wire[192];							inform_L[224][5] = l_cell_wire[193];							inform_L[193][5] = l_cell_wire[194];							inform_L[225][5] = l_cell_wire[195];							inform_L[194][5] = l_cell_wire[196];							inform_L[226][5] = l_cell_wire[197];							inform_L[195][5] = l_cell_wire[198];							inform_L[227][5] = l_cell_wire[199];							inform_L[196][5] = l_cell_wire[200];							inform_L[228][5] = l_cell_wire[201];							inform_L[197][5] = l_cell_wire[202];							inform_L[229][5] = l_cell_wire[203];							inform_L[198][5] = l_cell_wire[204];							inform_L[230][5] = l_cell_wire[205];							inform_L[199][5] = l_cell_wire[206];							inform_L[231][5] = l_cell_wire[207];							inform_L[200][5] = l_cell_wire[208];							inform_L[232][5] = l_cell_wire[209];							inform_L[201][5] = l_cell_wire[210];							inform_L[233][5] = l_cell_wire[211];							inform_L[202][5] = l_cell_wire[212];							inform_L[234][5] = l_cell_wire[213];							inform_L[203][5] = l_cell_wire[214];							inform_L[235][5] = l_cell_wire[215];							inform_L[204][5] = l_cell_wire[216];							inform_L[236][5] = l_cell_wire[217];							inform_L[205][5] = l_cell_wire[218];							inform_L[237][5] = l_cell_wire[219];							inform_L[206][5] = l_cell_wire[220];							inform_L[238][5] = l_cell_wire[221];							inform_L[207][5] = l_cell_wire[222];							inform_L[239][5] = l_cell_wire[223];							inform_L[208][5] = l_cell_wire[224];							inform_L[240][5] = l_cell_wire[225];							inform_L[209][5] = l_cell_wire[226];							inform_L[241][5] = l_cell_wire[227];							inform_L[210][5] = l_cell_wire[228];							inform_L[242][5] = l_cell_wire[229];							inform_L[211][5] = l_cell_wire[230];							inform_L[243][5] = l_cell_wire[231];							inform_L[212][5] = l_cell_wire[232];							inform_L[244][5] = l_cell_wire[233];							inform_L[213][5] = l_cell_wire[234];							inform_L[245][5] = l_cell_wire[235];							inform_L[214][5] = l_cell_wire[236];							inform_L[246][5] = l_cell_wire[237];							inform_L[215][5] = l_cell_wire[238];							inform_L[247][5] = l_cell_wire[239];							inform_L[216][5] = l_cell_wire[240];							inform_L[248][5] = l_cell_wire[241];							inform_L[217][5] = l_cell_wire[242];							inform_L[249][5] = l_cell_wire[243];							inform_L[218][5] = l_cell_wire[244];							inform_L[250][5] = l_cell_wire[245];							inform_L[219][5] = l_cell_wire[246];							inform_L[251][5] = l_cell_wire[247];							inform_L[220][5] = l_cell_wire[248];							inform_L[252][5] = l_cell_wire[249];							inform_L[221][5] = l_cell_wire[250];							inform_L[253][5] = l_cell_wire[251];							inform_L[222][5] = l_cell_wire[252];							inform_L[254][5] = l_cell_wire[253];							inform_L[223][5] = l_cell_wire[254];							inform_L[255][5] = l_cell_wire[255];							inform_L[256][5] = l_cell_wire[256];							inform_L[288][5] = l_cell_wire[257];							inform_L[257][5] = l_cell_wire[258];							inform_L[289][5] = l_cell_wire[259];							inform_L[258][5] = l_cell_wire[260];							inform_L[290][5] = l_cell_wire[261];							inform_L[259][5] = l_cell_wire[262];							inform_L[291][5] = l_cell_wire[263];							inform_L[260][5] = l_cell_wire[264];							inform_L[292][5] = l_cell_wire[265];							inform_L[261][5] = l_cell_wire[266];							inform_L[293][5] = l_cell_wire[267];							inform_L[262][5] = l_cell_wire[268];							inform_L[294][5] = l_cell_wire[269];							inform_L[263][5] = l_cell_wire[270];							inform_L[295][5] = l_cell_wire[271];							inform_L[264][5] = l_cell_wire[272];							inform_L[296][5] = l_cell_wire[273];							inform_L[265][5] = l_cell_wire[274];							inform_L[297][5] = l_cell_wire[275];							inform_L[266][5] = l_cell_wire[276];							inform_L[298][5] = l_cell_wire[277];							inform_L[267][5] = l_cell_wire[278];							inform_L[299][5] = l_cell_wire[279];							inform_L[268][5] = l_cell_wire[280];							inform_L[300][5] = l_cell_wire[281];							inform_L[269][5] = l_cell_wire[282];							inform_L[301][5] = l_cell_wire[283];							inform_L[270][5] = l_cell_wire[284];							inform_L[302][5] = l_cell_wire[285];							inform_L[271][5] = l_cell_wire[286];							inform_L[303][5] = l_cell_wire[287];							inform_L[272][5] = l_cell_wire[288];							inform_L[304][5] = l_cell_wire[289];							inform_L[273][5] = l_cell_wire[290];							inform_L[305][5] = l_cell_wire[291];							inform_L[274][5] = l_cell_wire[292];							inform_L[306][5] = l_cell_wire[293];							inform_L[275][5] = l_cell_wire[294];							inform_L[307][5] = l_cell_wire[295];							inform_L[276][5] = l_cell_wire[296];							inform_L[308][5] = l_cell_wire[297];							inform_L[277][5] = l_cell_wire[298];							inform_L[309][5] = l_cell_wire[299];							inform_L[278][5] = l_cell_wire[300];							inform_L[310][5] = l_cell_wire[301];							inform_L[279][5] = l_cell_wire[302];							inform_L[311][5] = l_cell_wire[303];							inform_L[280][5] = l_cell_wire[304];							inform_L[312][5] = l_cell_wire[305];							inform_L[281][5] = l_cell_wire[306];							inform_L[313][5] = l_cell_wire[307];							inform_L[282][5] = l_cell_wire[308];							inform_L[314][5] = l_cell_wire[309];							inform_L[283][5] = l_cell_wire[310];							inform_L[315][5] = l_cell_wire[311];							inform_L[284][5] = l_cell_wire[312];							inform_L[316][5] = l_cell_wire[313];							inform_L[285][5] = l_cell_wire[314];							inform_L[317][5] = l_cell_wire[315];							inform_L[286][5] = l_cell_wire[316];							inform_L[318][5] = l_cell_wire[317];							inform_L[287][5] = l_cell_wire[318];							inform_L[319][5] = l_cell_wire[319];							inform_L[320][5] = l_cell_wire[320];							inform_L[352][5] = l_cell_wire[321];							inform_L[321][5] = l_cell_wire[322];							inform_L[353][5] = l_cell_wire[323];							inform_L[322][5] = l_cell_wire[324];							inform_L[354][5] = l_cell_wire[325];							inform_L[323][5] = l_cell_wire[326];							inform_L[355][5] = l_cell_wire[327];							inform_L[324][5] = l_cell_wire[328];							inform_L[356][5] = l_cell_wire[329];							inform_L[325][5] = l_cell_wire[330];							inform_L[357][5] = l_cell_wire[331];							inform_L[326][5] = l_cell_wire[332];							inform_L[358][5] = l_cell_wire[333];							inform_L[327][5] = l_cell_wire[334];							inform_L[359][5] = l_cell_wire[335];							inform_L[328][5] = l_cell_wire[336];							inform_L[360][5] = l_cell_wire[337];							inform_L[329][5] = l_cell_wire[338];							inform_L[361][5] = l_cell_wire[339];							inform_L[330][5] = l_cell_wire[340];							inform_L[362][5] = l_cell_wire[341];							inform_L[331][5] = l_cell_wire[342];							inform_L[363][5] = l_cell_wire[343];							inform_L[332][5] = l_cell_wire[344];							inform_L[364][5] = l_cell_wire[345];							inform_L[333][5] = l_cell_wire[346];							inform_L[365][5] = l_cell_wire[347];							inform_L[334][5] = l_cell_wire[348];							inform_L[366][5] = l_cell_wire[349];							inform_L[335][5] = l_cell_wire[350];							inform_L[367][5] = l_cell_wire[351];							inform_L[336][5] = l_cell_wire[352];							inform_L[368][5] = l_cell_wire[353];							inform_L[337][5] = l_cell_wire[354];							inform_L[369][5] = l_cell_wire[355];							inform_L[338][5] = l_cell_wire[356];							inform_L[370][5] = l_cell_wire[357];							inform_L[339][5] = l_cell_wire[358];							inform_L[371][5] = l_cell_wire[359];							inform_L[340][5] = l_cell_wire[360];							inform_L[372][5] = l_cell_wire[361];							inform_L[341][5] = l_cell_wire[362];							inform_L[373][5] = l_cell_wire[363];							inform_L[342][5] = l_cell_wire[364];							inform_L[374][5] = l_cell_wire[365];							inform_L[343][5] = l_cell_wire[366];							inform_L[375][5] = l_cell_wire[367];							inform_L[344][5] = l_cell_wire[368];							inform_L[376][5] = l_cell_wire[369];							inform_L[345][5] = l_cell_wire[370];							inform_L[377][5] = l_cell_wire[371];							inform_L[346][5] = l_cell_wire[372];							inform_L[378][5] = l_cell_wire[373];							inform_L[347][5] = l_cell_wire[374];							inform_L[379][5] = l_cell_wire[375];							inform_L[348][5] = l_cell_wire[376];							inform_L[380][5] = l_cell_wire[377];							inform_L[349][5] = l_cell_wire[378];							inform_L[381][5] = l_cell_wire[379];							inform_L[350][5] = l_cell_wire[380];							inform_L[382][5] = l_cell_wire[381];							inform_L[351][5] = l_cell_wire[382];							inform_L[383][5] = l_cell_wire[383];							inform_L[384][5] = l_cell_wire[384];							inform_L[416][5] = l_cell_wire[385];							inform_L[385][5] = l_cell_wire[386];							inform_L[417][5] = l_cell_wire[387];							inform_L[386][5] = l_cell_wire[388];							inform_L[418][5] = l_cell_wire[389];							inform_L[387][5] = l_cell_wire[390];							inform_L[419][5] = l_cell_wire[391];							inform_L[388][5] = l_cell_wire[392];							inform_L[420][5] = l_cell_wire[393];							inform_L[389][5] = l_cell_wire[394];							inform_L[421][5] = l_cell_wire[395];							inform_L[390][5] = l_cell_wire[396];							inform_L[422][5] = l_cell_wire[397];							inform_L[391][5] = l_cell_wire[398];							inform_L[423][5] = l_cell_wire[399];							inform_L[392][5] = l_cell_wire[400];							inform_L[424][5] = l_cell_wire[401];							inform_L[393][5] = l_cell_wire[402];							inform_L[425][5] = l_cell_wire[403];							inform_L[394][5] = l_cell_wire[404];							inform_L[426][5] = l_cell_wire[405];							inform_L[395][5] = l_cell_wire[406];							inform_L[427][5] = l_cell_wire[407];							inform_L[396][5] = l_cell_wire[408];							inform_L[428][5] = l_cell_wire[409];							inform_L[397][5] = l_cell_wire[410];							inform_L[429][5] = l_cell_wire[411];							inform_L[398][5] = l_cell_wire[412];							inform_L[430][5] = l_cell_wire[413];							inform_L[399][5] = l_cell_wire[414];							inform_L[431][5] = l_cell_wire[415];							inform_L[400][5] = l_cell_wire[416];							inform_L[432][5] = l_cell_wire[417];							inform_L[401][5] = l_cell_wire[418];							inform_L[433][5] = l_cell_wire[419];							inform_L[402][5] = l_cell_wire[420];							inform_L[434][5] = l_cell_wire[421];							inform_L[403][5] = l_cell_wire[422];							inform_L[435][5] = l_cell_wire[423];							inform_L[404][5] = l_cell_wire[424];							inform_L[436][5] = l_cell_wire[425];							inform_L[405][5] = l_cell_wire[426];							inform_L[437][5] = l_cell_wire[427];							inform_L[406][5] = l_cell_wire[428];							inform_L[438][5] = l_cell_wire[429];							inform_L[407][5] = l_cell_wire[430];							inform_L[439][5] = l_cell_wire[431];							inform_L[408][5] = l_cell_wire[432];							inform_L[440][5] = l_cell_wire[433];							inform_L[409][5] = l_cell_wire[434];							inform_L[441][5] = l_cell_wire[435];							inform_L[410][5] = l_cell_wire[436];							inform_L[442][5] = l_cell_wire[437];							inform_L[411][5] = l_cell_wire[438];							inform_L[443][5] = l_cell_wire[439];							inform_L[412][5] = l_cell_wire[440];							inform_L[444][5] = l_cell_wire[441];							inform_L[413][5] = l_cell_wire[442];							inform_L[445][5] = l_cell_wire[443];							inform_L[414][5] = l_cell_wire[444];							inform_L[446][5] = l_cell_wire[445];							inform_L[415][5] = l_cell_wire[446];							inform_L[447][5] = l_cell_wire[447];							inform_L[448][5] = l_cell_wire[448];							inform_L[480][5] = l_cell_wire[449];							inform_L[449][5] = l_cell_wire[450];							inform_L[481][5] = l_cell_wire[451];							inform_L[450][5] = l_cell_wire[452];							inform_L[482][5] = l_cell_wire[453];							inform_L[451][5] = l_cell_wire[454];							inform_L[483][5] = l_cell_wire[455];							inform_L[452][5] = l_cell_wire[456];							inform_L[484][5] = l_cell_wire[457];							inform_L[453][5] = l_cell_wire[458];							inform_L[485][5] = l_cell_wire[459];							inform_L[454][5] = l_cell_wire[460];							inform_L[486][5] = l_cell_wire[461];							inform_L[455][5] = l_cell_wire[462];							inform_L[487][5] = l_cell_wire[463];							inform_L[456][5] = l_cell_wire[464];							inform_L[488][5] = l_cell_wire[465];							inform_L[457][5] = l_cell_wire[466];							inform_L[489][5] = l_cell_wire[467];							inform_L[458][5] = l_cell_wire[468];							inform_L[490][5] = l_cell_wire[469];							inform_L[459][5] = l_cell_wire[470];							inform_L[491][5] = l_cell_wire[471];							inform_L[460][5] = l_cell_wire[472];							inform_L[492][5] = l_cell_wire[473];							inform_L[461][5] = l_cell_wire[474];							inform_L[493][5] = l_cell_wire[475];							inform_L[462][5] = l_cell_wire[476];							inform_L[494][5] = l_cell_wire[477];							inform_L[463][5] = l_cell_wire[478];							inform_L[495][5] = l_cell_wire[479];							inform_L[464][5] = l_cell_wire[480];							inform_L[496][5] = l_cell_wire[481];							inform_L[465][5] = l_cell_wire[482];							inform_L[497][5] = l_cell_wire[483];							inform_L[466][5] = l_cell_wire[484];							inform_L[498][5] = l_cell_wire[485];							inform_L[467][5] = l_cell_wire[486];							inform_L[499][5] = l_cell_wire[487];							inform_L[468][5] = l_cell_wire[488];							inform_L[500][5] = l_cell_wire[489];							inform_L[469][5] = l_cell_wire[490];							inform_L[501][5] = l_cell_wire[491];							inform_L[470][5] = l_cell_wire[492];							inform_L[502][5] = l_cell_wire[493];							inform_L[471][5] = l_cell_wire[494];							inform_L[503][5] = l_cell_wire[495];							inform_L[472][5] = l_cell_wire[496];							inform_L[504][5] = l_cell_wire[497];							inform_L[473][5] = l_cell_wire[498];							inform_L[505][5] = l_cell_wire[499];							inform_L[474][5] = l_cell_wire[500];							inform_L[506][5] = l_cell_wire[501];							inform_L[475][5] = l_cell_wire[502];							inform_L[507][5] = l_cell_wire[503];							inform_L[476][5] = l_cell_wire[504];							inform_L[508][5] = l_cell_wire[505];							inform_L[477][5] = l_cell_wire[506];							inform_L[509][5] = l_cell_wire[507];							inform_L[478][5] = l_cell_wire[508];							inform_L[510][5] = l_cell_wire[509];							inform_L[479][5] = l_cell_wire[510];							inform_L[511][5] = l_cell_wire[511];							inform_L[512][5] = l_cell_wire[512];							inform_L[544][5] = l_cell_wire[513];							inform_L[513][5] = l_cell_wire[514];							inform_L[545][5] = l_cell_wire[515];							inform_L[514][5] = l_cell_wire[516];							inform_L[546][5] = l_cell_wire[517];							inform_L[515][5] = l_cell_wire[518];							inform_L[547][5] = l_cell_wire[519];							inform_L[516][5] = l_cell_wire[520];							inform_L[548][5] = l_cell_wire[521];							inform_L[517][5] = l_cell_wire[522];							inform_L[549][5] = l_cell_wire[523];							inform_L[518][5] = l_cell_wire[524];							inform_L[550][5] = l_cell_wire[525];							inform_L[519][5] = l_cell_wire[526];							inform_L[551][5] = l_cell_wire[527];							inform_L[520][5] = l_cell_wire[528];							inform_L[552][5] = l_cell_wire[529];							inform_L[521][5] = l_cell_wire[530];							inform_L[553][5] = l_cell_wire[531];							inform_L[522][5] = l_cell_wire[532];							inform_L[554][5] = l_cell_wire[533];							inform_L[523][5] = l_cell_wire[534];							inform_L[555][5] = l_cell_wire[535];							inform_L[524][5] = l_cell_wire[536];							inform_L[556][5] = l_cell_wire[537];							inform_L[525][5] = l_cell_wire[538];							inform_L[557][5] = l_cell_wire[539];							inform_L[526][5] = l_cell_wire[540];							inform_L[558][5] = l_cell_wire[541];							inform_L[527][5] = l_cell_wire[542];							inform_L[559][5] = l_cell_wire[543];							inform_L[528][5] = l_cell_wire[544];							inform_L[560][5] = l_cell_wire[545];							inform_L[529][5] = l_cell_wire[546];							inform_L[561][5] = l_cell_wire[547];							inform_L[530][5] = l_cell_wire[548];							inform_L[562][5] = l_cell_wire[549];							inform_L[531][5] = l_cell_wire[550];							inform_L[563][5] = l_cell_wire[551];							inform_L[532][5] = l_cell_wire[552];							inform_L[564][5] = l_cell_wire[553];							inform_L[533][5] = l_cell_wire[554];							inform_L[565][5] = l_cell_wire[555];							inform_L[534][5] = l_cell_wire[556];							inform_L[566][5] = l_cell_wire[557];							inform_L[535][5] = l_cell_wire[558];							inform_L[567][5] = l_cell_wire[559];							inform_L[536][5] = l_cell_wire[560];							inform_L[568][5] = l_cell_wire[561];							inform_L[537][5] = l_cell_wire[562];							inform_L[569][5] = l_cell_wire[563];							inform_L[538][5] = l_cell_wire[564];							inform_L[570][5] = l_cell_wire[565];							inform_L[539][5] = l_cell_wire[566];							inform_L[571][5] = l_cell_wire[567];							inform_L[540][5] = l_cell_wire[568];							inform_L[572][5] = l_cell_wire[569];							inform_L[541][5] = l_cell_wire[570];							inform_L[573][5] = l_cell_wire[571];							inform_L[542][5] = l_cell_wire[572];							inform_L[574][5] = l_cell_wire[573];							inform_L[543][5] = l_cell_wire[574];							inform_L[575][5] = l_cell_wire[575];							inform_L[576][5] = l_cell_wire[576];							inform_L[608][5] = l_cell_wire[577];							inform_L[577][5] = l_cell_wire[578];							inform_L[609][5] = l_cell_wire[579];							inform_L[578][5] = l_cell_wire[580];							inform_L[610][5] = l_cell_wire[581];							inform_L[579][5] = l_cell_wire[582];							inform_L[611][5] = l_cell_wire[583];							inform_L[580][5] = l_cell_wire[584];							inform_L[612][5] = l_cell_wire[585];							inform_L[581][5] = l_cell_wire[586];							inform_L[613][5] = l_cell_wire[587];							inform_L[582][5] = l_cell_wire[588];							inform_L[614][5] = l_cell_wire[589];							inform_L[583][5] = l_cell_wire[590];							inform_L[615][5] = l_cell_wire[591];							inform_L[584][5] = l_cell_wire[592];							inform_L[616][5] = l_cell_wire[593];							inform_L[585][5] = l_cell_wire[594];							inform_L[617][5] = l_cell_wire[595];							inform_L[586][5] = l_cell_wire[596];							inform_L[618][5] = l_cell_wire[597];							inform_L[587][5] = l_cell_wire[598];							inform_L[619][5] = l_cell_wire[599];							inform_L[588][5] = l_cell_wire[600];							inform_L[620][5] = l_cell_wire[601];							inform_L[589][5] = l_cell_wire[602];							inform_L[621][5] = l_cell_wire[603];							inform_L[590][5] = l_cell_wire[604];							inform_L[622][5] = l_cell_wire[605];							inform_L[591][5] = l_cell_wire[606];							inform_L[623][5] = l_cell_wire[607];							inform_L[592][5] = l_cell_wire[608];							inform_L[624][5] = l_cell_wire[609];							inform_L[593][5] = l_cell_wire[610];							inform_L[625][5] = l_cell_wire[611];							inform_L[594][5] = l_cell_wire[612];							inform_L[626][5] = l_cell_wire[613];							inform_L[595][5] = l_cell_wire[614];							inform_L[627][5] = l_cell_wire[615];							inform_L[596][5] = l_cell_wire[616];							inform_L[628][5] = l_cell_wire[617];							inform_L[597][5] = l_cell_wire[618];							inform_L[629][5] = l_cell_wire[619];							inform_L[598][5] = l_cell_wire[620];							inform_L[630][5] = l_cell_wire[621];							inform_L[599][5] = l_cell_wire[622];							inform_L[631][5] = l_cell_wire[623];							inform_L[600][5] = l_cell_wire[624];							inform_L[632][5] = l_cell_wire[625];							inform_L[601][5] = l_cell_wire[626];							inform_L[633][5] = l_cell_wire[627];							inform_L[602][5] = l_cell_wire[628];							inform_L[634][5] = l_cell_wire[629];							inform_L[603][5] = l_cell_wire[630];							inform_L[635][5] = l_cell_wire[631];							inform_L[604][5] = l_cell_wire[632];							inform_L[636][5] = l_cell_wire[633];							inform_L[605][5] = l_cell_wire[634];							inform_L[637][5] = l_cell_wire[635];							inform_L[606][5] = l_cell_wire[636];							inform_L[638][5] = l_cell_wire[637];							inform_L[607][5] = l_cell_wire[638];							inform_L[639][5] = l_cell_wire[639];							inform_L[640][5] = l_cell_wire[640];							inform_L[672][5] = l_cell_wire[641];							inform_L[641][5] = l_cell_wire[642];							inform_L[673][5] = l_cell_wire[643];							inform_L[642][5] = l_cell_wire[644];							inform_L[674][5] = l_cell_wire[645];							inform_L[643][5] = l_cell_wire[646];							inform_L[675][5] = l_cell_wire[647];							inform_L[644][5] = l_cell_wire[648];							inform_L[676][5] = l_cell_wire[649];							inform_L[645][5] = l_cell_wire[650];							inform_L[677][5] = l_cell_wire[651];							inform_L[646][5] = l_cell_wire[652];							inform_L[678][5] = l_cell_wire[653];							inform_L[647][5] = l_cell_wire[654];							inform_L[679][5] = l_cell_wire[655];							inform_L[648][5] = l_cell_wire[656];							inform_L[680][5] = l_cell_wire[657];							inform_L[649][5] = l_cell_wire[658];							inform_L[681][5] = l_cell_wire[659];							inform_L[650][5] = l_cell_wire[660];							inform_L[682][5] = l_cell_wire[661];							inform_L[651][5] = l_cell_wire[662];							inform_L[683][5] = l_cell_wire[663];							inform_L[652][5] = l_cell_wire[664];							inform_L[684][5] = l_cell_wire[665];							inform_L[653][5] = l_cell_wire[666];							inform_L[685][5] = l_cell_wire[667];							inform_L[654][5] = l_cell_wire[668];							inform_L[686][5] = l_cell_wire[669];							inform_L[655][5] = l_cell_wire[670];							inform_L[687][5] = l_cell_wire[671];							inform_L[656][5] = l_cell_wire[672];							inform_L[688][5] = l_cell_wire[673];							inform_L[657][5] = l_cell_wire[674];							inform_L[689][5] = l_cell_wire[675];							inform_L[658][5] = l_cell_wire[676];							inform_L[690][5] = l_cell_wire[677];							inform_L[659][5] = l_cell_wire[678];							inform_L[691][5] = l_cell_wire[679];							inform_L[660][5] = l_cell_wire[680];							inform_L[692][5] = l_cell_wire[681];							inform_L[661][5] = l_cell_wire[682];							inform_L[693][5] = l_cell_wire[683];							inform_L[662][5] = l_cell_wire[684];							inform_L[694][5] = l_cell_wire[685];							inform_L[663][5] = l_cell_wire[686];							inform_L[695][5] = l_cell_wire[687];							inform_L[664][5] = l_cell_wire[688];							inform_L[696][5] = l_cell_wire[689];							inform_L[665][5] = l_cell_wire[690];							inform_L[697][5] = l_cell_wire[691];							inform_L[666][5] = l_cell_wire[692];							inform_L[698][5] = l_cell_wire[693];							inform_L[667][5] = l_cell_wire[694];							inform_L[699][5] = l_cell_wire[695];							inform_L[668][5] = l_cell_wire[696];							inform_L[700][5] = l_cell_wire[697];							inform_L[669][5] = l_cell_wire[698];							inform_L[701][5] = l_cell_wire[699];							inform_L[670][5] = l_cell_wire[700];							inform_L[702][5] = l_cell_wire[701];							inform_L[671][5] = l_cell_wire[702];							inform_L[703][5] = l_cell_wire[703];							inform_L[704][5] = l_cell_wire[704];							inform_L[736][5] = l_cell_wire[705];							inform_L[705][5] = l_cell_wire[706];							inform_L[737][5] = l_cell_wire[707];							inform_L[706][5] = l_cell_wire[708];							inform_L[738][5] = l_cell_wire[709];							inform_L[707][5] = l_cell_wire[710];							inform_L[739][5] = l_cell_wire[711];							inform_L[708][5] = l_cell_wire[712];							inform_L[740][5] = l_cell_wire[713];							inform_L[709][5] = l_cell_wire[714];							inform_L[741][5] = l_cell_wire[715];							inform_L[710][5] = l_cell_wire[716];							inform_L[742][5] = l_cell_wire[717];							inform_L[711][5] = l_cell_wire[718];							inform_L[743][5] = l_cell_wire[719];							inform_L[712][5] = l_cell_wire[720];							inform_L[744][5] = l_cell_wire[721];							inform_L[713][5] = l_cell_wire[722];							inform_L[745][5] = l_cell_wire[723];							inform_L[714][5] = l_cell_wire[724];							inform_L[746][5] = l_cell_wire[725];							inform_L[715][5] = l_cell_wire[726];							inform_L[747][5] = l_cell_wire[727];							inform_L[716][5] = l_cell_wire[728];							inform_L[748][5] = l_cell_wire[729];							inform_L[717][5] = l_cell_wire[730];							inform_L[749][5] = l_cell_wire[731];							inform_L[718][5] = l_cell_wire[732];							inform_L[750][5] = l_cell_wire[733];							inform_L[719][5] = l_cell_wire[734];							inform_L[751][5] = l_cell_wire[735];							inform_L[720][5] = l_cell_wire[736];							inform_L[752][5] = l_cell_wire[737];							inform_L[721][5] = l_cell_wire[738];							inform_L[753][5] = l_cell_wire[739];							inform_L[722][5] = l_cell_wire[740];							inform_L[754][5] = l_cell_wire[741];							inform_L[723][5] = l_cell_wire[742];							inform_L[755][5] = l_cell_wire[743];							inform_L[724][5] = l_cell_wire[744];							inform_L[756][5] = l_cell_wire[745];							inform_L[725][5] = l_cell_wire[746];							inform_L[757][5] = l_cell_wire[747];							inform_L[726][5] = l_cell_wire[748];							inform_L[758][5] = l_cell_wire[749];							inform_L[727][5] = l_cell_wire[750];							inform_L[759][5] = l_cell_wire[751];							inform_L[728][5] = l_cell_wire[752];							inform_L[760][5] = l_cell_wire[753];							inform_L[729][5] = l_cell_wire[754];							inform_L[761][5] = l_cell_wire[755];							inform_L[730][5] = l_cell_wire[756];							inform_L[762][5] = l_cell_wire[757];							inform_L[731][5] = l_cell_wire[758];							inform_L[763][5] = l_cell_wire[759];							inform_L[732][5] = l_cell_wire[760];							inform_L[764][5] = l_cell_wire[761];							inform_L[733][5] = l_cell_wire[762];							inform_L[765][5] = l_cell_wire[763];							inform_L[734][5] = l_cell_wire[764];							inform_L[766][5] = l_cell_wire[765];							inform_L[735][5] = l_cell_wire[766];							inform_L[767][5] = l_cell_wire[767];							inform_L[768][5] = l_cell_wire[768];							inform_L[800][5] = l_cell_wire[769];							inform_L[769][5] = l_cell_wire[770];							inform_L[801][5] = l_cell_wire[771];							inform_L[770][5] = l_cell_wire[772];							inform_L[802][5] = l_cell_wire[773];							inform_L[771][5] = l_cell_wire[774];							inform_L[803][5] = l_cell_wire[775];							inform_L[772][5] = l_cell_wire[776];							inform_L[804][5] = l_cell_wire[777];							inform_L[773][5] = l_cell_wire[778];							inform_L[805][5] = l_cell_wire[779];							inform_L[774][5] = l_cell_wire[780];							inform_L[806][5] = l_cell_wire[781];							inform_L[775][5] = l_cell_wire[782];							inform_L[807][5] = l_cell_wire[783];							inform_L[776][5] = l_cell_wire[784];							inform_L[808][5] = l_cell_wire[785];							inform_L[777][5] = l_cell_wire[786];							inform_L[809][5] = l_cell_wire[787];							inform_L[778][5] = l_cell_wire[788];							inform_L[810][5] = l_cell_wire[789];							inform_L[779][5] = l_cell_wire[790];							inform_L[811][5] = l_cell_wire[791];							inform_L[780][5] = l_cell_wire[792];							inform_L[812][5] = l_cell_wire[793];							inform_L[781][5] = l_cell_wire[794];							inform_L[813][5] = l_cell_wire[795];							inform_L[782][5] = l_cell_wire[796];							inform_L[814][5] = l_cell_wire[797];							inform_L[783][5] = l_cell_wire[798];							inform_L[815][5] = l_cell_wire[799];							inform_L[784][5] = l_cell_wire[800];							inform_L[816][5] = l_cell_wire[801];							inform_L[785][5] = l_cell_wire[802];							inform_L[817][5] = l_cell_wire[803];							inform_L[786][5] = l_cell_wire[804];							inform_L[818][5] = l_cell_wire[805];							inform_L[787][5] = l_cell_wire[806];							inform_L[819][5] = l_cell_wire[807];							inform_L[788][5] = l_cell_wire[808];							inform_L[820][5] = l_cell_wire[809];							inform_L[789][5] = l_cell_wire[810];							inform_L[821][5] = l_cell_wire[811];							inform_L[790][5] = l_cell_wire[812];							inform_L[822][5] = l_cell_wire[813];							inform_L[791][5] = l_cell_wire[814];							inform_L[823][5] = l_cell_wire[815];							inform_L[792][5] = l_cell_wire[816];							inform_L[824][5] = l_cell_wire[817];							inform_L[793][5] = l_cell_wire[818];							inform_L[825][5] = l_cell_wire[819];							inform_L[794][5] = l_cell_wire[820];							inform_L[826][5] = l_cell_wire[821];							inform_L[795][5] = l_cell_wire[822];							inform_L[827][5] = l_cell_wire[823];							inform_L[796][5] = l_cell_wire[824];							inform_L[828][5] = l_cell_wire[825];							inform_L[797][5] = l_cell_wire[826];							inform_L[829][5] = l_cell_wire[827];							inform_L[798][5] = l_cell_wire[828];							inform_L[830][5] = l_cell_wire[829];							inform_L[799][5] = l_cell_wire[830];							inform_L[831][5] = l_cell_wire[831];							inform_L[832][5] = l_cell_wire[832];							inform_L[864][5] = l_cell_wire[833];							inform_L[833][5] = l_cell_wire[834];							inform_L[865][5] = l_cell_wire[835];							inform_L[834][5] = l_cell_wire[836];							inform_L[866][5] = l_cell_wire[837];							inform_L[835][5] = l_cell_wire[838];							inform_L[867][5] = l_cell_wire[839];							inform_L[836][5] = l_cell_wire[840];							inform_L[868][5] = l_cell_wire[841];							inform_L[837][5] = l_cell_wire[842];							inform_L[869][5] = l_cell_wire[843];							inform_L[838][5] = l_cell_wire[844];							inform_L[870][5] = l_cell_wire[845];							inform_L[839][5] = l_cell_wire[846];							inform_L[871][5] = l_cell_wire[847];							inform_L[840][5] = l_cell_wire[848];							inform_L[872][5] = l_cell_wire[849];							inform_L[841][5] = l_cell_wire[850];							inform_L[873][5] = l_cell_wire[851];							inform_L[842][5] = l_cell_wire[852];							inform_L[874][5] = l_cell_wire[853];							inform_L[843][5] = l_cell_wire[854];							inform_L[875][5] = l_cell_wire[855];							inform_L[844][5] = l_cell_wire[856];							inform_L[876][5] = l_cell_wire[857];							inform_L[845][5] = l_cell_wire[858];							inform_L[877][5] = l_cell_wire[859];							inform_L[846][5] = l_cell_wire[860];							inform_L[878][5] = l_cell_wire[861];							inform_L[847][5] = l_cell_wire[862];							inform_L[879][5] = l_cell_wire[863];							inform_L[848][5] = l_cell_wire[864];							inform_L[880][5] = l_cell_wire[865];							inform_L[849][5] = l_cell_wire[866];							inform_L[881][5] = l_cell_wire[867];							inform_L[850][5] = l_cell_wire[868];							inform_L[882][5] = l_cell_wire[869];							inform_L[851][5] = l_cell_wire[870];							inform_L[883][5] = l_cell_wire[871];							inform_L[852][5] = l_cell_wire[872];							inform_L[884][5] = l_cell_wire[873];							inform_L[853][5] = l_cell_wire[874];							inform_L[885][5] = l_cell_wire[875];							inform_L[854][5] = l_cell_wire[876];							inform_L[886][5] = l_cell_wire[877];							inform_L[855][5] = l_cell_wire[878];							inform_L[887][5] = l_cell_wire[879];							inform_L[856][5] = l_cell_wire[880];							inform_L[888][5] = l_cell_wire[881];							inform_L[857][5] = l_cell_wire[882];							inform_L[889][5] = l_cell_wire[883];							inform_L[858][5] = l_cell_wire[884];							inform_L[890][5] = l_cell_wire[885];							inform_L[859][5] = l_cell_wire[886];							inform_L[891][5] = l_cell_wire[887];							inform_L[860][5] = l_cell_wire[888];							inform_L[892][5] = l_cell_wire[889];							inform_L[861][5] = l_cell_wire[890];							inform_L[893][5] = l_cell_wire[891];							inform_L[862][5] = l_cell_wire[892];							inform_L[894][5] = l_cell_wire[893];							inform_L[863][5] = l_cell_wire[894];							inform_L[895][5] = l_cell_wire[895];							inform_L[896][5] = l_cell_wire[896];							inform_L[928][5] = l_cell_wire[897];							inform_L[897][5] = l_cell_wire[898];							inform_L[929][5] = l_cell_wire[899];							inform_L[898][5] = l_cell_wire[900];							inform_L[930][5] = l_cell_wire[901];							inform_L[899][5] = l_cell_wire[902];							inform_L[931][5] = l_cell_wire[903];							inform_L[900][5] = l_cell_wire[904];							inform_L[932][5] = l_cell_wire[905];							inform_L[901][5] = l_cell_wire[906];							inform_L[933][5] = l_cell_wire[907];							inform_L[902][5] = l_cell_wire[908];							inform_L[934][5] = l_cell_wire[909];							inform_L[903][5] = l_cell_wire[910];							inform_L[935][5] = l_cell_wire[911];							inform_L[904][5] = l_cell_wire[912];							inform_L[936][5] = l_cell_wire[913];							inform_L[905][5] = l_cell_wire[914];							inform_L[937][5] = l_cell_wire[915];							inform_L[906][5] = l_cell_wire[916];							inform_L[938][5] = l_cell_wire[917];							inform_L[907][5] = l_cell_wire[918];							inform_L[939][5] = l_cell_wire[919];							inform_L[908][5] = l_cell_wire[920];							inform_L[940][5] = l_cell_wire[921];							inform_L[909][5] = l_cell_wire[922];							inform_L[941][5] = l_cell_wire[923];							inform_L[910][5] = l_cell_wire[924];							inform_L[942][5] = l_cell_wire[925];							inform_L[911][5] = l_cell_wire[926];							inform_L[943][5] = l_cell_wire[927];							inform_L[912][5] = l_cell_wire[928];							inform_L[944][5] = l_cell_wire[929];							inform_L[913][5] = l_cell_wire[930];							inform_L[945][5] = l_cell_wire[931];							inform_L[914][5] = l_cell_wire[932];							inform_L[946][5] = l_cell_wire[933];							inform_L[915][5] = l_cell_wire[934];							inform_L[947][5] = l_cell_wire[935];							inform_L[916][5] = l_cell_wire[936];							inform_L[948][5] = l_cell_wire[937];							inform_L[917][5] = l_cell_wire[938];							inform_L[949][5] = l_cell_wire[939];							inform_L[918][5] = l_cell_wire[940];							inform_L[950][5] = l_cell_wire[941];							inform_L[919][5] = l_cell_wire[942];							inform_L[951][5] = l_cell_wire[943];							inform_L[920][5] = l_cell_wire[944];							inform_L[952][5] = l_cell_wire[945];							inform_L[921][5] = l_cell_wire[946];							inform_L[953][5] = l_cell_wire[947];							inform_L[922][5] = l_cell_wire[948];							inform_L[954][5] = l_cell_wire[949];							inform_L[923][5] = l_cell_wire[950];							inform_L[955][5] = l_cell_wire[951];							inform_L[924][5] = l_cell_wire[952];							inform_L[956][5] = l_cell_wire[953];							inform_L[925][5] = l_cell_wire[954];							inform_L[957][5] = l_cell_wire[955];							inform_L[926][5] = l_cell_wire[956];							inform_L[958][5] = l_cell_wire[957];							inform_L[927][5] = l_cell_wire[958];							inform_L[959][5] = l_cell_wire[959];							inform_L[960][5] = l_cell_wire[960];							inform_L[992][5] = l_cell_wire[961];							inform_L[961][5] = l_cell_wire[962];							inform_L[993][5] = l_cell_wire[963];							inform_L[962][5] = l_cell_wire[964];							inform_L[994][5] = l_cell_wire[965];							inform_L[963][5] = l_cell_wire[966];							inform_L[995][5] = l_cell_wire[967];							inform_L[964][5] = l_cell_wire[968];							inform_L[996][5] = l_cell_wire[969];							inform_L[965][5] = l_cell_wire[970];							inform_L[997][5] = l_cell_wire[971];							inform_L[966][5] = l_cell_wire[972];							inform_L[998][5] = l_cell_wire[973];							inform_L[967][5] = l_cell_wire[974];							inform_L[999][5] = l_cell_wire[975];							inform_L[968][5] = l_cell_wire[976];							inform_L[1000][5] = l_cell_wire[977];							inform_L[969][5] = l_cell_wire[978];							inform_L[1001][5] = l_cell_wire[979];							inform_L[970][5] = l_cell_wire[980];							inform_L[1002][5] = l_cell_wire[981];							inform_L[971][5] = l_cell_wire[982];							inform_L[1003][5] = l_cell_wire[983];							inform_L[972][5] = l_cell_wire[984];							inform_L[1004][5] = l_cell_wire[985];							inform_L[973][5] = l_cell_wire[986];							inform_L[1005][5] = l_cell_wire[987];							inform_L[974][5] = l_cell_wire[988];							inform_L[1006][5] = l_cell_wire[989];							inform_L[975][5] = l_cell_wire[990];							inform_L[1007][5] = l_cell_wire[991];							inform_L[976][5] = l_cell_wire[992];							inform_L[1008][5] = l_cell_wire[993];							inform_L[977][5] = l_cell_wire[994];							inform_L[1009][5] = l_cell_wire[995];							inform_L[978][5] = l_cell_wire[996];							inform_L[1010][5] = l_cell_wire[997];							inform_L[979][5] = l_cell_wire[998];							inform_L[1011][5] = l_cell_wire[999];							inform_L[980][5] = l_cell_wire[1000];							inform_L[1012][5] = l_cell_wire[1001];							inform_L[981][5] = l_cell_wire[1002];							inform_L[1013][5] = l_cell_wire[1003];							inform_L[982][5] = l_cell_wire[1004];							inform_L[1014][5] = l_cell_wire[1005];							inform_L[983][5] = l_cell_wire[1006];							inform_L[1015][5] = l_cell_wire[1007];							inform_L[984][5] = l_cell_wire[1008];							inform_L[1016][5] = l_cell_wire[1009];							inform_L[985][5] = l_cell_wire[1010];							inform_L[1017][5] = l_cell_wire[1011];							inform_L[986][5] = l_cell_wire[1012];							inform_L[1018][5] = l_cell_wire[1013];							inform_L[987][5] = l_cell_wire[1014];							inform_L[1019][5] = l_cell_wire[1015];							inform_L[988][5] = l_cell_wire[1016];							inform_L[1020][5] = l_cell_wire[1017];							inform_L[989][5] = l_cell_wire[1018];							inform_L[1021][5] = l_cell_wire[1019];							inform_L[990][5] = l_cell_wire[1020];							inform_L[1022][5] = l_cell_wire[1021];							inform_L[991][5] = l_cell_wire[1022];							inform_L[1023][5] = l_cell_wire[1023];						end
						7:						begin							inform_R[0][7] = r_cell_wire[0];							inform_R[64][7] = r_cell_wire[1];							inform_R[1][7] = r_cell_wire[2];							inform_R[65][7] = r_cell_wire[3];							inform_R[2][7] = r_cell_wire[4];							inform_R[66][7] = r_cell_wire[5];							inform_R[3][7] = r_cell_wire[6];							inform_R[67][7] = r_cell_wire[7];							inform_R[4][7] = r_cell_wire[8];							inform_R[68][7] = r_cell_wire[9];							inform_R[5][7] = r_cell_wire[10];							inform_R[69][7] = r_cell_wire[11];							inform_R[6][7] = r_cell_wire[12];							inform_R[70][7] = r_cell_wire[13];							inform_R[7][7] = r_cell_wire[14];							inform_R[71][7] = r_cell_wire[15];							inform_R[8][7] = r_cell_wire[16];							inform_R[72][7] = r_cell_wire[17];							inform_R[9][7] = r_cell_wire[18];							inform_R[73][7] = r_cell_wire[19];							inform_R[10][7] = r_cell_wire[20];							inform_R[74][7] = r_cell_wire[21];							inform_R[11][7] = r_cell_wire[22];							inform_R[75][7] = r_cell_wire[23];							inform_R[12][7] = r_cell_wire[24];							inform_R[76][7] = r_cell_wire[25];							inform_R[13][7] = r_cell_wire[26];							inform_R[77][7] = r_cell_wire[27];							inform_R[14][7] = r_cell_wire[28];							inform_R[78][7] = r_cell_wire[29];							inform_R[15][7] = r_cell_wire[30];							inform_R[79][7] = r_cell_wire[31];							inform_R[16][7] = r_cell_wire[32];							inform_R[80][7] = r_cell_wire[33];							inform_R[17][7] = r_cell_wire[34];							inform_R[81][7] = r_cell_wire[35];							inform_R[18][7] = r_cell_wire[36];							inform_R[82][7] = r_cell_wire[37];							inform_R[19][7] = r_cell_wire[38];							inform_R[83][7] = r_cell_wire[39];							inform_R[20][7] = r_cell_wire[40];							inform_R[84][7] = r_cell_wire[41];							inform_R[21][7] = r_cell_wire[42];							inform_R[85][7] = r_cell_wire[43];							inform_R[22][7] = r_cell_wire[44];							inform_R[86][7] = r_cell_wire[45];							inform_R[23][7] = r_cell_wire[46];							inform_R[87][7] = r_cell_wire[47];							inform_R[24][7] = r_cell_wire[48];							inform_R[88][7] = r_cell_wire[49];							inform_R[25][7] = r_cell_wire[50];							inform_R[89][7] = r_cell_wire[51];							inform_R[26][7] = r_cell_wire[52];							inform_R[90][7] = r_cell_wire[53];							inform_R[27][7] = r_cell_wire[54];							inform_R[91][7] = r_cell_wire[55];							inform_R[28][7] = r_cell_wire[56];							inform_R[92][7] = r_cell_wire[57];							inform_R[29][7] = r_cell_wire[58];							inform_R[93][7] = r_cell_wire[59];							inform_R[30][7] = r_cell_wire[60];							inform_R[94][7] = r_cell_wire[61];							inform_R[31][7] = r_cell_wire[62];							inform_R[95][7] = r_cell_wire[63];							inform_R[32][7] = r_cell_wire[64];							inform_R[96][7] = r_cell_wire[65];							inform_R[33][7] = r_cell_wire[66];							inform_R[97][7] = r_cell_wire[67];							inform_R[34][7] = r_cell_wire[68];							inform_R[98][7] = r_cell_wire[69];							inform_R[35][7] = r_cell_wire[70];							inform_R[99][7] = r_cell_wire[71];							inform_R[36][7] = r_cell_wire[72];							inform_R[100][7] = r_cell_wire[73];							inform_R[37][7] = r_cell_wire[74];							inform_R[101][7] = r_cell_wire[75];							inform_R[38][7] = r_cell_wire[76];							inform_R[102][7] = r_cell_wire[77];							inform_R[39][7] = r_cell_wire[78];							inform_R[103][7] = r_cell_wire[79];							inform_R[40][7] = r_cell_wire[80];							inform_R[104][7] = r_cell_wire[81];							inform_R[41][7] = r_cell_wire[82];							inform_R[105][7] = r_cell_wire[83];							inform_R[42][7] = r_cell_wire[84];							inform_R[106][7] = r_cell_wire[85];							inform_R[43][7] = r_cell_wire[86];							inform_R[107][7] = r_cell_wire[87];							inform_R[44][7] = r_cell_wire[88];							inform_R[108][7] = r_cell_wire[89];							inform_R[45][7] = r_cell_wire[90];							inform_R[109][7] = r_cell_wire[91];							inform_R[46][7] = r_cell_wire[92];							inform_R[110][7] = r_cell_wire[93];							inform_R[47][7] = r_cell_wire[94];							inform_R[111][7] = r_cell_wire[95];							inform_R[48][7] = r_cell_wire[96];							inform_R[112][7] = r_cell_wire[97];							inform_R[49][7] = r_cell_wire[98];							inform_R[113][7] = r_cell_wire[99];							inform_R[50][7] = r_cell_wire[100];							inform_R[114][7] = r_cell_wire[101];							inform_R[51][7] = r_cell_wire[102];							inform_R[115][7] = r_cell_wire[103];							inform_R[52][7] = r_cell_wire[104];							inform_R[116][7] = r_cell_wire[105];							inform_R[53][7] = r_cell_wire[106];							inform_R[117][7] = r_cell_wire[107];							inform_R[54][7] = r_cell_wire[108];							inform_R[118][7] = r_cell_wire[109];							inform_R[55][7] = r_cell_wire[110];							inform_R[119][7] = r_cell_wire[111];							inform_R[56][7] = r_cell_wire[112];							inform_R[120][7] = r_cell_wire[113];							inform_R[57][7] = r_cell_wire[114];							inform_R[121][7] = r_cell_wire[115];							inform_R[58][7] = r_cell_wire[116];							inform_R[122][7] = r_cell_wire[117];							inform_R[59][7] = r_cell_wire[118];							inform_R[123][7] = r_cell_wire[119];							inform_R[60][7] = r_cell_wire[120];							inform_R[124][7] = r_cell_wire[121];							inform_R[61][7] = r_cell_wire[122];							inform_R[125][7] = r_cell_wire[123];							inform_R[62][7] = r_cell_wire[124];							inform_R[126][7] = r_cell_wire[125];							inform_R[63][7] = r_cell_wire[126];							inform_R[127][7] = r_cell_wire[127];							inform_R[128][7] = r_cell_wire[128];							inform_R[192][7] = r_cell_wire[129];							inform_R[129][7] = r_cell_wire[130];							inform_R[193][7] = r_cell_wire[131];							inform_R[130][7] = r_cell_wire[132];							inform_R[194][7] = r_cell_wire[133];							inform_R[131][7] = r_cell_wire[134];							inform_R[195][7] = r_cell_wire[135];							inform_R[132][7] = r_cell_wire[136];							inform_R[196][7] = r_cell_wire[137];							inform_R[133][7] = r_cell_wire[138];							inform_R[197][7] = r_cell_wire[139];							inform_R[134][7] = r_cell_wire[140];							inform_R[198][7] = r_cell_wire[141];							inform_R[135][7] = r_cell_wire[142];							inform_R[199][7] = r_cell_wire[143];							inform_R[136][7] = r_cell_wire[144];							inform_R[200][7] = r_cell_wire[145];							inform_R[137][7] = r_cell_wire[146];							inform_R[201][7] = r_cell_wire[147];							inform_R[138][7] = r_cell_wire[148];							inform_R[202][7] = r_cell_wire[149];							inform_R[139][7] = r_cell_wire[150];							inform_R[203][7] = r_cell_wire[151];							inform_R[140][7] = r_cell_wire[152];							inform_R[204][7] = r_cell_wire[153];							inform_R[141][7] = r_cell_wire[154];							inform_R[205][7] = r_cell_wire[155];							inform_R[142][7] = r_cell_wire[156];							inform_R[206][7] = r_cell_wire[157];							inform_R[143][7] = r_cell_wire[158];							inform_R[207][7] = r_cell_wire[159];							inform_R[144][7] = r_cell_wire[160];							inform_R[208][7] = r_cell_wire[161];							inform_R[145][7] = r_cell_wire[162];							inform_R[209][7] = r_cell_wire[163];							inform_R[146][7] = r_cell_wire[164];							inform_R[210][7] = r_cell_wire[165];							inform_R[147][7] = r_cell_wire[166];							inform_R[211][7] = r_cell_wire[167];							inform_R[148][7] = r_cell_wire[168];							inform_R[212][7] = r_cell_wire[169];							inform_R[149][7] = r_cell_wire[170];							inform_R[213][7] = r_cell_wire[171];							inform_R[150][7] = r_cell_wire[172];							inform_R[214][7] = r_cell_wire[173];							inform_R[151][7] = r_cell_wire[174];							inform_R[215][7] = r_cell_wire[175];							inform_R[152][7] = r_cell_wire[176];							inform_R[216][7] = r_cell_wire[177];							inform_R[153][7] = r_cell_wire[178];							inform_R[217][7] = r_cell_wire[179];							inform_R[154][7] = r_cell_wire[180];							inform_R[218][7] = r_cell_wire[181];							inform_R[155][7] = r_cell_wire[182];							inform_R[219][7] = r_cell_wire[183];							inform_R[156][7] = r_cell_wire[184];							inform_R[220][7] = r_cell_wire[185];							inform_R[157][7] = r_cell_wire[186];							inform_R[221][7] = r_cell_wire[187];							inform_R[158][7] = r_cell_wire[188];							inform_R[222][7] = r_cell_wire[189];							inform_R[159][7] = r_cell_wire[190];							inform_R[223][7] = r_cell_wire[191];							inform_R[160][7] = r_cell_wire[192];							inform_R[224][7] = r_cell_wire[193];							inform_R[161][7] = r_cell_wire[194];							inform_R[225][7] = r_cell_wire[195];							inform_R[162][7] = r_cell_wire[196];							inform_R[226][7] = r_cell_wire[197];							inform_R[163][7] = r_cell_wire[198];							inform_R[227][7] = r_cell_wire[199];							inform_R[164][7] = r_cell_wire[200];							inform_R[228][7] = r_cell_wire[201];							inform_R[165][7] = r_cell_wire[202];							inform_R[229][7] = r_cell_wire[203];							inform_R[166][7] = r_cell_wire[204];							inform_R[230][7] = r_cell_wire[205];							inform_R[167][7] = r_cell_wire[206];							inform_R[231][7] = r_cell_wire[207];							inform_R[168][7] = r_cell_wire[208];							inform_R[232][7] = r_cell_wire[209];							inform_R[169][7] = r_cell_wire[210];							inform_R[233][7] = r_cell_wire[211];							inform_R[170][7] = r_cell_wire[212];							inform_R[234][7] = r_cell_wire[213];							inform_R[171][7] = r_cell_wire[214];							inform_R[235][7] = r_cell_wire[215];							inform_R[172][7] = r_cell_wire[216];							inform_R[236][7] = r_cell_wire[217];							inform_R[173][7] = r_cell_wire[218];							inform_R[237][7] = r_cell_wire[219];							inform_R[174][7] = r_cell_wire[220];							inform_R[238][7] = r_cell_wire[221];							inform_R[175][7] = r_cell_wire[222];							inform_R[239][7] = r_cell_wire[223];							inform_R[176][7] = r_cell_wire[224];							inform_R[240][7] = r_cell_wire[225];							inform_R[177][7] = r_cell_wire[226];							inform_R[241][7] = r_cell_wire[227];							inform_R[178][7] = r_cell_wire[228];							inform_R[242][7] = r_cell_wire[229];							inform_R[179][7] = r_cell_wire[230];							inform_R[243][7] = r_cell_wire[231];							inform_R[180][7] = r_cell_wire[232];							inform_R[244][7] = r_cell_wire[233];							inform_R[181][7] = r_cell_wire[234];							inform_R[245][7] = r_cell_wire[235];							inform_R[182][7] = r_cell_wire[236];							inform_R[246][7] = r_cell_wire[237];							inform_R[183][7] = r_cell_wire[238];							inform_R[247][7] = r_cell_wire[239];							inform_R[184][7] = r_cell_wire[240];							inform_R[248][7] = r_cell_wire[241];							inform_R[185][7] = r_cell_wire[242];							inform_R[249][7] = r_cell_wire[243];							inform_R[186][7] = r_cell_wire[244];							inform_R[250][7] = r_cell_wire[245];							inform_R[187][7] = r_cell_wire[246];							inform_R[251][7] = r_cell_wire[247];							inform_R[188][7] = r_cell_wire[248];							inform_R[252][7] = r_cell_wire[249];							inform_R[189][7] = r_cell_wire[250];							inform_R[253][7] = r_cell_wire[251];							inform_R[190][7] = r_cell_wire[252];							inform_R[254][7] = r_cell_wire[253];							inform_R[191][7] = r_cell_wire[254];							inform_R[255][7] = r_cell_wire[255];							inform_R[256][7] = r_cell_wire[256];							inform_R[320][7] = r_cell_wire[257];							inform_R[257][7] = r_cell_wire[258];							inform_R[321][7] = r_cell_wire[259];							inform_R[258][7] = r_cell_wire[260];							inform_R[322][7] = r_cell_wire[261];							inform_R[259][7] = r_cell_wire[262];							inform_R[323][7] = r_cell_wire[263];							inform_R[260][7] = r_cell_wire[264];							inform_R[324][7] = r_cell_wire[265];							inform_R[261][7] = r_cell_wire[266];							inform_R[325][7] = r_cell_wire[267];							inform_R[262][7] = r_cell_wire[268];							inform_R[326][7] = r_cell_wire[269];							inform_R[263][7] = r_cell_wire[270];							inform_R[327][7] = r_cell_wire[271];							inform_R[264][7] = r_cell_wire[272];							inform_R[328][7] = r_cell_wire[273];							inform_R[265][7] = r_cell_wire[274];							inform_R[329][7] = r_cell_wire[275];							inform_R[266][7] = r_cell_wire[276];							inform_R[330][7] = r_cell_wire[277];							inform_R[267][7] = r_cell_wire[278];							inform_R[331][7] = r_cell_wire[279];							inform_R[268][7] = r_cell_wire[280];							inform_R[332][7] = r_cell_wire[281];							inform_R[269][7] = r_cell_wire[282];							inform_R[333][7] = r_cell_wire[283];							inform_R[270][7] = r_cell_wire[284];							inform_R[334][7] = r_cell_wire[285];							inform_R[271][7] = r_cell_wire[286];							inform_R[335][7] = r_cell_wire[287];							inform_R[272][7] = r_cell_wire[288];							inform_R[336][7] = r_cell_wire[289];							inform_R[273][7] = r_cell_wire[290];							inform_R[337][7] = r_cell_wire[291];							inform_R[274][7] = r_cell_wire[292];							inform_R[338][7] = r_cell_wire[293];							inform_R[275][7] = r_cell_wire[294];							inform_R[339][7] = r_cell_wire[295];							inform_R[276][7] = r_cell_wire[296];							inform_R[340][7] = r_cell_wire[297];							inform_R[277][7] = r_cell_wire[298];							inform_R[341][7] = r_cell_wire[299];							inform_R[278][7] = r_cell_wire[300];							inform_R[342][7] = r_cell_wire[301];							inform_R[279][7] = r_cell_wire[302];							inform_R[343][7] = r_cell_wire[303];							inform_R[280][7] = r_cell_wire[304];							inform_R[344][7] = r_cell_wire[305];							inform_R[281][7] = r_cell_wire[306];							inform_R[345][7] = r_cell_wire[307];							inform_R[282][7] = r_cell_wire[308];							inform_R[346][7] = r_cell_wire[309];							inform_R[283][7] = r_cell_wire[310];							inform_R[347][7] = r_cell_wire[311];							inform_R[284][7] = r_cell_wire[312];							inform_R[348][7] = r_cell_wire[313];							inform_R[285][7] = r_cell_wire[314];							inform_R[349][7] = r_cell_wire[315];							inform_R[286][7] = r_cell_wire[316];							inform_R[350][7] = r_cell_wire[317];							inform_R[287][7] = r_cell_wire[318];							inform_R[351][7] = r_cell_wire[319];							inform_R[288][7] = r_cell_wire[320];							inform_R[352][7] = r_cell_wire[321];							inform_R[289][7] = r_cell_wire[322];							inform_R[353][7] = r_cell_wire[323];							inform_R[290][7] = r_cell_wire[324];							inform_R[354][7] = r_cell_wire[325];							inform_R[291][7] = r_cell_wire[326];							inform_R[355][7] = r_cell_wire[327];							inform_R[292][7] = r_cell_wire[328];							inform_R[356][7] = r_cell_wire[329];							inform_R[293][7] = r_cell_wire[330];							inform_R[357][7] = r_cell_wire[331];							inform_R[294][7] = r_cell_wire[332];							inform_R[358][7] = r_cell_wire[333];							inform_R[295][7] = r_cell_wire[334];							inform_R[359][7] = r_cell_wire[335];							inform_R[296][7] = r_cell_wire[336];							inform_R[360][7] = r_cell_wire[337];							inform_R[297][7] = r_cell_wire[338];							inform_R[361][7] = r_cell_wire[339];							inform_R[298][7] = r_cell_wire[340];							inform_R[362][7] = r_cell_wire[341];							inform_R[299][7] = r_cell_wire[342];							inform_R[363][7] = r_cell_wire[343];							inform_R[300][7] = r_cell_wire[344];							inform_R[364][7] = r_cell_wire[345];							inform_R[301][7] = r_cell_wire[346];							inform_R[365][7] = r_cell_wire[347];							inform_R[302][7] = r_cell_wire[348];							inform_R[366][7] = r_cell_wire[349];							inform_R[303][7] = r_cell_wire[350];							inform_R[367][7] = r_cell_wire[351];							inform_R[304][7] = r_cell_wire[352];							inform_R[368][7] = r_cell_wire[353];							inform_R[305][7] = r_cell_wire[354];							inform_R[369][7] = r_cell_wire[355];							inform_R[306][7] = r_cell_wire[356];							inform_R[370][7] = r_cell_wire[357];							inform_R[307][7] = r_cell_wire[358];							inform_R[371][7] = r_cell_wire[359];							inform_R[308][7] = r_cell_wire[360];							inform_R[372][7] = r_cell_wire[361];							inform_R[309][7] = r_cell_wire[362];							inform_R[373][7] = r_cell_wire[363];							inform_R[310][7] = r_cell_wire[364];							inform_R[374][7] = r_cell_wire[365];							inform_R[311][7] = r_cell_wire[366];							inform_R[375][7] = r_cell_wire[367];							inform_R[312][7] = r_cell_wire[368];							inform_R[376][7] = r_cell_wire[369];							inform_R[313][7] = r_cell_wire[370];							inform_R[377][7] = r_cell_wire[371];							inform_R[314][7] = r_cell_wire[372];							inform_R[378][7] = r_cell_wire[373];							inform_R[315][7] = r_cell_wire[374];							inform_R[379][7] = r_cell_wire[375];							inform_R[316][7] = r_cell_wire[376];							inform_R[380][7] = r_cell_wire[377];							inform_R[317][7] = r_cell_wire[378];							inform_R[381][7] = r_cell_wire[379];							inform_R[318][7] = r_cell_wire[380];							inform_R[382][7] = r_cell_wire[381];							inform_R[319][7] = r_cell_wire[382];							inform_R[383][7] = r_cell_wire[383];							inform_R[384][7] = r_cell_wire[384];							inform_R[448][7] = r_cell_wire[385];							inform_R[385][7] = r_cell_wire[386];							inform_R[449][7] = r_cell_wire[387];							inform_R[386][7] = r_cell_wire[388];							inform_R[450][7] = r_cell_wire[389];							inform_R[387][7] = r_cell_wire[390];							inform_R[451][7] = r_cell_wire[391];							inform_R[388][7] = r_cell_wire[392];							inform_R[452][7] = r_cell_wire[393];							inform_R[389][7] = r_cell_wire[394];							inform_R[453][7] = r_cell_wire[395];							inform_R[390][7] = r_cell_wire[396];							inform_R[454][7] = r_cell_wire[397];							inform_R[391][7] = r_cell_wire[398];							inform_R[455][7] = r_cell_wire[399];							inform_R[392][7] = r_cell_wire[400];							inform_R[456][7] = r_cell_wire[401];							inform_R[393][7] = r_cell_wire[402];							inform_R[457][7] = r_cell_wire[403];							inform_R[394][7] = r_cell_wire[404];							inform_R[458][7] = r_cell_wire[405];							inform_R[395][7] = r_cell_wire[406];							inform_R[459][7] = r_cell_wire[407];							inform_R[396][7] = r_cell_wire[408];							inform_R[460][7] = r_cell_wire[409];							inform_R[397][7] = r_cell_wire[410];							inform_R[461][7] = r_cell_wire[411];							inform_R[398][7] = r_cell_wire[412];							inform_R[462][7] = r_cell_wire[413];							inform_R[399][7] = r_cell_wire[414];							inform_R[463][7] = r_cell_wire[415];							inform_R[400][7] = r_cell_wire[416];							inform_R[464][7] = r_cell_wire[417];							inform_R[401][7] = r_cell_wire[418];							inform_R[465][7] = r_cell_wire[419];							inform_R[402][7] = r_cell_wire[420];							inform_R[466][7] = r_cell_wire[421];							inform_R[403][7] = r_cell_wire[422];							inform_R[467][7] = r_cell_wire[423];							inform_R[404][7] = r_cell_wire[424];							inform_R[468][7] = r_cell_wire[425];							inform_R[405][7] = r_cell_wire[426];							inform_R[469][7] = r_cell_wire[427];							inform_R[406][7] = r_cell_wire[428];							inform_R[470][7] = r_cell_wire[429];							inform_R[407][7] = r_cell_wire[430];							inform_R[471][7] = r_cell_wire[431];							inform_R[408][7] = r_cell_wire[432];							inform_R[472][7] = r_cell_wire[433];							inform_R[409][7] = r_cell_wire[434];							inform_R[473][7] = r_cell_wire[435];							inform_R[410][7] = r_cell_wire[436];							inform_R[474][7] = r_cell_wire[437];							inform_R[411][7] = r_cell_wire[438];							inform_R[475][7] = r_cell_wire[439];							inform_R[412][7] = r_cell_wire[440];							inform_R[476][7] = r_cell_wire[441];							inform_R[413][7] = r_cell_wire[442];							inform_R[477][7] = r_cell_wire[443];							inform_R[414][7] = r_cell_wire[444];							inform_R[478][7] = r_cell_wire[445];							inform_R[415][7] = r_cell_wire[446];							inform_R[479][7] = r_cell_wire[447];							inform_R[416][7] = r_cell_wire[448];							inform_R[480][7] = r_cell_wire[449];							inform_R[417][7] = r_cell_wire[450];							inform_R[481][7] = r_cell_wire[451];							inform_R[418][7] = r_cell_wire[452];							inform_R[482][7] = r_cell_wire[453];							inform_R[419][7] = r_cell_wire[454];							inform_R[483][7] = r_cell_wire[455];							inform_R[420][7] = r_cell_wire[456];							inform_R[484][7] = r_cell_wire[457];							inform_R[421][7] = r_cell_wire[458];							inform_R[485][7] = r_cell_wire[459];							inform_R[422][7] = r_cell_wire[460];							inform_R[486][7] = r_cell_wire[461];							inform_R[423][7] = r_cell_wire[462];							inform_R[487][7] = r_cell_wire[463];							inform_R[424][7] = r_cell_wire[464];							inform_R[488][7] = r_cell_wire[465];							inform_R[425][7] = r_cell_wire[466];							inform_R[489][7] = r_cell_wire[467];							inform_R[426][7] = r_cell_wire[468];							inform_R[490][7] = r_cell_wire[469];							inform_R[427][7] = r_cell_wire[470];							inform_R[491][7] = r_cell_wire[471];							inform_R[428][7] = r_cell_wire[472];							inform_R[492][7] = r_cell_wire[473];							inform_R[429][7] = r_cell_wire[474];							inform_R[493][7] = r_cell_wire[475];							inform_R[430][7] = r_cell_wire[476];							inform_R[494][7] = r_cell_wire[477];							inform_R[431][7] = r_cell_wire[478];							inform_R[495][7] = r_cell_wire[479];							inform_R[432][7] = r_cell_wire[480];							inform_R[496][7] = r_cell_wire[481];							inform_R[433][7] = r_cell_wire[482];							inform_R[497][7] = r_cell_wire[483];							inform_R[434][7] = r_cell_wire[484];							inform_R[498][7] = r_cell_wire[485];							inform_R[435][7] = r_cell_wire[486];							inform_R[499][7] = r_cell_wire[487];							inform_R[436][7] = r_cell_wire[488];							inform_R[500][7] = r_cell_wire[489];							inform_R[437][7] = r_cell_wire[490];							inform_R[501][7] = r_cell_wire[491];							inform_R[438][7] = r_cell_wire[492];							inform_R[502][7] = r_cell_wire[493];							inform_R[439][7] = r_cell_wire[494];							inform_R[503][7] = r_cell_wire[495];							inform_R[440][7] = r_cell_wire[496];							inform_R[504][7] = r_cell_wire[497];							inform_R[441][7] = r_cell_wire[498];							inform_R[505][7] = r_cell_wire[499];							inform_R[442][7] = r_cell_wire[500];							inform_R[506][7] = r_cell_wire[501];							inform_R[443][7] = r_cell_wire[502];							inform_R[507][7] = r_cell_wire[503];							inform_R[444][7] = r_cell_wire[504];							inform_R[508][7] = r_cell_wire[505];							inform_R[445][7] = r_cell_wire[506];							inform_R[509][7] = r_cell_wire[507];							inform_R[446][7] = r_cell_wire[508];							inform_R[510][7] = r_cell_wire[509];							inform_R[447][7] = r_cell_wire[510];							inform_R[511][7] = r_cell_wire[511];							inform_R[512][7] = r_cell_wire[512];							inform_R[576][7] = r_cell_wire[513];							inform_R[513][7] = r_cell_wire[514];							inform_R[577][7] = r_cell_wire[515];							inform_R[514][7] = r_cell_wire[516];							inform_R[578][7] = r_cell_wire[517];							inform_R[515][7] = r_cell_wire[518];							inform_R[579][7] = r_cell_wire[519];							inform_R[516][7] = r_cell_wire[520];							inform_R[580][7] = r_cell_wire[521];							inform_R[517][7] = r_cell_wire[522];							inform_R[581][7] = r_cell_wire[523];							inform_R[518][7] = r_cell_wire[524];							inform_R[582][7] = r_cell_wire[525];							inform_R[519][7] = r_cell_wire[526];							inform_R[583][7] = r_cell_wire[527];							inform_R[520][7] = r_cell_wire[528];							inform_R[584][7] = r_cell_wire[529];							inform_R[521][7] = r_cell_wire[530];							inform_R[585][7] = r_cell_wire[531];							inform_R[522][7] = r_cell_wire[532];							inform_R[586][7] = r_cell_wire[533];							inform_R[523][7] = r_cell_wire[534];							inform_R[587][7] = r_cell_wire[535];							inform_R[524][7] = r_cell_wire[536];							inform_R[588][7] = r_cell_wire[537];							inform_R[525][7] = r_cell_wire[538];							inform_R[589][7] = r_cell_wire[539];							inform_R[526][7] = r_cell_wire[540];							inform_R[590][7] = r_cell_wire[541];							inform_R[527][7] = r_cell_wire[542];							inform_R[591][7] = r_cell_wire[543];							inform_R[528][7] = r_cell_wire[544];							inform_R[592][7] = r_cell_wire[545];							inform_R[529][7] = r_cell_wire[546];							inform_R[593][7] = r_cell_wire[547];							inform_R[530][7] = r_cell_wire[548];							inform_R[594][7] = r_cell_wire[549];							inform_R[531][7] = r_cell_wire[550];							inform_R[595][7] = r_cell_wire[551];							inform_R[532][7] = r_cell_wire[552];							inform_R[596][7] = r_cell_wire[553];							inform_R[533][7] = r_cell_wire[554];							inform_R[597][7] = r_cell_wire[555];							inform_R[534][7] = r_cell_wire[556];							inform_R[598][7] = r_cell_wire[557];							inform_R[535][7] = r_cell_wire[558];							inform_R[599][7] = r_cell_wire[559];							inform_R[536][7] = r_cell_wire[560];							inform_R[600][7] = r_cell_wire[561];							inform_R[537][7] = r_cell_wire[562];							inform_R[601][7] = r_cell_wire[563];							inform_R[538][7] = r_cell_wire[564];							inform_R[602][7] = r_cell_wire[565];							inform_R[539][7] = r_cell_wire[566];							inform_R[603][7] = r_cell_wire[567];							inform_R[540][7] = r_cell_wire[568];							inform_R[604][7] = r_cell_wire[569];							inform_R[541][7] = r_cell_wire[570];							inform_R[605][7] = r_cell_wire[571];							inform_R[542][7] = r_cell_wire[572];							inform_R[606][7] = r_cell_wire[573];							inform_R[543][7] = r_cell_wire[574];							inform_R[607][7] = r_cell_wire[575];							inform_R[544][7] = r_cell_wire[576];							inform_R[608][7] = r_cell_wire[577];							inform_R[545][7] = r_cell_wire[578];							inform_R[609][7] = r_cell_wire[579];							inform_R[546][7] = r_cell_wire[580];							inform_R[610][7] = r_cell_wire[581];							inform_R[547][7] = r_cell_wire[582];							inform_R[611][7] = r_cell_wire[583];							inform_R[548][7] = r_cell_wire[584];							inform_R[612][7] = r_cell_wire[585];							inform_R[549][7] = r_cell_wire[586];							inform_R[613][7] = r_cell_wire[587];							inform_R[550][7] = r_cell_wire[588];							inform_R[614][7] = r_cell_wire[589];							inform_R[551][7] = r_cell_wire[590];							inform_R[615][7] = r_cell_wire[591];							inform_R[552][7] = r_cell_wire[592];							inform_R[616][7] = r_cell_wire[593];							inform_R[553][7] = r_cell_wire[594];							inform_R[617][7] = r_cell_wire[595];							inform_R[554][7] = r_cell_wire[596];							inform_R[618][7] = r_cell_wire[597];							inform_R[555][7] = r_cell_wire[598];							inform_R[619][7] = r_cell_wire[599];							inform_R[556][7] = r_cell_wire[600];							inform_R[620][7] = r_cell_wire[601];							inform_R[557][7] = r_cell_wire[602];							inform_R[621][7] = r_cell_wire[603];							inform_R[558][7] = r_cell_wire[604];							inform_R[622][7] = r_cell_wire[605];							inform_R[559][7] = r_cell_wire[606];							inform_R[623][7] = r_cell_wire[607];							inform_R[560][7] = r_cell_wire[608];							inform_R[624][7] = r_cell_wire[609];							inform_R[561][7] = r_cell_wire[610];							inform_R[625][7] = r_cell_wire[611];							inform_R[562][7] = r_cell_wire[612];							inform_R[626][7] = r_cell_wire[613];							inform_R[563][7] = r_cell_wire[614];							inform_R[627][7] = r_cell_wire[615];							inform_R[564][7] = r_cell_wire[616];							inform_R[628][7] = r_cell_wire[617];							inform_R[565][7] = r_cell_wire[618];							inform_R[629][7] = r_cell_wire[619];							inform_R[566][7] = r_cell_wire[620];							inform_R[630][7] = r_cell_wire[621];							inform_R[567][7] = r_cell_wire[622];							inform_R[631][7] = r_cell_wire[623];							inform_R[568][7] = r_cell_wire[624];							inform_R[632][7] = r_cell_wire[625];							inform_R[569][7] = r_cell_wire[626];							inform_R[633][7] = r_cell_wire[627];							inform_R[570][7] = r_cell_wire[628];							inform_R[634][7] = r_cell_wire[629];							inform_R[571][7] = r_cell_wire[630];							inform_R[635][7] = r_cell_wire[631];							inform_R[572][7] = r_cell_wire[632];							inform_R[636][7] = r_cell_wire[633];							inform_R[573][7] = r_cell_wire[634];							inform_R[637][7] = r_cell_wire[635];							inform_R[574][7] = r_cell_wire[636];							inform_R[638][7] = r_cell_wire[637];							inform_R[575][7] = r_cell_wire[638];							inform_R[639][7] = r_cell_wire[639];							inform_R[640][7] = r_cell_wire[640];							inform_R[704][7] = r_cell_wire[641];							inform_R[641][7] = r_cell_wire[642];							inform_R[705][7] = r_cell_wire[643];							inform_R[642][7] = r_cell_wire[644];							inform_R[706][7] = r_cell_wire[645];							inform_R[643][7] = r_cell_wire[646];							inform_R[707][7] = r_cell_wire[647];							inform_R[644][7] = r_cell_wire[648];							inform_R[708][7] = r_cell_wire[649];							inform_R[645][7] = r_cell_wire[650];							inform_R[709][7] = r_cell_wire[651];							inform_R[646][7] = r_cell_wire[652];							inform_R[710][7] = r_cell_wire[653];							inform_R[647][7] = r_cell_wire[654];							inform_R[711][7] = r_cell_wire[655];							inform_R[648][7] = r_cell_wire[656];							inform_R[712][7] = r_cell_wire[657];							inform_R[649][7] = r_cell_wire[658];							inform_R[713][7] = r_cell_wire[659];							inform_R[650][7] = r_cell_wire[660];							inform_R[714][7] = r_cell_wire[661];							inform_R[651][7] = r_cell_wire[662];							inform_R[715][7] = r_cell_wire[663];							inform_R[652][7] = r_cell_wire[664];							inform_R[716][7] = r_cell_wire[665];							inform_R[653][7] = r_cell_wire[666];							inform_R[717][7] = r_cell_wire[667];							inform_R[654][7] = r_cell_wire[668];							inform_R[718][7] = r_cell_wire[669];							inform_R[655][7] = r_cell_wire[670];							inform_R[719][7] = r_cell_wire[671];							inform_R[656][7] = r_cell_wire[672];							inform_R[720][7] = r_cell_wire[673];							inform_R[657][7] = r_cell_wire[674];							inform_R[721][7] = r_cell_wire[675];							inform_R[658][7] = r_cell_wire[676];							inform_R[722][7] = r_cell_wire[677];							inform_R[659][7] = r_cell_wire[678];							inform_R[723][7] = r_cell_wire[679];							inform_R[660][7] = r_cell_wire[680];							inform_R[724][7] = r_cell_wire[681];							inform_R[661][7] = r_cell_wire[682];							inform_R[725][7] = r_cell_wire[683];							inform_R[662][7] = r_cell_wire[684];							inform_R[726][7] = r_cell_wire[685];							inform_R[663][7] = r_cell_wire[686];							inform_R[727][7] = r_cell_wire[687];							inform_R[664][7] = r_cell_wire[688];							inform_R[728][7] = r_cell_wire[689];							inform_R[665][7] = r_cell_wire[690];							inform_R[729][7] = r_cell_wire[691];							inform_R[666][7] = r_cell_wire[692];							inform_R[730][7] = r_cell_wire[693];							inform_R[667][7] = r_cell_wire[694];							inform_R[731][7] = r_cell_wire[695];							inform_R[668][7] = r_cell_wire[696];							inform_R[732][7] = r_cell_wire[697];							inform_R[669][7] = r_cell_wire[698];							inform_R[733][7] = r_cell_wire[699];							inform_R[670][7] = r_cell_wire[700];							inform_R[734][7] = r_cell_wire[701];							inform_R[671][7] = r_cell_wire[702];							inform_R[735][7] = r_cell_wire[703];							inform_R[672][7] = r_cell_wire[704];							inform_R[736][7] = r_cell_wire[705];							inform_R[673][7] = r_cell_wire[706];							inform_R[737][7] = r_cell_wire[707];							inform_R[674][7] = r_cell_wire[708];							inform_R[738][7] = r_cell_wire[709];							inform_R[675][7] = r_cell_wire[710];							inform_R[739][7] = r_cell_wire[711];							inform_R[676][7] = r_cell_wire[712];							inform_R[740][7] = r_cell_wire[713];							inform_R[677][7] = r_cell_wire[714];							inform_R[741][7] = r_cell_wire[715];							inform_R[678][7] = r_cell_wire[716];							inform_R[742][7] = r_cell_wire[717];							inform_R[679][7] = r_cell_wire[718];							inform_R[743][7] = r_cell_wire[719];							inform_R[680][7] = r_cell_wire[720];							inform_R[744][7] = r_cell_wire[721];							inform_R[681][7] = r_cell_wire[722];							inform_R[745][7] = r_cell_wire[723];							inform_R[682][7] = r_cell_wire[724];							inform_R[746][7] = r_cell_wire[725];							inform_R[683][7] = r_cell_wire[726];							inform_R[747][7] = r_cell_wire[727];							inform_R[684][7] = r_cell_wire[728];							inform_R[748][7] = r_cell_wire[729];							inform_R[685][7] = r_cell_wire[730];							inform_R[749][7] = r_cell_wire[731];							inform_R[686][7] = r_cell_wire[732];							inform_R[750][7] = r_cell_wire[733];							inform_R[687][7] = r_cell_wire[734];							inform_R[751][7] = r_cell_wire[735];							inform_R[688][7] = r_cell_wire[736];							inform_R[752][7] = r_cell_wire[737];							inform_R[689][7] = r_cell_wire[738];							inform_R[753][7] = r_cell_wire[739];							inform_R[690][7] = r_cell_wire[740];							inform_R[754][7] = r_cell_wire[741];							inform_R[691][7] = r_cell_wire[742];							inform_R[755][7] = r_cell_wire[743];							inform_R[692][7] = r_cell_wire[744];							inform_R[756][7] = r_cell_wire[745];							inform_R[693][7] = r_cell_wire[746];							inform_R[757][7] = r_cell_wire[747];							inform_R[694][7] = r_cell_wire[748];							inform_R[758][7] = r_cell_wire[749];							inform_R[695][7] = r_cell_wire[750];							inform_R[759][7] = r_cell_wire[751];							inform_R[696][7] = r_cell_wire[752];							inform_R[760][7] = r_cell_wire[753];							inform_R[697][7] = r_cell_wire[754];							inform_R[761][7] = r_cell_wire[755];							inform_R[698][7] = r_cell_wire[756];							inform_R[762][7] = r_cell_wire[757];							inform_R[699][7] = r_cell_wire[758];							inform_R[763][7] = r_cell_wire[759];							inform_R[700][7] = r_cell_wire[760];							inform_R[764][7] = r_cell_wire[761];							inform_R[701][7] = r_cell_wire[762];							inform_R[765][7] = r_cell_wire[763];							inform_R[702][7] = r_cell_wire[764];							inform_R[766][7] = r_cell_wire[765];							inform_R[703][7] = r_cell_wire[766];							inform_R[767][7] = r_cell_wire[767];							inform_R[768][7] = r_cell_wire[768];							inform_R[832][7] = r_cell_wire[769];							inform_R[769][7] = r_cell_wire[770];							inform_R[833][7] = r_cell_wire[771];							inform_R[770][7] = r_cell_wire[772];							inform_R[834][7] = r_cell_wire[773];							inform_R[771][7] = r_cell_wire[774];							inform_R[835][7] = r_cell_wire[775];							inform_R[772][7] = r_cell_wire[776];							inform_R[836][7] = r_cell_wire[777];							inform_R[773][7] = r_cell_wire[778];							inform_R[837][7] = r_cell_wire[779];							inform_R[774][7] = r_cell_wire[780];							inform_R[838][7] = r_cell_wire[781];							inform_R[775][7] = r_cell_wire[782];							inform_R[839][7] = r_cell_wire[783];							inform_R[776][7] = r_cell_wire[784];							inform_R[840][7] = r_cell_wire[785];							inform_R[777][7] = r_cell_wire[786];							inform_R[841][7] = r_cell_wire[787];							inform_R[778][7] = r_cell_wire[788];							inform_R[842][7] = r_cell_wire[789];							inform_R[779][7] = r_cell_wire[790];							inform_R[843][7] = r_cell_wire[791];							inform_R[780][7] = r_cell_wire[792];							inform_R[844][7] = r_cell_wire[793];							inform_R[781][7] = r_cell_wire[794];							inform_R[845][7] = r_cell_wire[795];							inform_R[782][7] = r_cell_wire[796];							inform_R[846][7] = r_cell_wire[797];							inform_R[783][7] = r_cell_wire[798];							inform_R[847][7] = r_cell_wire[799];							inform_R[784][7] = r_cell_wire[800];							inform_R[848][7] = r_cell_wire[801];							inform_R[785][7] = r_cell_wire[802];							inform_R[849][7] = r_cell_wire[803];							inform_R[786][7] = r_cell_wire[804];							inform_R[850][7] = r_cell_wire[805];							inform_R[787][7] = r_cell_wire[806];							inform_R[851][7] = r_cell_wire[807];							inform_R[788][7] = r_cell_wire[808];							inform_R[852][7] = r_cell_wire[809];							inform_R[789][7] = r_cell_wire[810];							inform_R[853][7] = r_cell_wire[811];							inform_R[790][7] = r_cell_wire[812];							inform_R[854][7] = r_cell_wire[813];							inform_R[791][7] = r_cell_wire[814];							inform_R[855][7] = r_cell_wire[815];							inform_R[792][7] = r_cell_wire[816];							inform_R[856][7] = r_cell_wire[817];							inform_R[793][7] = r_cell_wire[818];							inform_R[857][7] = r_cell_wire[819];							inform_R[794][7] = r_cell_wire[820];							inform_R[858][7] = r_cell_wire[821];							inform_R[795][7] = r_cell_wire[822];							inform_R[859][7] = r_cell_wire[823];							inform_R[796][7] = r_cell_wire[824];							inform_R[860][7] = r_cell_wire[825];							inform_R[797][7] = r_cell_wire[826];							inform_R[861][7] = r_cell_wire[827];							inform_R[798][7] = r_cell_wire[828];							inform_R[862][7] = r_cell_wire[829];							inform_R[799][7] = r_cell_wire[830];							inform_R[863][7] = r_cell_wire[831];							inform_R[800][7] = r_cell_wire[832];							inform_R[864][7] = r_cell_wire[833];							inform_R[801][7] = r_cell_wire[834];							inform_R[865][7] = r_cell_wire[835];							inform_R[802][7] = r_cell_wire[836];							inform_R[866][7] = r_cell_wire[837];							inform_R[803][7] = r_cell_wire[838];							inform_R[867][7] = r_cell_wire[839];							inform_R[804][7] = r_cell_wire[840];							inform_R[868][7] = r_cell_wire[841];							inform_R[805][7] = r_cell_wire[842];							inform_R[869][7] = r_cell_wire[843];							inform_R[806][7] = r_cell_wire[844];							inform_R[870][7] = r_cell_wire[845];							inform_R[807][7] = r_cell_wire[846];							inform_R[871][7] = r_cell_wire[847];							inform_R[808][7] = r_cell_wire[848];							inform_R[872][7] = r_cell_wire[849];							inform_R[809][7] = r_cell_wire[850];							inform_R[873][7] = r_cell_wire[851];							inform_R[810][7] = r_cell_wire[852];							inform_R[874][7] = r_cell_wire[853];							inform_R[811][7] = r_cell_wire[854];							inform_R[875][7] = r_cell_wire[855];							inform_R[812][7] = r_cell_wire[856];							inform_R[876][7] = r_cell_wire[857];							inform_R[813][7] = r_cell_wire[858];							inform_R[877][7] = r_cell_wire[859];							inform_R[814][7] = r_cell_wire[860];							inform_R[878][7] = r_cell_wire[861];							inform_R[815][7] = r_cell_wire[862];							inform_R[879][7] = r_cell_wire[863];							inform_R[816][7] = r_cell_wire[864];							inform_R[880][7] = r_cell_wire[865];							inform_R[817][7] = r_cell_wire[866];							inform_R[881][7] = r_cell_wire[867];							inform_R[818][7] = r_cell_wire[868];							inform_R[882][7] = r_cell_wire[869];							inform_R[819][7] = r_cell_wire[870];							inform_R[883][7] = r_cell_wire[871];							inform_R[820][7] = r_cell_wire[872];							inform_R[884][7] = r_cell_wire[873];							inform_R[821][7] = r_cell_wire[874];							inform_R[885][7] = r_cell_wire[875];							inform_R[822][7] = r_cell_wire[876];							inform_R[886][7] = r_cell_wire[877];							inform_R[823][7] = r_cell_wire[878];							inform_R[887][7] = r_cell_wire[879];							inform_R[824][7] = r_cell_wire[880];							inform_R[888][7] = r_cell_wire[881];							inform_R[825][7] = r_cell_wire[882];							inform_R[889][7] = r_cell_wire[883];							inform_R[826][7] = r_cell_wire[884];							inform_R[890][7] = r_cell_wire[885];							inform_R[827][7] = r_cell_wire[886];							inform_R[891][7] = r_cell_wire[887];							inform_R[828][7] = r_cell_wire[888];							inform_R[892][7] = r_cell_wire[889];							inform_R[829][7] = r_cell_wire[890];							inform_R[893][7] = r_cell_wire[891];							inform_R[830][7] = r_cell_wire[892];							inform_R[894][7] = r_cell_wire[893];							inform_R[831][7] = r_cell_wire[894];							inform_R[895][7] = r_cell_wire[895];							inform_R[896][7] = r_cell_wire[896];							inform_R[960][7] = r_cell_wire[897];							inform_R[897][7] = r_cell_wire[898];							inform_R[961][7] = r_cell_wire[899];							inform_R[898][7] = r_cell_wire[900];							inform_R[962][7] = r_cell_wire[901];							inform_R[899][7] = r_cell_wire[902];							inform_R[963][7] = r_cell_wire[903];							inform_R[900][7] = r_cell_wire[904];							inform_R[964][7] = r_cell_wire[905];							inform_R[901][7] = r_cell_wire[906];							inform_R[965][7] = r_cell_wire[907];							inform_R[902][7] = r_cell_wire[908];							inform_R[966][7] = r_cell_wire[909];							inform_R[903][7] = r_cell_wire[910];							inform_R[967][7] = r_cell_wire[911];							inform_R[904][7] = r_cell_wire[912];							inform_R[968][7] = r_cell_wire[913];							inform_R[905][7] = r_cell_wire[914];							inform_R[969][7] = r_cell_wire[915];							inform_R[906][7] = r_cell_wire[916];							inform_R[970][7] = r_cell_wire[917];							inform_R[907][7] = r_cell_wire[918];							inform_R[971][7] = r_cell_wire[919];							inform_R[908][7] = r_cell_wire[920];							inform_R[972][7] = r_cell_wire[921];							inform_R[909][7] = r_cell_wire[922];							inform_R[973][7] = r_cell_wire[923];							inform_R[910][7] = r_cell_wire[924];							inform_R[974][7] = r_cell_wire[925];							inform_R[911][7] = r_cell_wire[926];							inform_R[975][7] = r_cell_wire[927];							inform_R[912][7] = r_cell_wire[928];							inform_R[976][7] = r_cell_wire[929];							inform_R[913][7] = r_cell_wire[930];							inform_R[977][7] = r_cell_wire[931];							inform_R[914][7] = r_cell_wire[932];							inform_R[978][7] = r_cell_wire[933];							inform_R[915][7] = r_cell_wire[934];							inform_R[979][7] = r_cell_wire[935];							inform_R[916][7] = r_cell_wire[936];							inform_R[980][7] = r_cell_wire[937];							inform_R[917][7] = r_cell_wire[938];							inform_R[981][7] = r_cell_wire[939];							inform_R[918][7] = r_cell_wire[940];							inform_R[982][7] = r_cell_wire[941];							inform_R[919][7] = r_cell_wire[942];							inform_R[983][7] = r_cell_wire[943];							inform_R[920][7] = r_cell_wire[944];							inform_R[984][7] = r_cell_wire[945];							inform_R[921][7] = r_cell_wire[946];							inform_R[985][7] = r_cell_wire[947];							inform_R[922][7] = r_cell_wire[948];							inform_R[986][7] = r_cell_wire[949];							inform_R[923][7] = r_cell_wire[950];							inform_R[987][7] = r_cell_wire[951];							inform_R[924][7] = r_cell_wire[952];							inform_R[988][7] = r_cell_wire[953];							inform_R[925][7] = r_cell_wire[954];							inform_R[989][7] = r_cell_wire[955];							inform_R[926][7] = r_cell_wire[956];							inform_R[990][7] = r_cell_wire[957];							inform_R[927][7] = r_cell_wire[958];							inform_R[991][7] = r_cell_wire[959];							inform_R[928][7] = r_cell_wire[960];							inform_R[992][7] = r_cell_wire[961];							inform_R[929][7] = r_cell_wire[962];							inform_R[993][7] = r_cell_wire[963];							inform_R[930][7] = r_cell_wire[964];							inform_R[994][7] = r_cell_wire[965];							inform_R[931][7] = r_cell_wire[966];							inform_R[995][7] = r_cell_wire[967];							inform_R[932][7] = r_cell_wire[968];							inform_R[996][7] = r_cell_wire[969];							inform_R[933][7] = r_cell_wire[970];							inform_R[997][7] = r_cell_wire[971];							inform_R[934][7] = r_cell_wire[972];							inform_R[998][7] = r_cell_wire[973];							inform_R[935][7] = r_cell_wire[974];							inform_R[999][7] = r_cell_wire[975];							inform_R[936][7] = r_cell_wire[976];							inform_R[1000][7] = r_cell_wire[977];							inform_R[937][7] = r_cell_wire[978];							inform_R[1001][7] = r_cell_wire[979];							inform_R[938][7] = r_cell_wire[980];							inform_R[1002][7] = r_cell_wire[981];							inform_R[939][7] = r_cell_wire[982];							inform_R[1003][7] = r_cell_wire[983];							inform_R[940][7] = r_cell_wire[984];							inform_R[1004][7] = r_cell_wire[985];							inform_R[941][7] = r_cell_wire[986];							inform_R[1005][7] = r_cell_wire[987];							inform_R[942][7] = r_cell_wire[988];							inform_R[1006][7] = r_cell_wire[989];							inform_R[943][7] = r_cell_wire[990];							inform_R[1007][7] = r_cell_wire[991];							inform_R[944][7] = r_cell_wire[992];							inform_R[1008][7] = r_cell_wire[993];							inform_R[945][7] = r_cell_wire[994];							inform_R[1009][7] = r_cell_wire[995];							inform_R[946][7] = r_cell_wire[996];							inform_R[1010][7] = r_cell_wire[997];							inform_R[947][7] = r_cell_wire[998];							inform_R[1011][7] = r_cell_wire[999];							inform_R[948][7] = r_cell_wire[1000];							inform_R[1012][7] = r_cell_wire[1001];							inform_R[949][7] = r_cell_wire[1002];							inform_R[1013][7] = r_cell_wire[1003];							inform_R[950][7] = r_cell_wire[1004];							inform_R[1014][7] = r_cell_wire[1005];							inform_R[951][7] = r_cell_wire[1006];							inform_R[1015][7] = r_cell_wire[1007];							inform_R[952][7] = r_cell_wire[1008];							inform_R[1016][7] = r_cell_wire[1009];							inform_R[953][7] = r_cell_wire[1010];							inform_R[1017][7] = r_cell_wire[1011];							inform_R[954][7] = r_cell_wire[1012];							inform_R[1018][7] = r_cell_wire[1013];							inform_R[955][7] = r_cell_wire[1014];							inform_R[1019][7] = r_cell_wire[1015];							inform_R[956][7] = r_cell_wire[1016];							inform_R[1020][7] = r_cell_wire[1017];							inform_R[957][7] = r_cell_wire[1018];							inform_R[1021][7] = r_cell_wire[1019];							inform_R[958][7] = r_cell_wire[1020];							inform_R[1022][7] = r_cell_wire[1021];							inform_R[959][7] = r_cell_wire[1022];							inform_R[1023][7] = r_cell_wire[1023];							inform_L[0][6] = l_cell_wire[0];							inform_L[64][6] = l_cell_wire[1];							inform_L[1][6] = l_cell_wire[2];							inform_L[65][6] = l_cell_wire[3];							inform_L[2][6] = l_cell_wire[4];							inform_L[66][6] = l_cell_wire[5];							inform_L[3][6] = l_cell_wire[6];							inform_L[67][6] = l_cell_wire[7];							inform_L[4][6] = l_cell_wire[8];							inform_L[68][6] = l_cell_wire[9];							inform_L[5][6] = l_cell_wire[10];							inform_L[69][6] = l_cell_wire[11];							inform_L[6][6] = l_cell_wire[12];							inform_L[70][6] = l_cell_wire[13];							inform_L[7][6] = l_cell_wire[14];							inform_L[71][6] = l_cell_wire[15];							inform_L[8][6] = l_cell_wire[16];							inform_L[72][6] = l_cell_wire[17];							inform_L[9][6] = l_cell_wire[18];							inform_L[73][6] = l_cell_wire[19];							inform_L[10][6] = l_cell_wire[20];							inform_L[74][6] = l_cell_wire[21];							inform_L[11][6] = l_cell_wire[22];							inform_L[75][6] = l_cell_wire[23];							inform_L[12][6] = l_cell_wire[24];							inform_L[76][6] = l_cell_wire[25];							inform_L[13][6] = l_cell_wire[26];							inform_L[77][6] = l_cell_wire[27];							inform_L[14][6] = l_cell_wire[28];							inform_L[78][6] = l_cell_wire[29];							inform_L[15][6] = l_cell_wire[30];							inform_L[79][6] = l_cell_wire[31];							inform_L[16][6] = l_cell_wire[32];							inform_L[80][6] = l_cell_wire[33];							inform_L[17][6] = l_cell_wire[34];							inform_L[81][6] = l_cell_wire[35];							inform_L[18][6] = l_cell_wire[36];							inform_L[82][6] = l_cell_wire[37];							inform_L[19][6] = l_cell_wire[38];							inform_L[83][6] = l_cell_wire[39];							inform_L[20][6] = l_cell_wire[40];							inform_L[84][6] = l_cell_wire[41];							inform_L[21][6] = l_cell_wire[42];							inform_L[85][6] = l_cell_wire[43];							inform_L[22][6] = l_cell_wire[44];							inform_L[86][6] = l_cell_wire[45];							inform_L[23][6] = l_cell_wire[46];							inform_L[87][6] = l_cell_wire[47];							inform_L[24][6] = l_cell_wire[48];							inform_L[88][6] = l_cell_wire[49];							inform_L[25][6] = l_cell_wire[50];							inform_L[89][6] = l_cell_wire[51];							inform_L[26][6] = l_cell_wire[52];							inform_L[90][6] = l_cell_wire[53];							inform_L[27][6] = l_cell_wire[54];							inform_L[91][6] = l_cell_wire[55];							inform_L[28][6] = l_cell_wire[56];							inform_L[92][6] = l_cell_wire[57];							inform_L[29][6] = l_cell_wire[58];							inform_L[93][6] = l_cell_wire[59];							inform_L[30][6] = l_cell_wire[60];							inform_L[94][6] = l_cell_wire[61];							inform_L[31][6] = l_cell_wire[62];							inform_L[95][6] = l_cell_wire[63];							inform_L[32][6] = l_cell_wire[64];							inform_L[96][6] = l_cell_wire[65];							inform_L[33][6] = l_cell_wire[66];							inform_L[97][6] = l_cell_wire[67];							inform_L[34][6] = l_cell_wire[68];							inform_L[98][6] = l_cell_wire[69];							inform_L[35][6] = l_cell_wire[70];							inform_L[99][6] = l_cell_wire[71];							inform_L[36][6] = l_cell_wire[72];							inform_L[100][6] = l_cell_wire[73];							inform_L[37][6] = l_cell_wire[74];							inform_L[101][6] = l_cell_wire[75];							inform_L[38][6] = l_cell_wire[76];							inform_L[102][6] = l_cell_wire[77];							inform_L[39][6] = l_cell_wire[78];							inform_L[103][6] = l_cell_wire[79];							inform_L[40][6] = l_cell_wire[80];							inform_L[104][6] = l_cell_wire[81];							inform_L[41][6] = l_cell_wire[82];							inform_L[105][6] = l_cell_wire[83];							inform_L[42][6] = l_cell_wire[84];							inform_L[106][6] = l_cell_wire[85];							inform_L[43][6] = l_cell_wire[86];							inform_L[107][6] = l_cell_wire[87];							inform_L[44][6] = l_cell_wire[88];							inform_L[108][6] = l_cell_wire[89];							inform_L[45][6] = l_cell_wire[90];							inform_L[109][6] = l_cell_wire[91];							inform_L[46][6] = l_cell_wire[92];							inform_L[110][6] = l_cell_wire[93];							inform_L[47][6] = l_cell_wire[94];							inform_L[111][6] = l_cell_wire[95];							inform_L[48][6] = l_cell_wire[96];							inform_L[112][6] = l_cell_wire[97];							inform_L[49][6] = l_cell_wire[98];							inform_L[113][6] = l_cell_wire[99];							inform_L[50][6] = l_cell_wire[100];							inform_L[114][6] = l_cell_wire[101];							inform_L[51][6] = l_cell_wire[102];							inform_L[115][6] = l_cell_wire[103];							inform_L[52][6] = l_cell_wire[104];							inform_L[116][6] = l_cell_wire[105];							inform_L[53][6] = l_cell_wire[106];							inform_L[117][6] = l_cell_wire[107];							inform_L[54][6] = l_cell_wire[108];							inform_L[118][6] = l_cell_wire[109];							inform_L[55][6] = l_cell_wire[110];							inform_L[119][6] = l_cell_wire[111];							inform_L[56][6] = l_cell_wire[112];							inform_L[120][6] = l_cell_wire[113];							inform_L[57][6] = l_cell_wire[114];							inform_L[121][6] = l_cell_wire[115];							inform_L[58][6] = l_cell_wire[116];							inform_L[122][6] = l_cell_wire[117];							inform_L[59][6] = l_cell_wire[118];							inform_L[123][6] = l_cell_wire[119];							inform_L[60][6] = l_cell_wire[120];							inform_L[124][6] = l_cell_wire[121];							inform_L[61][6] = l_cell_wire[122];							inform_L[125][6] = l_cell_wire[123];							inform_L[62][6] = l_cell_wire[124];							inform_L[126][6] = l_cell_wire[125];							inform_L[63][6] = l_cell_wire[126];							inform_L[127][6] = l_cell_wire[127];							inform_L[128][6] = l_cell_wire[128];							inform_L[192][6] = l_cell_wire[129];							inform_L[129][6] = l_cell_wire[130];							inform_L[193][6] = l_cell_wire[131];							inform_L[130][6] = l_cell_wire[132];							inform_L[194][6] = l_cell_wire[133];							inform_L[131][6] = l_cell_wire[134];							inform_L[195][6] = l_cell_wire[135];							inform_L[132][6] = l_cell_wire[136];							inform_L[196][6] = l_cell_wire[137];							inform_L[133][6] = l_cell_wire[138];							inform_L[197][6] = l_cell_wire[139];							inform_L[134][6] = l_cell_wire[140];							inform_L[198][6] = l_cell_wire[141];							inform_L[135][6] = l_cell_wire[142];							inform_L[199][6] = l_cell_wire[143];							inform_L[136][6] = l_cell_wire[144];							inform_L[200][6] = l_cell_wire[145];							inform_L[137][6] = l_cell_wire[146];							inform_L[201][6] = l_cell_wire[147];							inform_L[138][6] = l_cell_wire[148];							inform_L[202][6] = l_cell_wire[149];							inform_L[139][6] = l_cell_wire[150];							inform_L[203][6] = l_cell_wire[151];							inform_L[140][6] = l_cell_wire[152];							inform_L[204][6] = l_cell_wire[153];							inform_L[141][6] = l_cell_wire[154];							inform_L[205][6] = l_cell_wire[155];							inform_L[142][6] = l_cell_wire[156];							inform_L[206][6] = l_cell_wire[157];							inform_L[143][6] = l_cell_wire[158];							inform_L[207][6] = l_cell_wire[159];							inform_L[144][6] = l_cell_wire[160];							inform_L[208][6] = l_cell_wire[161];							inform_L[145][6] = l_cell_wire[162];							inform_L[209][6] = l_cell_wire[163];							inform_L[146][6] = l_cell_wire[164];							inform_L[210][6] = l_cell_wire[165];							inform_L[147][6] = l_cell_wire[166];							inform_L[211][6] = l_cell_wire[167];							inform_L[148][6] = l_cell_wire[168];							inform_L[212][6] = l_cell_wire[169];							inform_L[149][6] = l_cell_wire[170];							inform_L[213][6] = l_cell_wire[171];							inform_L[150][6] = l_cell_wire[172];							inform_L[214][6] = l_cell_wire[173];							inform_L[151][6] = l_cell_wire[174];							inform_L[215][6] = l_cell_wire[175];							inform_L[152][6] = l_cell_wire[176];							inform_L[216][6] = l_cell_wire[177];							inform_L[153][6] = l_cell_wire[178];							inform_L[217][6] = l_cell_wire[179];							inform_L[154][6] = l_cell_wire[180];							inform_L[218][6] = l_cell_wire[181];							inform_L[155][6] = l_cell_wire[182];							inform_L[219][6] = l_cell_wire[183];							inform_L[156][6] = l_cell_wire[184];							inform_L[220][6] = l_cell_wire[185];							inform_L[157][6] = l_cell_wire[186];							inform_L[221][6] = l_cell_wire[187];							inform_L[158][6] = l_cell_wire[188];							inform_L[222][6] = l_cell_wire[189];							inform_L[159][6] = l_cell_wire[190];							inform_L[223][6] = l_cell_wire[191];							inform_L[160][6] = l_cell_wire[192];							inform_L[224][6] = l_cell_wire[193];							inform_L[161][6] = l_cell_wire[194];							inform_L[225][6] = l_cell_wire[195];							inform_L[162][6] = l_cell_wire[196];							inform_L[226][6] = l_cell_wire[197];							inform_L[163][6] = l_cell_wire[198];							inform_L[227][6] = l_cell_wire[199];							inform_L[164][6] = l_cell_wire[200];							inform_L[228][6] = l_cell_wire[201];							inform_L[165][6] = l_cell_wire[202];							inform_L[229][6] = l_cell_wire[203];							inform_L[166][6] = l_cell_wire[204];							inform_L[230][6] = l_cell_wire[205];							inform_L[167][6] = l_cell_wire[206];							inform_L[231][6] = l_cell_wire[207];							inform_L[168][6] = l_cell_wire[208];							inform_L[232][6] = l_cell_wire[209];							inform_L[169][6] = l_cell_wire[210];							inform_L[233][6] = l_cell_wire[211];							inform_L[170][6] = l_cell_wire[212];							inform_L[234][6] = l_cell_wire[213];							inform_L[171][6] = l_cell_wire[214];							inform_L[235][6] = l_cell_wire[215];							inform_L[172][6] = l_cell_wire[216];							inform_L[236][6] = l_cell_wire[217];							inform_L[173][6] = l_cell_wire[218];							inform_L[237][6] = l_cell_wire[219];							inform_L[174][6] = l_cell_wire[220];							inform_L[238][6] = l_cell_wire[221];							inform_L[175][6] = l_cell_wire[222];							inform_L[239][6] = l_cell_wire[223];							inform_L[176][6] = l_cell_wire[224];							inform_L[240][6] = l_cell_wire[225];							inform_L[177][6] = l_cell_wire[226];							inform_L[241][6] = l_cell_wire[227];							inform_L[178][6] = l_cell_wire[228];							inform_L[242][6] = l_cell_wire[229];							inform_L[179][6] = l_cell_wire[230];							inform_L[243][6] = l_cell_wire[231];							inform_L[180][6] = l_cell_wire[232];							inform_L[244][6] = l_cell_wire[233];							inform_L[181][6] = l_cell_wire[234];							inform_L[245][6] = l_cell_wire[235];							inform_L[182][6] = l_cell_wire[236];							inform_L[246][6] = l_cell_wire[237];							inform_L[183][6] = l_cell_wire[238];							inform_L[247][6] = l_cell_wire[239];							inform_L[184][6] = l_cell_wire[240];							inform_L[248][6] = l_cell_wire[241];							inform_L[185][6] = l_cell_wire[242];							inform_L[249][6] = l_cell_wire[243];							inform_L[186][6] = l_cell_wire[244];							inform_L[250][6] = l_cell_wire[245];							inform_L[187][6] = l_cell_wire[246];							inform_L[251][6] = l_cell_wire[247];							inform_L[188][6] = l_cell_wire[248];							inform_L[252][6] = l_cell_wire[249];							inform_L[189][6] = l_cell_wire[250];							inform_L[253][6] = l_cell_wire[251];							inform_L[190][6] = l_cell_wire[252];							inform_L[254][6] = l_cell_wire[253];							inform_L[191][6] = l_cell_wire[254];							inform_L[255][6] = l_cell_wire[255];							inform_L[256][6] = l_cell_wire[256];							inform_L[320][6] = l_cell_wire[257];							inform_L[257][6] = l_cell_wire[258];							inform_L[321][6] = l_cell_wire[259];							inform_L[258][6] = l_cell_wire[260];							inform_L[322][6] = l_cell_wire[261];							inform_L[259][6] = l_cell_wire[262];							inform_L[323][6] = l_cell_wire[263];							inform_L[260][6] = l_cell_wire[264];							inform_L[324][6] = l_cell_wire[265];							inform_L[261][6] = l_cell_wire[266];							inform_L[325][6] = l_cell_wire[267];							inform_L[262][6] = l_cell_wire[268];							inform_L[326][6] = l_cell_wire[269];							inform_L[263][6] = l_cell_wire[270];							inform_L[327][6] = l_cell_wire[271];							inform_L[264][6] = l_cell_wire[272];							inform_L[328][6] = l_cell_wire[273];							inform_L[265][6] = l_cell_wire[274];							inform_L[329][6] = l_cell_wire[275];							inform_L[266][6] = l_cell_wire[276];							inform_L[330][6] = l_cell_wire[277];							inform_L[267][6] = l_cell_wire[278];							inform_L[331][6] = l_cell_wire[279];							inform_L[268][6] = l_cell_wire[280];							inform_L[332][6] = l_cell_wire[281];							inform_L[269][6] = l_cell_wire[282];							inform_L[333][6] = l_cell_wire[283];							inform_L[270][6] = l_cell_wire[284];							inform_L[334][6] = l_cell_wire[285];							inform_L[271][6] = l_cell_wire[286];							inform_L[335][6] = l_cell_wire[287];							inform_L[272][6] = l_cell_wire[288];							inform_L[336][6] = l_cell_wire[289];							inform_L[273][6] = l_cell_wire[290];							inform_L[337][6] = l_cell_wire[291];							inform_L[274][6] = l_cell_wire[292];							inform_L[338][6] = l_cell_wire[293];							inform_L[275][6] = l_cell_wire[294];							inform_L[339][6] = l_cell_wire[295];							inform_L[276][6] = l_cell_wire[296];							inform_L[340][6] = l_cell_wire[297];							inform_L[277][6] = l_cell_wire[298];							inform_L[341][6] = l_cell_wire[299];							inform_L[278][6] = l_cell_wire[300];							inform_L[342][6] = l_cell_wire[301];							inform_L[279][6] = l_cell_wire[302];							inform_L[343][6] = l_cell_wire[303];							inform_L[280][6] = l_cell_wire[304];							inform_L[344][6] = l_cell_wire[305];							inform_L[281][6] = l_cell_wire[306];							inform_L[345][6] = l_cell_wire[307];							inform_L[282][6] = l_cell_wire[308];							inform_L[346][6] = l_cell_wire[309];							inform_L[283][6] = l_cell_wire[310];							inform_L[347][6] = l_cell_wire[311];							inform_L[284][6] = l_cell_wire[312];							inform_L[348][6] = l_cell_wire[313];							inform_L[285][6] = l_cell_wire[314];							inform_L[349][6] = l_cell_wire[315];							inform_L[286][6] = l_cell_wire[316];							inform_L[350][6] = l_cell_wire[317];							inform_L[287][6] = l_cell_wire[318];							inform_L[351][6] = l_cell_wire[319];							inform_L[288][6] = l_cell_wire[320];							inform_L[352][6] = l_cell_wire[321];							inform_L[289][6] = l_cell_wire[322];							inform_L[353][6] = l_cell_wire[323];							inform_L[290][6] = l_cell_wire[324];							inform_L[354][6] = l_cell_wire[325];							inform_L[291][6] = l_cell_wire[326];							inform_L[355][6] = l_cell_wire[327];							inform_L[292][6] = l_cell_wire[328];							inform_L[356][6] = l_cell_wire[329];							inform_L[293][6] = l_cell_wire[330];							inform_L[357][6] = l_cell_wire[331];							inform_L[294][6] = l_cell_wire[332];							inform_L[358][6] = l_cell_wire[333];							inform_L[295][6] = l_cell_wire[334];							inform_L[359][6] = l_cell_wire[335];							inform_L[296][6] = l_cell_wire[336];							inform_L[360][6] = l_cell_wire[337];							inform_L[297][6] = l_cell_wire[338];							inform_L[361][6] = l_cell_wire[339];							inform_L[298][6] = l_cell_wire[340];							inform_L[362][6] = l_cell_wire[341];							inform_L[299][6] = l_cell_wire[342];							inform_L[363][6] = l_cell_wire[343];							inform_L[300][6] = l_cell_wire[344];							inform_L[364][6] = l_cell_wire[345];							inform_L[301][6] = l_cell_wire[346];							inform_L[365][6] = l_cell_wire[347];							inform_L[302][6] = l_cell_wire[348];							inform_L[366][6] = l_cell_wire[349];							inform_L[303][6] = l_cell_wire[350];							inform_L[367][6] = l_cell_wire[351];							inform_L[304][6] = l_cell_wire[352];							inform_L[368][6] = l_cell_wire[353];							inform_L[305][6] = l_cell_wire[354];							inform_L[369][6] = l_cell_wire[355];							inform_L[306][6] = l_cell_wire[356];							inform_L[370][6] = l_cell_wire[357];							inform_L[307][6] = l_cell_wire[358];							inform_L[371][6] = l_cell_wire[359];							inform_L[308][6] = l_cell_wire[360];							inform_L[372][6] = l_cell_wire[361];							inform_L[309][6] = l_cell_wire[362];							inform_L[373][6] = l_cell_wire[363];							inform_L[310][6] = l_cell_wire[364];							inform_L[374][6] = l_cell_wire[365];							inform_L[311][6] = l_cell_wire[366];							inform_L[375][6] = l_cell_wire[367];							inform_L[312][6] = l_cell_wire[368];							inform_L[376][6] = l_cell_wire[369];							inform_L[313][6] = l_cell_wire[370];							inform_L[377][6] = l_cell_wire[371];							inform_L[314][6] = l_cell_wire[372];							inform_L[378][6] = l_cell_wire[373];							inform_L[315][6] = l_cell_wire[374];							inform_L[379][6] = l_cell_wire[375];							inform_L[316][6] = l_cell_wire[376];							inform_L[380][6] = l_cell_wire[377];							inform_L[317][6] = l_cell_wire[378];							inform_L[381][6] = l_cell_wire[379];							inform_L[318][6] = l_cell_wire[380];							inform_L[382][6] = l_cell_wire[381];							inform_L[319][6] = l_cell_wire[382];							inform_L[383][6] = l_cell_wire[383];							inform_L[384][6] = l_cell_wire[384];							inform_L[448][6] = l_cell_wire[385];							inform_L[385][6] = l_cell_wire[386];							inform_L[449][6] = l_cell_wire[387];							inform_L[386][6] = l_cell_wire[388];							inform_L[450][6] = l_cell_wire[389];							inform_L[387][6] = l_cell_wire[390];							inform_L[451][6] = l_cell_wire[391];							inform_L[388][6] = l_cell_wire[392];							inform_L[452][6] = l_cell_wire[393];							inform_L[389][6] = l_cell_wire[394];							inform_L[453][6] = l_cell_wire[395];							inform_L[390][6] = l_cell_wire[396];							inform_L[454][6] = l_cell_wire[397];							inform_L[391][6] = l_cell_wire[398];							inform_L[455][6] = l_cell_wire[399];							inform_L[392][6] = l_cell_wire[400];							inform_L[456][6] = l_cell_wire[401];							inform_L[393][6] = l_cell_wire[402];							inform_L[457][6] = l_cell_wire[403];							inform_L[394][6] = l_cell_wire[404];							inform_L[458][6] = l_cell_wire[405];							inform_L[395][6] = l_cell_wire[406];							inform_L[459][6] = l_cell_wire[407];							inform_L[396][6] = l_cell_wire[408];							inform_L[460][6] = l_cell_wire[409];							inform_L[397][6] = l_cell_wire[410];							inform_L[461][6] = l_cell_wire[411];							inform_L[398][6] = l_cell_wire[412];							inform_L[462][6] = l_cell_wire[413];							inform_L[399][6] = l_cell_wire[414];							inform_L[463][6] = l_cell_wire[415];							inform_L[400][6] = l_cell_wire[416];							inform_L[464][6] = l_cell_wire[417];							inform_L[401][6] = l_cell_wire[418];							inform_L[465][6] = l_cell_wire[419];							inform_L[402][6] = l_cell_wire[420];							inform_L[466][6] = l_cell_wire[421];							inform_L[403][6] = l_cell_wire[422];							inform_L[467][6] = l_cell_wire[423];							inform_L[404][6] = l_cell_wire[424];							inform_L[468][6] = l_cell_wire[425];							inform_L[405][6] = l_cell_wire[426];							inform_L[469][6] = l_cell_wire[427];							inform_L[406][6] = l_cell_wire[428];							inform_L[470][6] = l_cell_wire[429];							inform_L[407][6] = l_cell_wire[430];							inform_L[471][6] = l_cell_wire[431];							inform_L[408][6] = l_cell_wire[432];							inform_L[472][6] = l_cell_wire[433];							inform_L[409][6] = l_cell_wire[434];							inform_L[473][6] = l_cell_wire[435];							inform_L[410][6] = l_cell_wire[436];							inform_L[474][6] = l_cell_wire[437];							inform_L[411][6] = l_cell_wire[438];							inform_L[475][6] = l_cell_wire[439];							inform_L[412][6] = l_cell_wire[440];							inform_L[476][6] = l_cell_wire[441];							inform_L[413][6] = l_cell_wire[442];							inform_L[477][6] = l_cell_wire[443];							inform_L[414][6] = l_cell_wire[444];							inform_L[478][6] = l_cell_wire[445];							inform_L[415][6] = l_cell_wire[446];							inform_L[479][6] = l_cell_wire[447];							inform_L[416][6] = l_cell_wire[448];							inform_L[480][6] = l_cell_wire[449];							inform_L[417][6] = l_cell_wire[450];							inform_L[481][6] = l_cell_wire[451];							inform_L[418][6] = l_cell_wire[452];							inform_L[482][6] = l_cell_wire[453];							inform_L[419][6] = l_cell_wire[454];							inform_L[483][6] = l_cell_wire[455];							inform_L[420][6] = l_cell_wire[456];							inform_L[484][6] = l_cell_wire[457];							inform_L[421][6] = l_cell_wire[458];							inform_L[485][6] = l_cell_wire[459];							inform_L[422][6] = l_cell_wire[460];							inform_L[486][6] = l_cell_wire[461];							inform_L[423][6] = l_cell_wire[462];							inform_L[487][6] = l_cell_wire[463];							inform_L[424][6] = l_cell_wire[464];							inform_L[488][6] = l_cell_wire[465];							inform_L[425][6] = l_cell_wire[466];							inform_L[489][6] = l_cell_wire[467];							inform_L[426][6] = l_cell_wire[468];							inform_L[490][6] = l_cell_wire[469];							inform_L[427][6] = l_cell_wire[470];							inform_L[491][6] = l_cell_wire[471];							inform_L[428][6] = l_cell_wire[472];							inform_L[492][6] = l_cell_wire[473];							inform_L[429][6] = l_cell_wire[474];							inform_L[493][6] = l_cell_wire[475];							inform_L[430][6] = l_cell_wire[476];							inform_L[494][6] = l_cell_wire[477];							inform_L[431][6] = l_cell_wire[478];							inform_L[495][6] = l_cell_wire[479];							inform_L[432][6] = l_cell_wire[480];							inform_L[496][6] = l_cell_wire[481];							inform_L[433][6] = l_cell_wire[482];							inform_L[497][6] = l_cell_wire[483];							inform_L[434][6] = l_cell_wire[484];							inform_L[498][6] = l_cell_wire[485];							inform_L[435][6] = l_cell_wire[486];							inform_L[499][6] = l_cell_wire[487];							inform_L[436][6] = l_cell_wire[488];							inform_L[500][6] = l_cell_wire[489];							inform_L[437][6] = l_cell_wire[490];							inform_L[501][6] = l_cell_wire[491];							inform_L[438][6] = l_cell_wire[492];							inform_L[502][6] = l_cell_wire[493];							inform_L[439][6] = l_cell_wire[494];							inform_L[503][6] = l_cell_wire[495];							inform_L[440][6] = l_cell_wire[496];							inform_L[504][6] = l_cell_wire[497];							inform_L[441][6] = l_cell_wire[498];							inform_L[505][6] = l_cell_wire[499];							inform_L[442][6] = l_cell_wire[500];							inform_L[506][6] = l_cell_wire[501];							inform_L[443][6] = l_cell_wire[502];							inform_L[507][6] = l_cell_wire[503];							inform_L[444][6] = l_cell_wire[504];							inform_L[508][6] = l_cell_wire[505];							inform_L[445][6] = l_cell_wire[506];							inform_L[509][6] = l_cell_wire[507];							inform_L[446][6] = l_cell_wire[508];							inform_L[510][6] = l_cell_wire[509];							inform_L[447][6] = l_cell_wire[510];							inform_L[511][6] = l_cell_wire[511];							inform_L[512][6] = l_cell_wire[512];							inform_L[576][6] = l_cell_wire[513];							inform_L[513][6] = l_cell_wire[514];							inform_L[577][6] = l_cell_wire[515];							inform_L[514][6] = l_cell_wire[516];							inform_L[578][6] = l_cell_wire[517];							inform_L[515][6] = l_cell_wire[518];							inform_L[579][6] = l_cell_wire[519];							inform_L[516][6] = l_cell_wire[520];							inform_L[580][6] = l_cell_wire[521];							inform_L[517][6] = l_cell_wire[522];							inform_L[581][6] = l_cell_wire[523];							inform_L[518][6] = l_cell_wire[524];							inform_L[582][6] = l_cell_wire[525];							inform_L[519][6] = l_cell_wire[526];							inform_L[583][6] = l_cell_wire[527];							inform_L[520][6] = l_cell_wire[528];							inform_L[584][6] = l_cell_wire[529];							inform_L[521][6] = l_cell_wire[530];							inform_L[585][6] = l_cell_wire[531];							inform_L[522][6] = l_cell_wire[532];							inform_L[586][6] = l_cell_wire[533];							inform_L[523][6] = l_cell_wire[534];							inform_L[587][6] = l_cell_wire[535];							inform_L[524][6] = l_cell_wire[536];							inform_L[588][6] = l_cell_wire[537];							inform_L[525][6] = l_cell_wire[538];							inform_L[589][6] = l_cell_wire[539];							inform_L[526][6] = l_cell_wire[540];							inform_L[590][6] = l_cell_wire[541];							inform_L[527][6] = l_cell_wire[542];							inform_L[591][6] = l_cell_wire[543];							inform_L[528][6] = l_cell_wire[544];							inform_L[592][6] = l_cell_wire[545];							inform_L[529][6] = l_cell_wire[546];							inform_L[593][6] = l_cell_wire[547];							inform_L[530][6] = l_cell_wire[548];							inform_L[594][6] = l_cell_wire[549];							inform_L[531][6] = l_cell_wire[550];							inform_L[595][6] = l_cell_wire[551];							inform_L[532][6] = l_cell_wire[552];							inform_L[596][6] = l_cell_wire[553];							inform_L[533][6] = l_cell_wire[554];							inform_L[597][6] = l_cell_wire[555];							inform_L[534][6] = l_cell_wire[556];							inform_L[598][6] = l_cell_wire[557];							inform_L[535][6] = l_cell_wire[558];							inform_L[599][6] = l_cell_wire[559];							inform_L[536][6] = l_cell_wire[560];							inform_L[600][6] = l_cell_wire[561];							inform_L[537][6] = l_cell_wire[562];							inform_L[601][6] = l_cell_wire[563];							inform_L[538][6] = l_cell_wire[564];							inform_L[602][6] = l_cell_wire[565];							inform_L[539][6] = l_cell_wire[566];							inform_L[603][6] = l_cell_wire[567];							inform_L[540][6] = l_cell_wire[568];							inform_L[604][6] = l_cell_wire[569];							inform_L[541][6] = l_cell_wire[570];							inform_L[605][6] = l_cell_wire[571];							inform_L[542][6] = l_cell_wire[572];							inform_L[606][6] = l_cell_wire[573];							inform_L[543][6] = l_cell_wire[574];							inform_L[607][6] = l_cell_wire[575];							inform_L[544][6] = l_cell_wire[576];							inform_L[608][6] = l_cell_wire[577];							inform_L[545][6] = l_cell_wire[578];							inform_L[609][6] = l_cell_wire[579];							inform_L[546][6] = l_cell_wire[580];							inform_L[610][6] = l_cell_wire[581];							inform_L[547][6] = l_cell_wire[582];							inform_L[611][6] = l_cell_wire[583];							inform_L[548][6] = l_cell_wire[584];							inform_L[612][6] = l_cell_wire[585];							inform_L[549][6] = l_cell_wire[586];							inform_L[613][6] = l_cell_wire[587];							inform_L[550][6] = l_cell_wire[588];							inform_L[614][6] = l_cell_wire[589];							inform_L[551][6] = l_cell_wire[590];							inform_L[615][6] = l_cell_wire[591];							inform_L[552][6] = l_cell_wire[592];							inform_L[616][6] = l_cell_wire[593];							inform_L[553][6] = l_cell_wire[594];							inform_L[617][6] = l_cell_wire[595];							inform_L[554][6] = l_cell_wire[596];							inform_L[618][6] = l_cell_wire[597];							inform_L[555][6] = l_cell_wire[598];							inform_L[619][6] = l_cell_wire[599];							inform_L[556][6] = l_cell_wire[600];							inform_L[620][6] = l_cell_wire[601];							inform_L[557][6] = l_cell_wire[602];							inform_L[621][6] = l_cell_wire[603];							inform_L[558][6] = l_cell_wire[604];							inform_L[622][6] = l_cell_wire[605];							inform_L[559][6] = l_cell_wire[606];							inform_L[623][6] = l_cell_wire[607];							inform_L[560][6] = l_cell_wire[608];							inform_L[624][6] = l_cell_wire[609];							inform_L[561][6] = l_cell_wire[610];							inform_L[625][6] = l_cell_wire[611];							inform_L[562][6] = l_cell_wire[612];							inform_L[626][6] = l_cell_wire[613];							inform_L[563][6] = l_cell_wire[614];							inform_L[627][6] = l_cell_wire[615];							inform_L[564][6] = l_cell_wire[616];							inform_L[628][6] = l_cell_wire[617];							inform_L[565][6] = l_cell_wire[618];							inform_L[629][6] = l_cell_wire[619];							inform_L[566][6] = l_cell_wire[620];							inform_L[630][6] = l_cell_wire[621];							inform_L[567][6] = l_cell_wire[622];							inform_L[631][6] = l_cell_wire[623];							inform_L[568][6] = l_cell_wire[624];							inform_L[632][6] = l_cell_wire[625];							inform_L[569][6] = l_cell_wire[626];							inform_L[633][6] = l_cell_wire[627];							inform_L[570][6] = l_cell_wire[628];							inform_L[634][6] = l_cell_wire[629];							inform_L[571][6] = l_cell_wire[630];							inform_L[635][6] = l_cell_wire[631];							inform_L[572][6] = l_cell_wire[632];							inform_L[636][6] = l_cell_wire[633];							inform_L[573][6] = l_cell_wire[634];							inform_L[637][6] = l_cell_wire[635];							inform_L[574][6] = l_cell_wire[636];							inform_L[638][6] = l_cell_wire[637];							inform_L[575][6] = l_cell_wire[638];							inform_L[639][6] = l_cell_wire[639];							inform_L[640][6] = l_cell_wire[640];							inform_L[704][6] = l_cell_wire[641];							inform_L[641][6] = l_cell_wire[642];							inform_L[705][6] = l_cell_wire[643];							inform_L[642][6] = l_cell_wire[644];							inform_L[706][6] = l_cell_wire[645];							inform_L[643][6] = l_cell_wire[646];							inform_L[707][6] = l_cell_wire[647];							inform_L[644][6] = l_cell_wire[648];							inform_L[708][6] = l_cell_wire[649];							inform_L[645][6] = l_cell_wire[650];							inform_L[709][6] = l_cell_wire[651];							inform_L[646][6] = l_cell_wire[652];							inform_L[710][6] = l_cell_wire[653];							inform_L[647][6] = l_cell_wire[654];							inform_L[711][6] = l_cell_wire[655];							inform_L[648][6] = l_cell_wire[656];							inform_L[712][6] = l_cell_wire[657];							inform_L[649][6] = l_cell_wire[658];							inform_L[713][6] = l_cell_wire[659];							inform_L[650][6] = l_cell_wire[660];							inform_L[714][6] = l_cell_wire[661];							inform_L[651][6] = l_cell_wire[662];							inform_L[715][6] = l_cell_wire[663];							inform_L[652][6] = l_cell_wire[664];							inform_L[716][6] = l_cell_wire[665];							inform_L[653][6] = l_cell_wire[666];							inform_L[717][6] = l_cell_wire[667];							inform_L[654][6] = l_cell_wire[668];							inform_L[718][6] = l_cell_wire[669];							inform_L[655][6] = l_cell_wire[670];							inform_L[719][6] = l_cell_wire[671];							inform_L[656][6] = l_cell_wire[672];							inform_L[720][6] = l_cell_wire[673];							inform_L[657][6] = l_cell_wire[674];							inform_L[721][6] = l_cell_wire[675];							inform_L[658][6] = l_cell_wire[676];							inform_L[722][6] = l_cell_wire[677];							inform_L[659][6] = l_cell_wire[678];							inform_L[723][6] = l_cell_wire[679];							inform_L[660][6] = l_cell_wire[680];							inform_L[724][6] = l_cell_wire[681];							inform_L[661][6] = l_cell_wire[682];							inform_L[725][6] = l_cell_wire[683];							inform_L[662][6] = l_cell_wire[684];							inform_L[726][6] = l_cell_wire[685];							inform_L[663][6] = l_cell_wire[686];							inform_L[727][6] = l_cell_wire[687];							inform_L[664][6] = l_cell_wire[688];							inform_L[728][6] = l_cell_wire[689];							inform_L[665][6] = l_cell_wire[690];							inform_L[729][6] = l_cell_wire[691];							inform_L[666][6] = l_cell_wire[692];							inform_L[730][6] = l_cell_wire[693];							inform_L[667][6] = l_cell_wire[694];							inform_L[731][6] = l_cell_wire[695];							inform_L[668][6] = l_cell_wire[696];							inform_L[732][6] = l_cell_wire[697];							inform_L[669][6] = l_cell_wire[698];							inform_L[733][6] = l_cell_wire[699];							inform_L[670][6] = l_cell_wire[700];							inform_L[734][6] = l_cell_wire[701];							inform_L[671][6] = l_cell_wire[702];							inform_L[735][6] = l_cell_wire[703];							inform_L[672][6] = l_cell_wire[704];							inform_L[736][6] = l_cell_wire[705];							inform_L[673][6] = l_cell_wire[706];							inform_L[737][6] = l_cell_wire[707];							inform_L[674][6] = l_cell_wire[708];							inform_L[738][6] = l_cell_wire[709];							inform_L[675][6] = l_cell_wire[710];							inform_L[739][6] = l_cell_wire[711];							inform_L[676][6] = l_cell_wire[712];							inform_L[740][6] = l_cell_wire[713];							inform_L[677][6] = l_cell_wire[714];							inform_L[741][6] = l_cell_wire[715];							inform_L[678][6] = l_cell_wire[716];							inform_L[742][6] = l_cell_wire[717];							inform_L[679][6] = l_cell_wire[718];							inform_L[743][6] = l_cell_wire[719];							inform_L[680][6] = l_cell_wire[720];							inform_L[744][6] = l_cell_wire[721];							inform_L[681][6] = l_cell_wire[722];							inform_L[745][6] = l_cell_wire[723];							inform_L[682][6] = l_cell_wire[724];							inform_L[746][6] = l_cell_wire[725];							inform_L[683][6] = l_cell_wire[726];							inform_L[747][6] = l_cell_wire[727];							inform_L[684][6] = l_cell_wire[728];							inform_L[748][6] = l_cell_wire[729];							inform_L[685][6] = l_cell_wire[730];							inform_L[749][6] = l_cell_wire[731];							inform_L[686][6] = l_cell_wire[732];							inform_L[750][6] = l_cell_wire[733];							inform_L[687][6] = l_cell_wire[734];							inform_L[751][6] = l_cell_wire[735];							inform_L[688][6] = l_cell_wire[736];							inform_L[752][6] = l_cell_wire[737];							inform_L[689][6] = l_cell_wire[738];							inform_L[753][6] = l_cell_wire[739];							inform_L[690][6] = l_cell_wire[740];							inform_L[754][6] = l_cell_wire[741];							inform_L[691][6] = l_cell_wire[742];							inform_L[755][6] = l_cell_wire[743];							inform_L[692][6] = l_cell_wire[744];							inform_L[756][6] = l_cell_wire[745];							inform_L[693][6] = l_cell_wire[746];							inform_L[757][6] = l_cell_wire[747];							inform_L[694][6] = l_cell_wire[748];							inform_L[758][6] = l_cell_wire[749];							inform_L[695][6] = l_cell_wire[750];							inform_L[759][6] = l_cell_wire[751];							inform_L[696][6] = l_cell_wire[752];							inform_L[760][6] = l_cell_wire[753];							inform_L[697][6] = l_cell_wire[754];							inform_L[761][6] = l_cell_wire[755];							inform_L[698][6] = l_cell_wire[756];							inform_L[762][6] = l_cell_wire[757];							inform_L[699][6] = l_cell_wire[758];							inform_L[763][6] = l_cell_wire[759];							inform_L[700][6] = l_cell_wire[760];							inform_L[764][6] = l_cell_wire[761];							inform_L[701][6] = l_cell_wire[762];							inform_L[765][6] = l_cell_wire[763];							inform_L[702][6] = l_cell_wire[764];							inform_L[766][6] = l_cell_wire[765];							inform_L[703][6] = l_cell_wire[766];							inform_L[767][6] = l_cell_wire[767];							inform_L[768][6] = l_cell_wire[768];							inform_L[832][6] = l_cell_wire[769];							inform_L[769][6] = l_cell_wire[770];							inform_L[833][6] = l_cell_wire[771];							inform_L[770][6] = l_cell_wire[772];							inform_L[834][6] = l_cell_wire[773];							inform_L[771][6] = l_cell_wire[774];							inform_L[835][6] = l_cell_wire[775];							inform_L[772][6] = l_cell_wire[776];							inform_L[836][6] = l_cell_wire[777];							inform_L[773][6] = l_cell_wire[778];							inform_L[837][6] = l_cell_wire[779];							inform_L[774][6] = l_cell_wire[780];							inform_L[838][6] = l_cell_wire[781];							inform_L[775][6] = l_cell_wire[782];							inform_L[839][6] = l_cell_wire[783];							inform_L[776][6] = l_cell_wire[784];							inform_L[840][6] = l_cell_wire[785];							inform_L[777][6] = l_cell_wire[786];							inform_L[841][6] = l_cell_wire[787];							inform_L[778][6] = l_cell_wire[788];							inform_L[842][6] = l_cell_wire[789];							inform_L[779][6] = l_cell_wire[790];							inform_L[843][6] = l_cell_wire[791];							inform_L[780][6] = l_cell_wire[792];							inform_L[844][6] = l_cell_wire[793];							inform_L[781][6] = l_cell_wire[794];							inform_L[845][6] = l_cell_wire[795];							inform_L[782][6] = l_cell_wire[796];							inform_L[846][6] = l_cell_wire[797];							inform_L[783][6] = l_cell_wire[798];							inform_L[847][6] = l_cell_wire[799];							inform_L[784][6] = l_cell_wire[800];							inform_L[848][6] = l_cell_wire[801];							inform_L[785][6] = l_cell_wire[802];							inform_L[849][6] = l_cell_wire[803];							inform_L[786][6] = l_cell_wire[804];							inform_L[850][6] = l_cell_wire[805];							inform_L[787][6] = l_cell_wire[806];							inform_L[851][6] = l_cell_wire[807];							inform_L[788][6] = l_cell_wire[808];							inform_L[852][6] = l_cell_wire[809];							inform_L[789][6] = l_cell_wire[810];							inform_L[853][6] = l_cell_wire[811];							inform_L[790][6] = l_cell_wire[812];							inform_L[854][6] = l_cell_wire[813];							inform_L[791][6] = l_cell_wire[814];							inform_L[855][6] = l_cell_wire[815];							inform_L[792][6] = l_cell_wire[816];							inform_L[856][6] = l_cell_wire[817];							inform_L[793][6] = l_cell_wire[818];							inform_L[857][6] = l_cell_wire[819];							inform_L[794][6] = l_cell_wire[820];							inform_L[858][6] = l_cell_wire[821];							inform_L[795][6] = l_cell_wire[822];							inform_L[859][6] = l_cell_wire[823];							inform_L[796][6] = l_cell_wire[824];							inform_L[860][6] = l_cell_wire[825];							inform_L[797][6] = l_cell_wire[826];							inform_L[861][6] = l_cell_wire[827];							inform_L[798][6] = l_cell_wire[828];							inform_L[862][6] = l_cell_wire[829];							inform_L[799][6] = l_cell_wire[830];							inform_L[863][6] = l_cell_wire[831];							inform_L[800][6] = l_cell_wire[832];							inform_L[864][6] = l_cell_wire[833];							inform_L[801][6] = l_cell_wire[834];							inform_L[865][6] = l_cell_wire[835];							inform_L[802][6] = l_cell_wire[836];							inform_L[866][6] = l_cell_wire[837];							inform_L[803][6] = l_cell_wire[838];							inform_L[867][6] = l_cell_wire[839];							inform_L[804][6] = l_cell_wire[840];							inform_L[868][6] = l_cell_wire[841];							inform_L[805][6] = l_cell_wire[842];							inform_L[869][6] = l_cell_wire[843];							inform_L[806][6] = l_cell_wire[844];							inform_L[870][6] = l_cell_wire[845];							inform_L[807][6] = l_cell_wire[846];							inform_L[871][6] = l_cell_wire[847];							inform_L[808][6] = l_cell_wire[848];							inform_L[872][6] = l_cell_wire[849];							inform_L[809][6] = l_cell_wire[850];							inform_L[873][6] = l_cell_wire[851];							inform_L[810][6] = l_cell_wire[852];							inform_L[874][6] = l_cell_wire[853];							inform_L[811][6] = l_cell_wire[854];							inform_L[875][6] = l_cell_wire[855];							inform_L[812][6] = l_cell_wire[856];							inform_L[876][6] = l_cell_wire[857];							inform_L[813][6] = l_cell_wire[858];							inform_L[877][6] = l_cell_wire[859];							inform_L[814][6] = l_cell_wire[860];							inform_L[878][6] = l_cell_wire[861];							inform_L[815][6] = l_cell_wire[862];							inform_L[879][6] = l_cell_wire[863];							inform_L[816][6] = l_cell_wire[864];							inform_L[880][6] = l_cell_wire[865];							inform_L[817][6] = l_cell_wire[866];							inform_L[881][6] = l_cell_wire[867];							inform_L[818][6] = l_cell_wire[868];							inform_L[882][6] = l_cell_wire[869];							inform_L[819][6] = l_cell_wire[870];							inform_L[883][6] = l_cell_wire[871];							inform_L[820][6] = l_cell_wire[872];							inform_L[884][6] = l_cell_wire[873];							inform_L[821][6] = l_cell_wire[874];							inform_L[885][6] = l_cell_wire[875];							inform_L[822][6] = l_cell_wire[876];							inform_L[886][6] = l_cell_wire[877];							inform_L[823][6] = l_cell_wire[878];							inform_L[887][6] = l_cell_wire[879];							inform_L[824][6] = l_cell_wire[880];							inform_L[888][6] = l_cell_wire[881];							inform_L[825][6] = l_cell_wire[882];							inform_L[889][6] = l_cell_wire[883];							inform_L[826][6] = l_cell_wire[884];							inform_L[890][6] = l_cell_wire[885];							inform_L[827][6] = l_cell_wire[886];							inform_L[891][6] = l_cell_wire[887];							inform_L[828][6] = l_cell_wire[888];							inform_L[892][6] = l_cell_wire[889];							inform_L[829][6] = l_cell_wire[890];							inform_L[893][6] = l_cell_wire[891];							inform_L[830][6] = l_cell_wire[892];							inform_L[894][6] = l_cell_wire[893];							inform_L[831][6] = l_cell_wire[894];							inform_L[895][6] = l_cell_wire[895];							inform_L[896][6] = l_cell_wire[896];							inform_L[960][6] = l_cell_wire[897];							inform_L[897][6] = l_cell_wire[898];							inform_L[961][6] = l_cell_wire[899];							inform_L[898][6] = l_cell_wire[900];							inform_L[962][6] = l_cell_wire[901];							inform_L[899][6] = l_cell_wire[902];							inform_L[963][6] = l_cell_wire[903];							inform_L[900][6] = l_cell_wire[904];							inform_L[964][6] = l_cell_wire[905];							inform_L[901][6] = l_cell_wire[906];							inform_L[965][6] = l_cell_wire[907];							inform_L[902][6] = l_cell_wire[908];							inform_L[966][6] = l_cell_wire[909];							inform_L[903][6] = l_cell_wire[910];							inform_L[967][6] = l_cell_wire[911];							inform_L[904][6] = l_cell_wire[912];							inform_L[968][6] = l_cell_wire[913];							inform_L[905][6] = l_cell_wire[914];							inform_L[969][6] = l_cell_wire[915];							inform_L[906][6] = l_cell_wire[916];							inform_L[970][6] = l_cell_wire[917];							inform_L[907][6] = l_cell_wire[918];							inform_L[971][6] = l_cell_wire[919];							inform_L[908][6] = l_cell_wire[920];							inform_L[972][6] = l_cell_wire[921];							inform_L[909][6] = l_cell_wire[922];							inform_L[973][6] = l_cell_wire[923];							inform_L[910][6] = l_cell_wire[924];							inform_L[974][6] = l_cell_wire[925];							inform_L[911][6] = l_cell_wire[926];							inform_L[975][6] = l_cell_wire[927];							inform_L[912][6] = l_cell_wire[928];							inform_L[976][6] = l_cell_wire[929];							inform_L[913][6] = l_cell_wire[930];							inform_L[977][6] = l_cell_wire[931];							inform_L[914][6] = l_cell_wire[932];							inform_L[978][6] = l_cell_wire[933];							inform_L[915][6] = l_cell_wire[934];							inform_L[979][6] = l_cell_wire[935];							inform_L[916][6] = l_cell_wire[936];							inform_L[980][6] = l_cell_wire[937];							inform_L[917][6] = l_cell_wire[938];							inform_L[981][6] = l_cell_wire[939];							inform_L[918][6] = l_cell_wire[940];							inform_L[982][6] = l_cell_wire[941];							inform_L[919][6] = l_cell_wire[942];							inform_L[983][6] = l_cell_wire[943];							inform_L[920][6] = l_cell_wire[944];							inform_L[984][6] = l_cell_wire[945];							inform_L[921][6] = l_cell_wire[946];							inform_L[985][6] = l_cell_wire[947];							inform_L[922][6] = l_cell_wire[948];							inform_L[986][6] = l_cell_wire[949];							inform_L[923][6] = l_cell_wire[950];							inform_L[987][6] = l_cell_wire[951];							inform_L[924][6] = l_cell_wire[952];							inform_L[988][6] = l_cell_wire[953];							inform_L[925][6] = l_cell_wire[954];							inform_L[989][6] = l_cell_wire[955];							inform_L[926][6] = l_cell_wire[956];							inform_L[990][6] = l_cell_wire[957];							inform_L[927][6] = l_cell_wire[958];							inform_L[991][6] = l_cell_wire[959];							inform_L[928][6] = l_cell_wire[960];							inform_L[992][6] = l_cell_wire[961];							inform_L[929][6] = l_cell_wire[962];							inform_L[993][6] = l_cell_wire[963];							inform_L[930][6] = l_cell_wire[964];							inform_L[994][6] = l_cell_wire[965];							inform_L[931][6] = l_cell_wire[966];							inform_L[995][6] = l_cell_wire[967];							inform_L[932][6] = l_cell_wire[968];							inform_L[996][6] = l_cell_wire[969];							inform_L[933][6] = l_cell_wire[970];							inform_L[997][6] = l_cell_wire[971];							inform_L[934][6] = l_cell_wire[972];							inform_L[998][6] = l_cell_wire[973];							inform_L[935][6] = l_cell_wire[974];							inform_L[999][6] = l_cell_wire[975];							inform_L[936][6] = l_cell_wire[976];							inform_L[1000][6] = l_cell_wire[977];							inform_L[937][6] = l_cell_wire[978];							inform_L[1001][6] = l_cell_wire[979];							inform_L[938][6] = l_cell_wire[980];							inform_L[1002][6] = l_cell_wire[981];							inform_L[939][6] = l_cell_wire[982];							inform_L[1003][6] = l_cell_wire[983];							inform_L[940][6] = l_cell_wire[984];							inform_L[1004][6] = l_cell_wire[985];							inform_L[941][6] = l_cell_wire[986];							inform_L[1005][6] = l_cell_wire[987];							inform_L[942][6] = l_cell_wire[988];							inform_L[1006][6] = l_cell_wire[989];							inform_L[943][6] = l_cell_wire[990];							inform_L[1007][6] = l_cell_wire[991];							inform_L[944][6] = l_cell_wire[992];							inform_L[1008][6] = l_cell_wire[993];							inform_L[945][6] = l_cell_wire[994];							inform_L[1009][6] = l_cell_wire[995];							inform_L[946][6] = l_cell_wire[996];							inform_L[1010][6] = l_cell_wire[997];							inform_L[947][6] = l_cell_wire[998];							inform_L[1011][6] = l_cell_wire[999];							inform_L[948][6] = l_cell_wire[1000];							inform_L[1012][6] = l_cell_wire[1001];							inform_L[949][6] = l_cell_wire[1002];							inform_L[1013][6] = l_cell_wire[1003];							inform_L[950][6] = l_cell_wire[1004];							inform_L[1014][6] = l_cell_wire[1005];							inform_L[951][6] = l_cell_wire[1006];							inform_L[1015][6] = l_cell_wire[1007];							inform_L[952][6] = l_cell_wire[1008];							inform_L[1016][6] = l_cell_wire[1009];							inform_L[953][6] = l_cell_wire[1010];							inform_L[1017][6] = l_cell_wire[1011];							inform_L[954][6] = l_cell_wire[1012];							inform_L[1018][6] = l_cell_wire[1013];							inform_L[955][6] = l_cell_wire[1014];							inform_L[1019][6] = l_cell_wire[1015];							inform_L[956][6] = l_cell_wire[1016];							inform_L[1020][6] = l_cell_wire[1017];							inform_L[957][6] = l_cell_wire[1018];							inform_L[1021][6] = l_cell_wire[1019];							inform_L[958][6] = l_cell_wire[1020];							inform_L[1022][6] = l_cell_wire[1021];							inform_L[959][6] = l_cell_wire[1022];							inform_L[1023][6] = l_cell_wire[1023];						end
						8:						begin							inform_R[0][8] = r_cell_wire[0];							inform_R[128][8] = r_cell_wire[1];							inform_R[1][8] = r_cell_wire[2];							inform_R[129][8] = r_cell_wire[3];							inform_R[2][8] = r_cell_wire[4];							inform_R[130][8] = r_cell_wire[5];							inform_R[3][8] = r_cell_wire[6];							inform_R[131][8] = r_cell_wire[7];							inform_R[4][8] = r_cell_wire[8];							inform_R[132][8] = r_cell_wire[9];							inform_R[5][8] = r_cell_wire[10];							inform_R[133][8] = r_cell_wire[11];							inform_R[6][8] = r_cell_wire[12];							inform_R[134][8] = r_cell_wire[13];							inform_R[7][8] = r_cell_wire[14];							inform_R[135][8] = r_cell_wire[15];							inform_R[8][8] = r_cell_wire[16];							inform_R[136][8] = r_cell_wire[17];							inform_R[9][8] = r_cell_wire[18];							inform_R[137][8] = r_cell_wire[19];							inform_R[10][8] = r_cell_wire[20];							inform_R[138][8] = r_cell_wire[21];							inform_R[11][8] = r_cell_wire[22];							inform_R[139][8] = r_cell_wire[23];							inform_R[12][8] = r_cell_wire[24];							inform_R[140][8] = r_cell_wire[25];							inform_R[13][8] = r_cell_wire[26];							inform_R[141][8] = r_cell_wire[27];							inform_R[14][8] = r_cell_wire[28];							inform_R[142][8] = r_cell_wire[29];							inform_R[15][8] = r_cell_wire[30];							inform_R[143][8] = r_cell_wire[31];							inform_R[16][8] = r_cell_wire[32];							inform_R[144][8] = r_cell_wire[33];							inform_R[17][8] = r_cell_wire[34];							inform_R[145][8] = r_cell_wire[35];							inform_R[18][8] = r_cell_wire[36];							inform_R[146][8] = r_cell_wire[37];							inform_R[19][8] = r_cell_wire[38];							inform_R[147][8] = r_cell_wire[39];							inform_R[20][8] = r_cell_wire[40];							inform_R[148][8] = r_cell_wire[41];							inform_R[21][8] = r_cell_wire[42];							inform_R[149][8] = r_cell_wire[43];							inform_R[22][8] = r_cell_wire[44];							inform_R[150][8] = r_cell_wire[45];							inform_R[23][8] = r_cell_wire[46];							inform_R[151][8] = r_cell_wire[47];							inform_R[24][8] = r_cell_wire[48];							inform_R[152][8] = r_cell_wire[49];							inform_R[25][8] = r_cell_wire[50];							inform_R[153][8] = r_cell_wire[51];							inform_R[26][8] = r_cell_wire[52];							inform_R[154][8] = r_cell_wire[53];							inform_R[27][8] = r_cell_wire[54];							inform_R[155][8] = r_cell_wire[55];							inform_R[28][8] = r_cell_wire[56];							inform_R[156][8] = r_cell_wire[57];							inform_R[29][8] = r_cell_wire[58];							inform_R[157][8] = r_cell_wire[59];							inform_R[30][8] = r_cell_wire[60];							inform_R[158][8] = r_cell_wire[61];							inform_R[31][8] = r_cell_wire[62];							inform_R[159][8] = r_cell_wire[63];							inform_R[32][8] = r_cell_wire[64];							inform_R[160][8] = r_cell_wire[65];							inform_R[33][8] = r_cell_wire[66];							inform_R[161][8] = r_cell_wire[67];							inform_R[34][8] = r_cell_wire[68];							inform_R[162][8] = r_cell_wire[69];							inform_R[35][8] = r_cell_wire[70];							inform_R[163][8] = r_cell_wire[71];							inform_R[36][8] = r_cell_wire[72];							inform_R[164][8] = r_cell_wire[73];							inform_R[37][8] = r_cell_wire[74];							inform_R[165][8] = r_cell_wire[75];							inform_R[38][8] = r_cell_wire[76];							inform_R[166][8] = r_cell_wire[77];							inform_R[39][8] = r_cell_wire[78];							inform_R[167][8] = r_cell_wire[79];							inform_R[40][8] = r_cell_wire[80];							inform_R[168][8] = r_cell_wire[81];							inform_R[41][8] = r_cell_wire[82];							inform_R[169][8] = r_cell_wire[83];							inform_R[42][8] = r_cell_wire[84];							inform_R[170][8] = r_cell_wire[85];							inform_R[43][8] = r_cell_wire[86];							inform_R[171][8] = r_cell_wire[87];							inform_R[44][8] = r_cell_wire[88];							inform_R[172][8] = r_cell_wire[89];							inform_R[45][8] = r_cell_wire[90];							inform_R[173][8] = r_cell_wire[91];							inform_R[46][8] = r_cell_wire[92];							inform_R[174][8] = r_cell_wire[93];							inform_R[47][8] = r_cell_wire[94];							inform_R[175][8] = r_cell_wire[95];							inform_R[48][8] = r_cell_wire[96];							inform_R[176][8] = r_cell_wire[97];							inform_R[49][8] = r_cell_wire[98];							inform_R[177][8] = r_cell_wire[99];							inform_R[50][8] = r_cell_wire[100];							inform_R[178][8] = r_cell_wire[101];							inform_R[51][8] = r_cell_wire[102];							inform_R[179][8] = r_cell_wire[103];							inform_R[52][8] = r_cell_wire[104];							inform_R[180][8] = r_cell_wire[105];							inform_R[53][8] = r_cell_wire[106];							inform_R[181][8] = r_cell_wire[107];							inform_R[54][8] = r_cell_wire[108];							inform_R[182][8] = r_cell_wire[109];							inform_R[55][8] = r_cell_wire[110];							inform_R[183][8] = r_cell_wire[111];							inform_R[56][8] = r_cell_wire[112];							inform_R[184][8] = r_cell_wire[113];							inform_R[57][8] = r_cell_wire[114];							inform_R[185][8] = r_cell_wire[115];							inform_R[58][8] = r_cell_wire[116];							inform_R[186][8] = r_cell_wire[117];							inform_R[59][8] = r_cell_wire[118];							inform_R[187][8] = r_cell_wire[119];							inform_R[60][8] = r_cell_wire[120];							inform_R[188][8] = r_cell_wire[121];							inform_R[61][8] = r_cell_wire[122];							inform_R[189][8] = r_cell_wire[123];							inform_R[62][8] = r_cell_wire[124];							inform_R[190][8] = r_cell_wire[125];							inform_R[63][8] = r_cell_wire[126];							inform_R[191][8] = r_cell_wire[127];							inform_R[64][8] = r_cell_wire[128];							inform_R[192][8] = r_cell_wire[129];							inform_R[65][8] = r_cell_wire[130];							inform_R[193][8] = r_cell_wire[131];							inform_R[66][8] = r_cell_wire[132];							inform_R[194][8] = r_cell_wire[133];							inform_R[67][8] = r_cell_wire[134];							inform_R[195][8] = r_cell_wire[135];							inform_R[68][8] = r_cell_wire[136];							inform_R[196][8] = r_cell_wire[137];							inform_R[69][8] = r_cell_wire[138];							inform_R[197][8] = r_cell_wire[139];							inform_R[70][8] = r_cell_wire[140];							inform_R[198][8] = r_cell_wire[141];							inform_R[71][8] = r_cell_wire[142];							inform_R[199][8] = r_cell_wire[143];							inform_R[72][8] = r_cell_wire[144];							inform_R[200][8] = r_cell_wire[145];							inform_R[73][8] = r_cell_wire[146];							inform_R[201][8] = r_cell_wire[147];							inform_R[74][8] = r_cell_wire[148];							inform_R[202][8] = r_cell_wire[149];							inform_R[75][8] = r_cell_wire[150];							inform_R[203][8] = r_cell_wire[151];							inform_R[76][8] = r_cell_wire[152];							inform_R[204][8] = r_cell_wire[153];							inform_R[77][8] = r_cell_wire[154];							inform_R[205][8] = r_cell_wire[155];							inform_R[78][8] = r_cell_wire[156];							inform_R[206][8] = r_cell_wire[157];							inform_R[79][8] = r_cell_wire[158];							inform_R[207][8] = r_cell_wire[159];							inform_R[80][8] = r_cell_wire[160];							inform_R[208][8] = r_cell_wire[161];							inform_R[81][8] = r_cell_wire[162];							inform_R[209][8] = r_cell_wire[163];							inform_R[82][8] = r_cell_wire[164];							inform_R[210][8] = r_cell_wire[165];							inform_R[83][8] = r_cell_wire[166];							inform_R[211][8] = r_cell_wire[167];							inform_R[84][8] = r_cell_wire[168];							inform_R[212][8] = r_cell_wire[169];							inform_R[85][8] = r_cell_wire[170];							inform_R[213][8] = r_cell_wire[171];							inform_R[86][8] = r_cell_wire[172];							inform_R[214][8] = r_cell_wire[173];							inform_R[87][8] = r_cell_wire[174];							inform_R[215][8] = r_cell_wire[175];							inform_R[88][8] = r_cell_wire[176];							inform_R[216][8] = r_cell_wire[177];							inform_R[89][8] = r_cell_wire[178];							inform_R[217][8] = r_cell_wire[179];							inform_R[90][8] = r_cell_wire[180];							inform_R[218][8] = r_cell_wire[181];							inform_R[91][8] = r_cell_wire[182];							inform_R[219][8] = r_cell_wire[183];							inform_R[92][8] = r_cell_wire[184];							inform_R[220][8] = r_cell_wire[185];							inform_R[93][8] = r_cell_wire[186];							inform_R[221][8] = r_cell_wire[187];							inform_R[94][8] = r_cell_wire[188];							inform_R[222][8] = r_cell_wire[189];							inform_R[95][8] = r_cell_wire[190];							inform_R[223][8] = r_cell_wire[191];							inform_R[96][8] = r_cell_wire[192];							inform_R[224][8] = r_cell_wire[193];							inform_R[97][8] = r_cell_wire[194];							inform_R[225][8] = r_cell_wire[195];							inform_R[98][8] = r_cell_wire[196];							inform_R[226][8] = r_cell_wire[197];							inform_R[99][8] = r_cell_wire[198];							inform_R[227][8] = r_cell_wire[199];							inform_R[100][8] = r_cell_wire[200];							inform_R[228][8] = r_cell_wire[201];							inform_R[101][8] = r_cell_wire[202];							inform_R[229][8] = r_cell_wire[203];							inform_R[102][8] = r_cell_wire[204];							inform_R[230][8] = r_cell_wire[205];							inform_R[103][8] = r_cell_wire[206];							inform_R[231][8] = r_cell_wire[207];							inform_R[104][8] = r_cell_wire[208];							inform_R[232][8] = r_cell_wire[209];							inform_R[105][8] = r_cell_wire[210];							inform_R[233][8] = r_cell_wire[211];							inform_R[106][8] = r_cell_wire[212];							inform_R[234][8] = r_cell_wire[213];							inform_R[107][8] = r_cell_wire[214];							inform_R[235][8] = r_cell_wire[215];							inform_R[108][8] = r_cell_wire[216];							inform_R[236][8] = r_cell_wire[217];							inform_R[109][8] = r_cell_wire[218];							inform_R[237][8] = r_cell_wire[219];							inform_R[110][8] = r_cell_wire[220];							inform_R[238][8] = r_cell_wire[221];							inform_R[111][8] = r_cell_wire[222];							inform_R[239][8] = r_cell_wire[223];							inform_R[112][8] = r_cell_wire[224];							inform_R[240][8] = r_cell_wire[225];							inform_R[113][8] = r_cell_wire[226];							inform_R[241][8] = r_cell_wire[227];							inform_R[114][8] = r_cell_wire[228];							inform_R[242][8] = r_cell_wire[229];							inform_R[115][8] = r_cell_wire[230];							inform_R[243][8] = r_cell_wire[231];							inform_R[116][8] = r_cell_wire[232];							inform_R[244][8] = r_cell_wire[233];							inform_R[117][8] = r_cell_wire[234];							inform_R[245][8] = r_cell_wire[235];							inform_R[118][8] = r_cell_wire[236];							inform_R[246][8] = r_cell_wire[237];							inform_R[119][8] = r_cell_wire[238];							inform_R[247][8] = r_cell_wire[239];							inform_R[120][8] = r_cell_wire[240];							inform_R[248][8] = r_cell_wire[241];							inform_R[121][8] = r_cell_wire[242];							inform_R[249][8] = r_cell_wire[243];							inform_R[122][8] = r_cell_wire[244];							inform_R[250][8] = r_cell_wire[245];							inform_R[123][8] = r_cell_wire[246];							inform_R[251][8] = r_cell_wire[247];							inform_R[124][8] = r_cell_wire[248];							inform_R[252][8] = r_cell_wire[249];							inform_R[125][8] = r_cell_wire[250];							inform_R[253][8] = r_cell_wire[251];							inform_R[126][8] = r_cell_wire[252];							inform_R[254][8] = r_cell_wire[253];							inform_R[127][8] = r_cell_wire[254];							inform_R[255][8] = r_cell_wire[255];							inform_R[256][8] = r_cell_wire[256];							inform_R[384][8] = r_cell_wire[257];							inform_R[257][8] = r_cell_wire[258];							inform_R[385][8] = r_cell_wire[259];							inform_R[258][8] = r_cell_wire[260];							inform_R[386][8] = r_cell_wire[261];							inform_R[259][8] = r_cell_wire[262];							inform_R[387][8] = r_cell_wire[263];							inform_R[260][8] = r_cell_wire[264];							inform_R[388][8] = r_cell_wire[265];							inform_R[261][8] = r_cell_wire[266];							inform_R[389][8] = r_cell_wire[267];							inform_R[262][8] = r_cell_wire[268];							inform_R[390][8] = r_cell_wire[269];							inform_R[263][8] = r_cell_wire[270];							inform_R[391][8] = r_cell_wire[271];							inform_R[264][8] = r_cell_wire[272];							inform_R[392][8] = r_cell_wire[273];							inform_R[265][8] = r_cell_wire[274];							inform_R[393][8] = r_cell_wire[275];							inform_R[266][8] = r_cell_wire[276];							inform_R[394][8] = r_cell_wire[277];							inform_R[267][8] = r_cell_wire[278];							inform_R[395][8] = r_cell_wire[279];							inform_R[268][8] = r_cell_wire[280];							inform_R[396][8] = r_cell_wire[281];							inform_R[269][8] = r_cell_wire[282];							inform_R[397][8] = r_cell_wire[283];							inform_R[270][8] = r_cell_wire[284];							inform_R[398][8] = r_cell_wire[285];							inform_R[271][8] = r_cell_wire[286];							inform_R[399][8] = r_cell_wire[287];							inform_R[272][8] = r_cell_wire[288];							inform_R[400][8] = r_cell_wire[289];							inform_R[273][8] = r_cell_wire[290];							inform_R[401][8] = r_cell_wire[291];							inform_R[274][8] = r_cell_wire[292];							inform_R[402][8] = r_cell_wire[293];							inform_R[275][8] = r_cell_wire[294];							inform_R[403][8] = r_cell_wire[295];							inform_R[276][8] = r_cell_wire[296];							inform_R[404][8] = r_cell_wire[297];							inform_R[277][8] = r_cell_wire[298];							inform_R[405][8] = r_cell_wire[299];							inform_R[278][8] = r_cell_wire[300];							inform_R[406][8] = r_cell_wire[301];							inform_R[279][8] = r_cell_wire[302];							inform_R[407][8] = r_cell_wire[303];							inform_R[280][8] = r_cell_wire[304];							inform_R[408][8] = r_cell_wire[305];							inform_R[281][8] = r_cell_wire[306];							inform_R[409][8] = r_cell_wire[307];							inform_R[282][8] = r_cell_wire[308];							inform_R[410][8] = r_cell_wire[309];							inform_R[283][8] = r_cell_wire[310];							inform_R[411][8] = r_cell_wire[311];							inform_R[284][8] = r_cell_wire[312];							inform_R[412][8] = r_cell_wire[313];							inform_R[285][8] = r_cell_wire[314];							inform_R[413][8] = r_cell_wire[315];							inform_R[286][8] = r_cell_wire[316];							inform_R[414][8] = r_cell_wire[317];							inform_R[287][8] = r_cell_wire[318];							inform_R[415][8] = r_cell_wire[319];							inform_R[288][8] = r_cell_wire[320];							inform_R[416][8] = r_cell_wire[321];							inform_R[289][8] = r_cell_wire[322];							inform_R[417][8] = r_cell_wire[323];							inform_R[290][8] = r_cell_wire[324];							inform_R[418][8] = r_cell_wire[325];							inform_R[291][8] = r_cell_wire[326];							inform_R[419][8] = r_cell_wire[327];							inform_R[292][8] = r_cell_wire[328];							inform_R[420][8] = r_cell_wire[329];							inform_R[293][8] = r_cell_wire[330];							inform_R[421][8] = r_cell_wire[331];							inform_R[294][8] = r_cell_wire[332];							inform_R[422][8] = r_cell_wire[333];							inform_R[295][8] = r_cell_wire[334];							inform_R[423][8] = r_cell_wire[335];							inform_R[296][8] = r_cell_wire[336];							inform_R[424][8] = r_cell_wire[337];							inform_R[297][8] = r_cell_wire[338];							inform_R[425][8] = r_cell_wire[339];							inform_R[298][8] = r_cell_wire[340];							inform_R[426][8] = r_cell_wire[341];							inform_R[299][8] = r_cell_wire[342];							inform_R[427][8] = r_cell_wire[343];							inform_R[300][8] = r_cell_wire[344];							inform_R[428][8] = r_cell_wire[345];							inform_R[301][8] = r_cell_wire[346];							inform_R[429][8] = r_cell_wire[347];							inform_R[302][8] = r_cell_wire[348];							inform_R[430][8] = r_cell_wire[349];							inform_R[303][8] = r_cell_wire[350];							inform_R[431][8] = r_cell_wire[351];							inform_R[304][8] = r_cell_wire[352];							inform_R[432][8] = r_cell_wire[353];							inform_R[305][8] = r_cell_wire[354];							inform_R[433][8] = r_cell_wire[355];							inform_R[306][8] = r_cell_wire[356];							inform_R[434][8] = r_cell_wire[357];							inform_R[307][8] = r_cell_wire[358];							inform_R[435][8] = r_cell_wire[359];							inform_R[308][8] = r_cell_wire[360];							inform_R[436][8] = r_cell_wire[361];							inform_R[309][8] = r_cell_wire[362];							inform_R[437][8] = r_cell_wire[363];							inform_R[310][8] = r_cell_wire[364];							inform_R[438][8] = r_cell_wire[365];							inform_R[311][8] = r_cell_wire[366];							inform_R[439][8] = r_cell_wire[367];							inform_R[312][8] = r_cell_wire[368];							inform_R[440][8] = r_cell_wire[369];							inform_R[313][8] = r_cell_wire[370];							inform_R[441][8] = r_cell_wire[371];							inform_R[314][8] = r_cell_wire[372];							inform_R[442][8] = r_cell_wire[373];							inform_R[315][8] = r_cell_wire[374];							inform_R[443][8] = r_cell_wire[375];							inform_R[316][8] = r_cell_wire[376];							inform_R[444][8] = r_cell_wire[377];							inform_R[317][8] = r_cell_wire[378];							inform_R[445][8] = r_cell_wire[379];							inform_R[318][8] = r_cell_wire[380];							inform_R[446][8] = r_cell_wire[381];							inform_R[319][8] = r_cell_wire[382];							inform_R[447][8] = r_cell_wire[383];							inform_R[320][8] = r_cell_wire[384];							inform_R[448][8] = r_cell_wire[385];							inform_R[321][8] = r_cell_wire[386];							inform_R[449][8] = r_cell_wire[387];							inform_R[322][8] = r_cell_wire[388];							inform_R[450][8] = r_cell_wire[389];							inform_R[323][8] = r_cell_wire[390];							inform_R[451][8] = r_cell_wire[391];							inform_R[324][8] = r_cell_wire[392];							inform_R[452][8] = r_cell_wire[393];							inform_R[325][8] = r_cell_wire[394];							inform_R[453][8] = r_cell_wire[395];							inform_R[326][8] = r_cell_wire[396];							inform_R[454][8] = r_cell_wire[397];							inform_R[327][8] = r_cell_wire[398];							inform_R[455][8] = r_cell_wire[399];							inform_R[328][8] = r_cell_wire[400];							inform_R[456][8] = r_cell_wire[401];							inform_R[329][8] = r_cell_wire[402];							inform_R[457][8] = r_cell_wire[403];							inform_R[330][8] = r_cell_wire[404];							inform_R[458][8] = r_cell_wire[405];							inform_R[331][8] = r_cell_wire[406];							inform_R[459][8] = r_cell_wire[407];							inform_R[332][8] = r_cell_wire[408];							inform_R[460][8] = r_cell_wire[409];							inform_R[333][8] = r_cell_wire[410];							inform_R[461][8] = r_cell_wire[411];							inform_R[334][8] = r_cell_wire[412];							inform_R[462][8] = r_cell_wire[413];							inform_R[335][8] = r_cell_wire[414];							inform_R[463][8] = r_cell_wire[415];							inform_R[336][8] = r_cell_wire[416];							inform_R[464][8] = r_cell_wire[417];							inform_R[337][8] = r_cell_wire[418];							inform_R[465][8] = r_cell_wire[419];							inform_R[338][8] = r_cell_wire[420];							inform_R[466][8] = r_cell_wire[421];							inform_R[339][8] = r_cell_wire[422];							inform_R[467][8] = r_cell_wire[423];							inform_R[340][8] = r_cell_wire[424];							inform_R[468][8] = r_cell_wire[425];							inform_R[341][8] = r_cell_wire[426];							inform_R[469][8] = r_cell_wire[427];							inform_R[342][8] = r_cell_wire[428];							inform_R[470][8] = r_cell_wire[429];							inform_R[343][8] = r_cell_wire[430];							inform_R[471][8] = r_cell_wire[431];							inform_R[344][8] = r_cell_wire[432];							inform_R[472][8] = r_cell_wire[433];							inform_R[345][8] = r_cell_wire[434];							inform_R[473][8] = r_cell_wire[435];							inform_R[346][8] = r_cell_wire[436];							inform_R[474][8] = r_cell_wire[437];							inform_R[347][8] = r_cell_wire[438];							inform_R[475][8] = r_cell_wire[439];							inform_R[348][8] = r_cell_wire[440];							inform_R[476][8] = r_cell_wire[441];							inform_R[349][8] = r_cell_wire[442];							inform_R[477][8] = r_cell_wire[443];							inform_R[350][8] = r_cell_wire[444];							inform_R[478][8] = r_cell_wire[445];							inform_R[351][8] = r_cell_wire[446];							inform_R[479][8] = r_cell_wire[447];							inform_R[352][8] = r_cell_wire[448];							inform_R[480][8] = r_cell_wire[449];							inform_R[353][8] = r_cell_wire[450];							inform_R[481][8] = r_cell_wire[451];							inform_R[354][8] = r_cell_wire[452];							inform_R[482][8] = r_cell_wire[453];							inform_R[355][8] = r_cell_wire[454];							inform_R[483][8] = r_cell_wire[455];							inform_R[356][8] = r_cell_wire[456];							inform_R[484][8] = r_cell_wire[457];							inform_R[357][8] = r_cell_wire[458];							inform_R[485][8] = r_cell_wire[459];							inform_R[358][8] = r_cell_wire[460];							inform_R[486][8] = r_cell_wire[461];							inform_R[359][8] = r_cell_wire[462];							inform_R[487][8] = r_cell_wire[463];							inform_R[360][8] = r_cell_wire[464];							inform_R[488][8] = r_cell_wire[465];							inform_R[361][8] = r_cell_wire[466];							inform_R[489][8] = r_cell_wire[467];							inform_R[362][8] = r_cell_wire[468];							inform_R[490][8] = r_cell_wire[469];							inform_R[363][8] = r_cell_wire[470];							inform_R[491][8] = r_cell_wire[471];							inform_R[364][8] = r_cell_wire[472];							inform_R[492][8] = r_cell_wire[473];							inform_R[365][8] = r_cell_wire[474];							inform_R[493][8] = r_cell_wire[475];							inform_R[366][8] = r_cell_wire[476];							inform_R[494][8] = r_cell_wire[477];							inform_R[367][8] = r_cell_wire[478];							inform_R[495][8] = r_cell_wire[479];							inform_R[368][8] = r_cell_wire[480];							inform_R[496][8] = r_cell_wire[481];							inform_R[369][8] = r_cell_wire[482];							inform_R[497][8] = r_cell_wire[483];							inform_R[370][8] = r_cell_wire[484];							inform_R[498][8] = r_cell_wire[485];							inform_R[371][8] = r_cell_wire[486];							inform_R[499][8] = r_cell_wire[487];							inform_R[372][8] = r_cell_wire[488];							inform_R[500][8] = r_cell_wire[489];							inform_R[373][8] = r_cell_wire[490];							inform_R[501][8] = r_cell_wire[491];							inform_R[374][8] = r_cell_wire[492];							inform_R[502][8] = r_cell_wire[493];							inform_R[375][8] = r_cell_wire[494];							inform_R[503][8] = r_cell_wire[495];							inform_R[376][8] = r_cell_wire[496];							inform_R[504][8] = r_cell_wire[497];							inform_R[377][8] = r_cell_wire[498];							inform_R[505][8] = r_cell_wire[499];							inform_R[378][8] = r_cell_wire[500];							inform_R[506][8] = r_cell_wire[501];							inform_R[379][8] = r_cell_wire[502];							inform_R[507][8] = r_cell_wire[503];							inform_R[380][8] = r_cell_wire[504];							inform_R[508][8] = r_cell_wire[505];							inform_R[381][8] = r_cell_wire[506];							inform_R[509][8] = r_cell_wire[507];							inform_R[382][8] = r_cell_wire[508];							inform_R[510][8] = r_cell_wire[509];							inform_R[383][8] = r_cell_wire[510];							inform_R[511][8] = r_cell_wire[511];							inform_R[512][8] = r_cell_wire[512];							inform_R[640][8] = r_cell_wire[513];							inform_R[513][8] = r_cell_wire[514];							inform_R[641][8] = r_cell_wire[515];							inform_R[514][8] = r_cell_wire[516];							inform_R[642][8] = r_cell_wire[517];							inform_R[515][8] = r_cell_wire[518];							inform_R[643][8] = r_cell_wire[519];							inform_R[516][8] = r_cell_wire[520];							inform_R[644][8] = r_cell_wire[521];							inform_R[517][8] = r_cell_wire[522];							inform_R[645][8] = r_cell_wire[523];							inform_R[518][8] = r_cell_wire[524];							inform_R[646][8] = r_cell_wire[525];							inform_R[519][8] = r_cell_wire[526];							inform_R[647][8] = r_cell_wire[527];							inform_R[520][8] = r_cell_wire[528];							inform_R[648][8] = r_cell_wire[529];							inform_R[521][8] = r_cell_wire[530];							inform_R[649][8] = r_cell_wire[531];							inform_R[522][8] = r_cell_wire[532];							inform_R[650][8] = r_cell_wire[533];							inform_R[523][8] = r_cell_wire[534];							inform_R[651][8] = r_cell_wire[535];							inform_R[524][8] = r_cell_wire[536];							inform_R[652][8] = r_cell_wire[537];							inform_R[525][8] = r_cell_wire[538];							inform_R[653][8] = r_cell_wire[539];							inform_R[526][8] = r_cell_wire[540];							inform_R[654][8] = r_cell_wire[541];							inform_R[527][8] = r_cell_wire[542];							inform_R[655][8] = r_cell_wire[543];							inform_R[528][8] = r_cell_wire[544];							inform_R[656][8] = r_cell_wire[545];							inform_R[529][8] = r_cell_wire[546];							inform_R[657][8] = r_cell_wire[547];							inform_R[530][8] = r_cell_wire[548];							inform_R[658][8] = r_cell_wire[549];							inform_R[531][8] = r_cell_wire[550];							inform_R[659][8] = r_cell_wire[551];							inform_R[532][8] = r_cell_wire[552];							inform_R[660][8] = r_cell_wire[553];							inform_R[533][8] = r_cell_wire[554];							inform_R[661][8] = r_cell_wire[555];							inform_R[534][8] = r_cell_wire[556];							inform_R[662][8] = r_cell_wire[557];							inform_R[535][8] = r_cell_wire[558];							inform_R[663][8] = r_cell_wire[559];							inform_R[536][8] = r_cell_wire[560];							inform_R[664][8] = r_cell_wire[561];							inform_R[537][8] = r_cell_wire[562];							inform_R[665][8] = r_cell_wire[563];							inform_R[538][8] = r_cell_wire[564];							inform_R[666][8] = r_cell_wire[565];							inform_R[539][8] = r_cell_wire[566];							inform_R[667][8] = r_cell_wire[567];							inform_R[540][8] = r_cell_wire[568];							inform_R[668][8] = r_cell_wire[569];							inform_R[541][8] = r_cell_wire[570];							inform_R[669][8] = r_cell_wire[571];							inform_R[542][8] = r_cell_wire[572];							inform_R[670][8] = r_cell_wire[573];							inform_R[543][8] = r_cell_wire[574];							inform_R[671][8] = r_cell_wire[575];							inform_R[544][8] = r_cell_wire[576];							inform_R[672][8] = r_cell_wire[577];							inform_R[545][8] = r_cell_wire[578];							inform_R[673][8] = r_cell_wire[579];							inform_R[546][8] = r_cell_wire[580];							inform_R[674][8] = r_cell_wire[581];							inform_R[547][8] = r_cell_wire[582];							inform_R[675][8] = r_cell_wire[583];							inform_R[548][8] = r_cell_wire[584];							inform_R[676][8] = r_cell_wire[585];							inform_R[549][8] = r_cell_wire[586];							inform_R[677][8] = r_cell_wire[587];							inform_R[550][8] = r_cell_wire[588];							inform_R[678][8] = r_cell_wire[589];							inform_R[551][8] = r_cell_wire[590];							inform_R[679][8] = r_cell_wire[591];							inform_R[552][8] = r_cell_wire[592];							inform_R[680][8] = r_cell_wire[593];							inform_R[553][8] = r_cell_wire[594];							inform_R[681][8] = r_cell_wire[595];							inform_R[554][8] = r_cell_wire[596];							inform_R[682][8] = r_cell_wire[597];							inform_R[555][8] = r_cell_wire[598];							inform_R[683][8] = r_cell_wire[599];							inform_R[556][8] = r_cell_wire[600];							inform_R[684][8] = r_cell_wire[601];							inform_R[557][8] = r_cell_wire[602];							inform_R[685][8] = r_cell_wire[603];							inform_R[558][8] = r_cell_wire[604];							inform_R[686][8] = r_cell_wire[605];							inform_R[559][8] = r_cell_wire[606];							inform_R[687][8] = r_cell_wire[607];							inform_R[560][8] = r_cell_wire[608];							inform_R[688][8] = r_cell_wire[609];							inform_R[561][8] = r_cell_wire[610];							inform_R[689][8] = r_cell_wire[611];							inform_R[562][8] = r_cell_wire[612];							inform_R[690][8] = r_cell_wire[613];							inform_R[563][8] = r_cell_wire[614];							inform_R[691][8] = r_cell_wire[615];							inform_R[564][8] = r_cell_wire[616];							inform_R[692][8] = r_cell_wire[617];							inform_R[565][8] = r_cell_wire[618];							inform_R[693][8] = r_cell_wire[619];							inform_R[566][8] = r_cell_wire[620];							inform_R[694][8] = r_cell_wire[621];							inform_R[567][8] = r_cell_wire[622];							inform_R[695][8] = r_cell_wire[623];							inform_R[568][8] = r_cell_wire[624];							inform_R[696][8] = r_cell_wire[625];							inform_R[569][8] = r_cell_wire[626];							inform_R[697][8] = r_cell_wire[627];							inform_R[570][8] = r_cell_wire[628];							inform_R[698][8] = r_cell_wire[629];							inform_R[571][8] = r_cell_wire[630];							inform_R[699][8] = r_cell_wire[631];							inform_R[572][8] = r_cell_wire[632];							inform_R[700][8] = r_cell_wire[633];							inform_R[573][8] = r_cell_wire[634];							inform_R[701][8] = r_cell_wire[635];							inform_R[574][8] = r_cell_wire[636];							inform_R[702][8] = r_cell_wire[637];							inform_R[575][8] = r_cell_wire[638];							inform_R[703][8] = r_cell_wire[639];							inform_R[576][8] = r_cell_wire[640];							inform_R[704][8] = r_cell_wire[641];							inform_R[577][8] = r_cell_wire[642];							inform_R[705][8] = r_cell_wire[643];							inform_R[578][8] = r_cell_wire[644];							inform_R[706][8] = r_cell_wire[645];							inform_R[579][8] = r_cell_wire[646];							inform_R[707][8] = r_cell_wire[647];							inform_R[580][8] = r_cell_wire[648];							inform_R[708][8] = r_cell_wire[649];							inform_R[581][8] = r_cell_wire[650];							inform_R[709][8] = r_cell_wire[651];							inform_R[582][8] = r_cell_wire[652];							inform_R[710][8] = r_cell_wire[653];							inform_R[583][8] = r_cell_wire[654];							inform_R[711][8] = r_cell_wire[655];							inform_R[584][8] = r_cell_wire[656];							inform_R[712][8] = r_cell_wire[657];							inform_R[585][8] = r_cell_wire[658];							inform_R[713][8] = r_cell_wire[659];							inform_R[586][8] = r_cell_wire[660];							inform_R[714][8] = r_cell_wire[661];							inform_R[587][8] = r_cell_wire[662];							inform_R[715][8] = r_cell_wire[663];							inform_R[588][8] = r_cell_wire[664];							inform_R[716][8] = r_cell_wire[665];							inform_R[589][8] = r_cell_wire[666];							inform_R[717][8] = r_cell_wire[667];							inform_R[590][8] = r_cell_wire[668];							inform_R[718][8] = r_cell_wire[669];							inform_R[591][8] = r_cell_wire[670];							inform_R[719][8] = r_cell_wire[671];							inform_R[592][8] = r_cell_wire[672];							inform_R[720][8] = r_cell_wire[673];							inform_R[593][8] = r_cell_wire[674];							inform_R[721][8] = r_cell_wire[675];							inform_R[594][8] = r_cell_wire[676];							inform_R[722][8] = r_cell_wire[677];							inform_R[595][8] = r_cell_wire[678];							inform_R[723][8] = r_cell_wire[679];							inform_R[596][8] = r_cell_wire[680];							inform_R[724][8] = r_cell_wire[681];							inform_R[597][8] = r_cell_wire[682];							inform_R[725][8] = r_cell_wire[683];							inform_R[598][8] = r_cell_wire[684];							inform_R[726][8] = r_cell_wire[685];							inform_R[599][8] = r_cell_wire[686];							inform_R[727][8] = r_cell_wire[687];							inform_R[600][8] = r_cell_wire[688];							inform_R[728][8] = r_cell_wire[689];							inform_R[601][8] = r_cell_wire[690];							inform_R[729][8] = r_cell_wire[691];							inform_R[602][8] = r_cell_wire[692];							inform_R[730][8] = r_cell_wire[693];							inform_R[603][8] = r_cell_wire[694];							inform_R[731][8] = r_cell_wire[695];							inform_R[604][8] = r_cell_wire[696];							inform_R[732][8] = r_cell_wire[697];							inform_R[605][8] = r_cell_wire[698];							inform_R[733][8] = r_cell_wire[699];							inform_R[606][8] = r_cell_wire[700];							inform_R[734][8] = r_cell_wire[701];							inform_R[607][8] = r_cell_wire[702];							inform_R[735][8] = r_cell_wire[703];							inform_R[608][8] = r_cell_wire[704];							inform_R[736][8] = r_cell_wire[705];							inform_R[609][8] = r_cell_wire[706];							inform_R[737][8] = r_cell_wire[707];							inform_R[610][8] = r_cell_wire[708];							inform_R[738][8] = r_cell_wire[709];							inform_R[611][8] = r_cell_wire[710];							inform_R[739][8] = r_cell_wire[711];							inform_R[612][8] = r_cell_wire[712];							inform_R[740][8] = r_cell_wire[713];							inform_R[613][8] = r_cell_wire[714];							inform_R[741][8] = r_cell_wire[715];							inform_R[614][8] = r_cell_wire[716];							inform_R[742][8] = r_cell_wire[717];							inform_R[615][8] = r_cell_wire[718];							inform_R[743][8] = r_cell_wire[719];							inform_R[616][8] = r_cell_wire[720];							inform_R[744][8] = r_cell_wire[721];							inform_R[617][8] = r_cell_wire[722];							inform_R[745][8] = r_cell_wire[723];							inform_R[618][8] = r_cell_wire[724];							inform_R[746][8] = r_cell_wire[725];							inform_R[619][8] = r_cell_wire[726];							inform_R[747][8] = r_cell_wire[727];							inform_R[620][8] = r_cell_wire[728];							inform_R[748][8] = r_cell_wire[729];							inform_R[621][8] = r_cell_wire[730];							inform_R[749][8] = r_cell_wire[731];							inform_R[622][8] = r_cell_wire[732];							inform_R[750][8] = r_cell_wire[733];							inform_R[623][8] = r_cell_wire[734];							inform_R[751][8] = r_cell_wire[735];							inform_R[624][8] = r_cell_wire[736];							inform_R[752][8] = r_cell_wire[737];							inform_R[625][8] = r_cell_wire[738];							inform_R[753][8] = r_cell_wire[739];							inform_R[626][8] = r_cell_wire[740];							inform_R[754][8] = r_cell_wire[741];							inform_R[627][8] = r_cell_wire[742];							inform_R[755][8] = r_cell_wire[743];							inform_R[628][8] = r_cell_wire[744];							inform_R[756][8] = r_cell_wire[745];							inform_R[629][8] = r_cell_wire[746];							inform_R[757][8] = r_cell_wire[747];							inform_R[630][8] = r_cell_wire[748];							inform_R[758][8] = r_cell_wire[749];							inform_R[631][8] = r_cell_wire[750];							inform_R[759][8] = r_cell_wire[751];							inform_R[632][8] = r_cell_wire[752];							inform_R[760][8] = r_cell_wire[753];							inform_R[633][8] = r_cell_wire[754];							inform_R[761][8] = r_cell_wire[755];							inform_R[634][8] = r_cell_wire[756];							inform_R[762][8] = r_cell_wire[757];							inform_R[635][8] = r_cell_wire[758];							inform_R[763][8] = r_cell_wire[759];							inform_R[636][8] = r_cell_wire[760];							inform_R[764][8] = r_cell_wire[761];							inform_R[637][8] = r_cell_wire[762];							inform_R[765][8] = r_cell_wire[763];							inform_R[638][8] = r_cell_wire[764];							inform_R[766][8] = r_cell_wire[765];							inform_R[639][8] = r_cell_wire[766];							inform_R[767][8] = r_cell_wire[767];							inform_R[768][8] = r_cell_wire[768];							inform_R[896][8] = r_cell_wire[769];							inform_R[769][8] = r_cell_wire[770];							inform_R[897][8] = r_cell_wire[771];							inform_R[770][8] = r_cell_wire[772];							inform_R[898][8] = r_cell_wire[773];							inform_R[771][8] = r_cell_wire[774];							inform_R[899][8] = r_cell_wire[775];							inform_R[772][8] = r_cell_wire[776];							inform_R[900][8] = r_cell_wire[777];							inform_R[773][8] = r_cell_wire[778];							inform_R[901][8] = r_cell_wire[779];							inform_R[774][8] = r_cell_wire[780];							inform_R[902][8] = r_cell_wire[781];							inform_R[775][8] = r_cell_wire[782];							inform_R[903][8] = r_cell_wire[783];							inform_R[776][8] = r_cell_wire[784];							inform_R[904][8] = r_cell_wire[785];							inform_R[777][8] = r_cell_wire[786];							inform_R[905][8] = r_cell_wire[787];							inform_R[778][8] = r_cell_wire[788];							inform_R[906][8] = r_cell_wire[789];							inform_R[779][8] = r_cell_wire[790];							inform_R[907][8] = r_cell_wire[791];							inform_R[780][8] = r_cell_wire[792];							inform_R[908][8] = r_cell_wire[793];							inform_R[781][8] = r_cell_wire[794];							inform_R[909][8] = r_cell_wire[795];							inform_R[782][8] = r_cell_wire[796];							inform_R[910][8] = r_cell_wire[797];							inform_R[783][8] = r_cell_wire[798];							inform_R[911][8] = r_cell_wire[799];							inform_R[784][8] = r_cell_wire[800];							inform_R[912][8] = r_cell_wire[801];							inform_R[785][8] = r_cell_wire[802];							inform_R[913][8] = r_cell_wire[803];							inform_R[786][8] = r_cell_wire[804];							inform_R[914][8] = r_cell_wire[805];							inform_R[787][8] = r_cell_wire[806];							inform_R[915][8] = r_cell_wire[807];							inform_R[788][8] = r_cell_wire[808];							inform_R[916][8] = r_cell_wire[809];							inform_R[789][8] = r_cell_wire[810];							inform_R[917][8] = r_cell_wire[811];							inform_R[790][8] = r_cell_wire[812];							inform_R[918][8] = r_cell_wire[813];							inform_R[791][8] = r_cell_wire[814];							inform_R[919][8] = r_cell_wire[815];							inform_R[792][8] = r_cell_wire[816];							inform_R[920][8] = r_cell_wire[817];							inform_R[793][8] = r_cell_wire[818];							inform_R[921][8] = r_cell_wire[819];							inform_R[794][8] = r_cell_wire[820];							inform_R[922][8] = r_cell_wire[821];							inform_R[795][8] = r_cell_wire[822];							inform_R[923][8] = r_cell_wire[823];							inform_R[796][8] = r_cell_wire[824];							inform_R[924][8] = r_cell_wire[825];							inform_R[797][8] = r_cell_wire[826];							inform_R[925][8] = r_cell_wire[827];							inform_R[798][8] = r_cell_wire[828];							inform_R[926][8] = r_cell_wire[829];							inform_R[799][8] = r_cell_wire[830];							inform_R[927][8] = r_cell_wire[831];							inform_R[800][8] = r_cell_wire[832];							inform_R[928][8] = r_cell_wire[833];							inform_R[801][8] = r_cell_wire[834];							inform_R[929][8] = r_cell_wire[835];							inform_R[802][8] = r_cell_wire[836];							inform_R[930][8] = r_cell_wire[837];							inform_R[803][8] = r_cell_wire[838];							inform_R[931][8] = r_cell_wire[839];							inform_R[804][8] = r_cell_wire[840];							inform_R[932][8] = r_cell_wire[841];							inform_R[805][8] = r_cell_wire[842];							inform_R[933][8] = r_cell_wire[843];							inform_R[806][8] = r_cell_wire[844];							inform_R[934][8] = r_cell_wire[845];							inform_R[807][8] = r_cell_wire[846];							inform_R[935][8] = r_cell_wire[847];							inform_R[808][8] = r_cell_wire[848];							inform_R[936][8] = r_cell_wire[849];							inform_R[809][8] = r_cell_wire[850];							inform_R[937][8] = r_cell_wire[851];							inform_R[810][8] = r_cell_wire[852];							inform_R[938][8] = r_cell_wire[853];							inform_R[811][8] = r_cell_wire[854];							inform_R[939][8] = r_cell_wire[855];							inform_R[812][8] = r_cell_wire[856];							inform_R[940][8] = r_cell_wire[857];							inform_R[813][8] = r_cell_wire[858];							inform_R[941][8] = r_cell_wire[859];							inform_R[814][8] = r_cell_wire[860];							inform_R[942][8] = r_cell_wire[861];							inform_R[815][8] = r_cell_wire[862];							inform_R[943][8] = r_cell_wire[863];							inform_R[816][8] = r_cell_wire[864];							inform_R[944][8] = r_cell_wire[865];							inform_R[817][8] = r_cell_wire[866];							inform_R[945][8] = r_cell_wire[867];							inform_R[818][8] = r_cell_wire[868];							inform_R[946][8] = r_cell_wire[869];							inform_R[819][8] = r_cell_wire[870];							inform_R[947][8] = r_cell_wire[871];							inform_R[820][8] = r_cell_wire[872];							inform_R[948][8] = r_cell_wire[873];							inform_R[821][8] = r_cell_wire[874];							inform_R[949][8] = r_cell_wire[875];							inform_R[822][8] = r_cell_wire[876];							inform_R[950][8] = r_cell_wire[877];							inform_R[823][8] = r_cell_wire[878];							inform_R[951][8] = r_cell_wire[879];							inform_R[824][8] = r_cell_wire[880];							inform_R[952][8] = r_cell_wire[881];							inform_R[825][8] = r_cell_wire[882];							inform_R[953][8] = r_cell_wire[883];							inform_R[826][8] = r_cell_wire[884];							inform_R[954][8] = r_cell_wire[885];							inform_R[827][8] = r_cell_wire[886];							inform_R[955][8] = r_cell_wire[887];							inform_R[828][8] = r_cell_wire[888];							inform_R[956][8] = r_cell_wire[889];							inform_R[829][8] = r_cell_wire[890];							inform_R[957][8] = r_cell_wire[891];							inform_R[830][8] = r_cell_wire[892];							inform_R[958][8] = r_cell_wire[893];							inform_R[831][8] = r_cell_wire[894];							inform_R[959][8] = r_cell_wire[895];							inform_R[832][8] = r_cell_wire[896];							inform_R[960][8] = r_cell_wire[897];							inform_R[833][8] = r_cell_wire[898];							inform_R[961][8] = r_cell_wire[899];							inform_R[834][8] = r_cell_wire[900];							inform_R[962][8] = r_cell_wire[901];							inform_R[835][8] = r_cell_wire[902];							inform_R[963][8] = r_cell_wire[903];							inform_R[836][8] = r_cell_wire[904];							inform_R[964][8] = r_cell_wire[905];							inform_R[837][8] = r_cell_wire[906];							inform_R[965][8] = r_cell_wire[907];							inform_R[838][8] = r_cell_wire[908];							inform_R[966][8] = r_cell_wire[909];							inform_R[839][8] = r_cell_wire[910];							inform_R[967][8] = r_cell_wire[911];							inform_R[840][8] = r_cell_wire[912];							inform_R[968][8] = r_cell_wire[913];							inform_R[841][8] = r_cell_wire[914];							inform_R[969][8] = r_cell_wire[915];							inform_R[842][8] = r_cell_wire[916];							inform_R[970][8] = r_cell_wire[917];							inform_R[843][8] = r_cell_wire[918];							inform_R[971][8] = r_cell_wire[919];							inform_R[844][8] = r_cell_wire[920];							inform_R[972][8] = r_cell_wire[921];							inform_R[845][8] = r_cell_wire[922];							inform_R[973][8] = r_cell_wire[923];							inform_R[846][8] = r_cell_wire[924];							inform_R[974][8] = r_cell_wire[925];							inform_R[847][8] = r_cell_wire[926];							inform_R[975][8] = r_cell_wire[927];							inform_R[848][8] = r_cell_wire[928];							inform_R[976][8] = r_cell_wire[929];							inform_R[849][8] = r_cell_wire[930];							inform_R[977][8] = r_cell_wire[931];							inform_R[850][8] = r_cell_wire[932];							inform_R[978][8] = r_cell_wire[933];							inform_R[851][8] = r_cell_wire[934];							inform_R[979][8] = r_cell_wire[935];							inform_R[852][8] = r_cell_wire[936];							inform_R[980][8] = r_cell_wire[937];							inform_R[853][8] = r_cell_wire[938];							inform_R[981][8] = r_cell_wire[939];							inform_R[854][8] = r_cell_wire[940];							inform_R[982][8] = r_cell_wire[941];							inform_R[855][8] = r_cell_wire[942];							inform_R[983][8] = r_cell_wire[943];							inform_R[856][8] = r_cell_wire[944];							inform_R[984][8] = r_cell_wire[945];							inform_R[857][8] = r_cell_wire[946];							inform_R[985][8] = r_cell_wire[947];							inform_R[858][8] = r_cell_wire[948];							inform_R[986][8] = r_cell_wire[949];							inform_R[859][8] = r_cell_wire[950];							inform_R[987][8] = r_cell_wire[951];							inform_R[860][8] = r_cell_wire[952];							inform_R[988][8] = r_cell_wire[953];							inform_R[861][8] = r_cell_wire[954];							inform_R[989][8] = r_cell_wire[955];							inform_R[862][8] = r_cell_wire[956];							inform_R[990][8] = r_cell_wire[957];							inform_R[863][8] = r_cell_wire[958];							inform_R[991][8] = r_cell_wire[959];							inform_R[864][8] = r_cell_wire[960];							inform_R[992][8] = r_cell_wire[961];							inform_R[865][8] = r_cell_wire[962];							inform_R[993][8] = r_cell_wire[963];							inform_R[866][8] = r_cell_wire[964];							inform_R[994][8] = r_cell_wire[965];							inform_R[867][8] = r_cell_wire[966];							inform_R[995][8] = r_cell_wire[967];							inform_R[868][8] = r_cell_wire[968];							inform_R[996][8] = r_cell_wire[969];							inform_R[869][8] = r_cell_wire[970];							inform_R[997][8] = r_cell_wire[971];							inform_R[870][8] = r_cell_wire[972];							inform_R[998][8] = r_cell_wire[973];							inform_R[871][8] = r_cell_wire[974];							inform_R[999][8] = r_cell_wire[975];							inform_R[872][8] = r_cell_wire[976];							inform_R[1000][8] = r_cell_wire[977];							inform_R[873][8] = r_cell_wire[978];							inform_R[1001][8] = r_cell_wire[979];							inform_R[874][8] = r_cell_wire[980];							inform_R[1002][8] = r_cell_wire[981];							inform_R[875][8] = r_cell_wire[982];							inform_R[1003][8] = r_cell_wire[983];							inform_R[876][8] = r_cell_wire[984];							inform_R[1004][8] = r_cell_wire[985];							inform_R[877][8] = r_cell_wire[986];							inform_R[1005][8] = r_cell_wire[987];							inform_R[878][8] = r_cell_wire[988];							inform_R[1006][8] = r_cell_wire[989];							inform_R[879][8] = r_cell_wire[990];							inform_R[1007][8] = r_cell_wire[991];							inform_R[880][8] = r_cell_wire[992];							inform_R[1008][8] = r_cell_wire[993];							inform_R[881][8] = r_cell_wire[994];							inform_R[1009][8] = r_cell_wire[995];							inform_R[882][8] = r_cell_wire[996];							inform_R[1010][8] = r_cell_wire[997];							inform_R[883][8] = r_cell_wire[998];							inform_R[1011][8] = r_cell_wire[999];							inform_R[884][8] = r_cell_wire[1000];							inform_R[1012][8] = r_cell_wire[1001];							inform_R[885][8] = r_cell_wire[1002];							inform_R[1013][8] = r_cell_wire[1003];							inform_R[886][8] = r_cell_wire[1004];							inform_R[1014][8] = r_cell_wire[1005];							inform_R[887][8] = r_cell_wire[1006];							inform_R[1015][8] = r_cell_wire[1007];							inform_R[888][8] = r_cell_wire[1008];							inform_R[1016][8] = r_cell_wire[1009];							inform_R[889][8] = r_cell_wire[1010];							inform_R[1017][8] = r_cell_wire[1011];							inform_R[890][8] = r_cell_wire[1012];							inform_R[1018][8] = r_cell_wire[1013];							inform_R[891][8] = r_cell_wire[1014];							inform_R[1019][8] = r_cell_wire[1015];							inform_R[892][8] = r_cell_wire[1016];							inform_R[1020][8] = r_cell_wire[1017];							inform_R[893][8] = r_cell_wire[1018];							inform_R[1021][8] = r_cell_wire[1019];							inform_R[894][8] = r_cell_wire[1020];							inform_R[1022][8] = r_cell_wire[1021];							inform_R[895][8] = r_cell_wire[1022];							inform_R[1023][8] = r_cell_wire[1023];							inform_L[0][7] = l_cell_wire[0];							inform_L[128][7] = l_cell_wire[1];							inform_L[1][7] = l_cell_wire[2];							inform_L[129][7] = l_cell_wire[3];							inform_L[2][7] = l_cell_wire[4];							inform_L[130][7] = l_cell_wire[5];							inform_L[3][7] = l_cell_wire[6];							inform_L[131][7] = l_cell_wire[7];							inform_L[4][7] = l_cell_wire[8];							inform_L[132][7] = l_cell_wire[9];							inform_L[5][7] = l_cell_wire[10];							inform_L[133][7] = l_cell_wire[11];							inform_L[6][7] = l_cell_wire[12];							inform_L[134][7] = l_cell_wire[13];							inform_L[7][7] = l_cell_wire[14];							inform_L[135][7] = l_cell_wire[15];							inform_L[8][7] = l_cell_wire[16];							inform_L[136][7] = l_cell_wire[17];							inform_L[9][7] = l_cell_wire[18];							inform_L[137][7] = l_cell_wire[19];							inform_L[10][7] = l_cell_wire[20];							inform_L[138][7] = l_cell_wire[21];							inform_L[11][7] = l_cell_wire[22];							inform_L[139][7] = l_cell_wire[23];							inform_L[12][7] = l_cell_wire[24];							inform_L[140][7] = l_cell_wire[25];							inform_L[13][7] = l_cell_wire[26];							inform_L[141][7] = l_cell_wire[27];							inform_L[14][7] = l_cell_wire[28];							inform_L[142][7] = l_cell_wire[29];							inform_L[15][7] = l_cell_wire[30];							inform_L[143][7] = l_cell_wire[31];							inform_L[16][7] = l_cell_wire[32];							inform_L[144][7] = l_cell_wire[33];							inform_L[17][7] = l_cell_wire[34];							inform_L[145][7] = l_cell_wire[35];							inform_L[18][7] = l_cell_wire[36];							inform_L[146][7] = l_cell_wire[37];							inform_L[19][7] = l_cell_wire[38];							inform_L[147][7] = l_cell_wire[39];							inform_L[20][7] = l_cell_wire[40];							inform_L[148][7] = l_cell_wire[41];							inform_L[21][7] = l_cell_wire[42];							inform_L[149][7] = l_cell_wire[43];							inform_L[22][7] = l_cell_wire[44];							inform_L[150][7] = l_cell_wire[45];							inform_L[23][7] = l_cell_wire[46];							inform_L[151][7] = l_cell_wire[47];							inform_L[24][7] = l_cell_wire[48];							inform_L[152][7] = l_cell_wire[49];							inform_L[25][7] = l_cell_wire[50];							inform_L[153][7] = l_cell_wire[51];							inform_L[26][7] = l_cell_wire[52];							inform_L[154][7] = l_cell_wire[53];							inform_L[27][7] = l_cell_wire[54];							inform_L[155][7] = l_cell_wire[55];							inform_L[28][7] = l_cell_wire[56];							inform_L[156][7] = l_cell_wire[57];							inform_L[29][7] = l_cell_wire[58];							inform_L[157][7] = l_cell_wire[59];							inform_L[30][7] = l_cell_wire[60];							inform_L[158][7] = l_cell_wire[61];							inform_L[31][7] = l_cell_wire[62];							inform_L[159][7] = l_cell_wire[63];							inform_L[32][7] = l_cell_wire[64];							inform_L[160][7] = l_cell_wire[65];							inform_L[33][7] = l_cell_wire[66];							inform_L[161][7] = l_cell_wire[67];							inform_L[34][7] = l_cell_wire[68];							inform_L[162][7] = l_cell_wire[69];							inform_L[35][7] = l_cell_wire[70];							inform_L[163][7] = l_cell_wire[71];							inform_L[36][7] = l_cell_wire[72];							inform_L[164][7] = l_cell_wire[73];							inform_L[37][7] = l_cell_wire[74];							inform_L[165][7] = l_cell_wire[75];							inform_L[38][7] = l_cell_wire[76];							inform_L[166][7] = l_cell_wire[77];							inform_L[39][7] = l_cell_wire[78];							inform_L[167][7] = l_cell_wire[79];							inform_L[40][7] = l_cell_wire[80];							inform_L[168][7] = l_cell_wire[81];							inform_L[41][7] = l_cell_wire[82];							inform_L[169][7] = l_cell_wire[83];							inform_L[42][7] = l_cell_wire[84];							inform_L[170][7] = l_cell_wire[85];							inform_L[43][7] = l_cell_wire[86];							inform_L[171][7] = l_cell_wire[87];							inform_L[44][7] = l_cell_wire[88];							inform_L[172][7] = l_cell_wire[89];							inform_L[45][7] = l_cell_wire[90];							inform_L[173][7] = l_cell_wire[91];							inform_L[46][7] = l_cell_wire[92];							inform_L[174][7] = l_cell_wire[93];							inform_L[47][7] = l_cell_wire[94];							inform_L[175][7] = l_cell_wire[95];							inform_L[48][7] = l_cell_wire[96];							inform_L[176][7] = l_cell_wire[97];							inform_L[49][7] = l_cell_wire[98];							inform_L[177][7] = l_cell_wire[99];							inform_L[50][7] = l_cell_wire[100];							inform_L[178][7] = l_cell_wire[101];							inform_L[51][7] = l_cell_wire[102];							inform_L[179][7] = l_cell_wire[103];							inform_L[52][7] = l_cell_wire[104];							inform_L[180][7] = l_cell_wire[105];							inform_L[53][7] = l_cell_wire[106];							inform_L[181][7] = l_cell_wire[107];							inform_L[54][7] = l_cell_wire[108];							inform_L[182][7] = l_cell_wire[109];							inform_L[55][7] = l_cell_wire[110];							inform_L[183][7] = l_cell_wire[111];							inform_L[56][7] = l_cell_wire[112];							inform_L[184][7] = l_cell_wire[113];							inform_L[57][7] = l_cell_wire[114];							inform_L[185][7] = l_cell_wire[115];							inform_L[58][7] = l_cell_wire[116];							inform_L[186][7] = l_cell_wire[117];							inform_L[59][7] = l_cell_wire[118];							inform_L[187][7] = l_cell_wire[119];							inform_L[60][7] = l_cell_wire[120];							inform_L[188][7] = l_cell_wire[121];							inform_L[61][7] = l_cell_wire[122];							inform_L[189][7] = l_cell_wire[123];							inform_L[62][7] = l_cell_wire[124];							inform_L[190][7] = l_cell_wire[125];							inform_L[63][7] = l_cell_wire[126];							inform_L[191][7] = l_cell_wire[127];							inform_L[64][7] = l_cell_wire[128];							inform_L[192][7] = l_cell_wire[129];							inform_L[65][7] = l_cell_wire[130];							inform_L[193][7] = l_cell_wire[131];							inform_L[66][7] = l_cell_wire[132];							inform_L[194][7] = l_cell_wire[133];							inform_L[67][7] = l_cell_wire[134];							inform_L[195][7] = l_cell_wire[135];							inform_L[68][7] = l_cell_wire[136];							inform_L[196][7] = l_cell_wire[137];							inform_L[69][7] = l_cell_wire[138];							inform_L[197][7] = l_cell_wire[139];							inform_L[70][7] = l_cell_wire[140];							inform_L[198][7] = l_cell_wire[141];							inform_L[71][7] = l_cell_wire[142];							inform_L[199][7] = l_cell_wire[143];							inform_L[72][7] = l_cell_wire[144];							inform_L[200][7] = l_cell_wire[145];							inform_L[73][7] = l_cell_wire[146];							inform_L[201][7] = l_cell_wire[147];							inform_L[74][7] = l_cell_wire[148];							inform_L[202][7] = l_cell_wire[149];							inform_L[75][7] = l_cell_wire[150];							inform_L[203][7] = l_cell_wire[151];							inform_L[76][7] = l_cell_wire[152];							inform_L[204][7] = l_cell_wire[153];							inform_L[77][7] = l_cell_wire[154];							inform_L[205][7] = l_cell_wire[155];							inform_L[78][7] = l_cell_wire[156];							inform_L[206][7] = l_cell_wire[157];							inform_L[79][7] = l_cell_wire[158];							inform_L[207][7] = l_cell_wire[159];							inform_L[80][7] = l_cell_wire[160];							inform_L[208][7] = l_cell_wire[161];							inform_L[81][7] = l_cell_wire[162];							inform_L[209][7] = l_cell_wire[163];							inform_L[82][7] = l_cell_wire[164];							inform_L[210][7] = l_cell_wire[165];							inform_L[83][7] = l_cell_wire[166];							inform_L[211][7] = l_cell_wire[167];							inform_L[84][7] = l_cell_wire[168];							inform_L[212][7] = l_cell_wire[169];							inform_L[85][7] = l_cell_wire[170];							inform_L[213][7] = l_cell_wire[171];							inform_L[86][7] = l_cell_wire[172];							inform_L[214][7] = l_cell_wire[173];							inform_L[87][7] = l_cell_wire[174];							inform_L[215][7] = l_cell_wire[175];							inform_L[88][7] = l_cell_wire[176];							inform_L[216][7] = l_cell_wire[177];							inform_L[89][7] = l_cell_wire[178];							inform_L[217][7] = l_cell_wire[179];							inform_L[90][7] = l_cell_wire[180];							inform_L[218][7] = l_cell_wire[181];							inform_L[91][7] = l_cell_wire[182];							inform_L[219][7] = l_cell_wire[183];							inform_L[92][7] = l_cell_wire[184];							inform_L[220][7] = l_cell_wire[185];							inform_L[93][7] = l_cell_wire[186];							inform_L[221][7] = l_cell_wire[187];							inform_L[94][7] = l_cell_wire[188];							inform_L[222][7] = l_cell_wire[189];							inform_L[95][7] = l_cell_wire[190];							inform_L[223][7] = l_cell_wire[191];							inform_L[96][7] = l_cell_wire[192];							inform_L[224][7] = l_cell_wire[193];							inform_L[97][7] = l_cell_wire[194];							inform_L[225][7] = l_cell_wire[195];							inform_L[98][7] = l_cell_wire[196];							inform_L[226][7] = l_cell_wire[197];							inform_L[99][7] = l_cell_wire[198];							inform_L[227][7] = l_cell_wire[199];							inform_L[100][7] = l_cell_wire[200];							inform_L[228][7] = l_cell_wire[201];							inform_L[101][7] = l_cell_wire[202];							inform_L[229][7] = l_cell_wire[203];							inform_L[102][7] = l_cell_wire[204];							inform_L[230][7] = l_cell_wire[205];							inform_L[103][7] = l_cell_wire[206];							inform_L[231][7] = l_cell_wire[207];							inform_L[104][7] = l_cell_wire[208];							inform_L[232][7] = l_cell_wire[209];							inform_L[105][7] = l_cell_wire[210];							inform_L[233][7] = l_cell_wire[211];							inform_L[106][7] = l_cell_wire[212];							inform_L[234][7] = l_cell_wire[213];							inform_L[107][7] = l_cell_wire[214];							inform_L[235][7] = l_cell_wire[215];							inform_L[108][7] = l_cell_wire[216];							inform_L[236][7] = l_cell_wire[217];							inform_L[109][7] = l_cell_wire[218];							inform_L[237][7] = l_cell_wire[219];							inform_L[110][7] = l_cell_wire[220];							inform_L[238][7] = l_cell_wire[221];							inform_L[111][7] = l_cell_wire[222];							inform_L[239][7] = l_cell_wire[223];							inform_L[112][7] = l_cell_wire[224];							inform_L[240][7] = l_cell_wire[225];							inform_L[113][7] = l_cell_wire[226];							inform_L[241][7] = l_cell_wire[227];							inform_L[114][7] = l_cell_wire[228];							inform_L[242][7] = l_cell_wire[229];							inform_L[115][7] = l_cell_wire[230];							inform_L[243][7] = l_cell_wire[231];							inform_L[116][7] = l_cell_wire[232];							inform_L[244][7] = l_cell_wire[233];							inform_L[117][7] = l_cell_wire[234];							inform_L[245][7] = l_cell_wire[235];							inform_L[118][7] = l_cell_wire[236];							inform_L[246][7] = l_cell_wire[237];							inform_L[119][7] = l_cell_wire[238];							inform_L[247][7] = l_cell_wire[239];							inform_L[120][7] = l_cell_wire[240];							inform_L[248][7] = l_cell_wire[241];							inform_L[121][7] = l_cell_wire[242];							inform_L[249][7] = l_cell_wire[243];							inform_L[122][7] = l_cell_wire[244];							inform_L[250][7] = l_cell_wire[245];							inform_L[123][7] = l_cell_wire[246];							inform_L[251][7] = l_cell_wire[247];							inform_L[124][7] = l_cell_wire[248];							inform_L[252][7] = l_cell_wire[249];							inform_L[125][7] = l_cell_wire[250];							inform_L[253][7] = l_cell_wire[251];							inform_L[126][7] = l_cell_wire[252];							inform_L[254][7] = l_cell_wire[253];							inform_L[127][7] = l_cell_wire[254];							inform_L[255][7] = l_cell_wire[255];							inform_L[256][7] = l_cell_wire[256];							inform_L[384][7] = l_cell_wire[257];							inform_L[257][7] = l_cell_wire[258];							inform_L[385][7] = l_cell_wire[259];							inform_L[258][7] = l_cell_wire[260];							inform_L[386][7] = l_cell_wire[261];							inform_L[259][7] = l_cell_wire[262];							inform_L[387][7] = l_cell_wire[263];							inform_L[260][7] = l_cell_wire[264];							inform_L[388][7] = l_cell_wire[265];							inform_L[261][7] = l_cell_wire[266];							inform_L[389][7] = l_cell_wire[267];							inform_L[262][7] = l_cell_wire[268];							inform_L[390][7] = l_cell_wire[269];							inform_L[263][7] = l_cell_wire[270];							inform_L[391][7] = l_cell_wire[271];							inform_L[264][7] = l_cell_wire[272];							inform_L[392][7] = l_cell_wire[273];							inform_L[265][7] = l_cell_wire[274];							inform_L[393][7] = l_cell_wire[275];							inform_L[266][7] = l_cell_wire[276];							inform_L[394][7] = l_cell_wire[277];							inform_L[267][7] = l_cell_wire[278];							inform_L[395][7] = l_cell_wire[279];							inform_L[268][7] = l_cell_wire[280];							inform_L[396][7] = l_cell_wire[281];							inform_L[269][7] = l_cell_wire[282];							inform_L[397][7] = l_cell_wire[283];							inform_L[270][7] = l_cell_wire[284];							inform_L[398][7] = l_cell_wire[285];							inform_L[271][7] = l_cell_wire[286];							inform_L[399][7] = l_cell_wire[287];							inform_L[272][7] = l_cell_wire[288];							inform_L[400][7] = l_cell_wire[289];							inform_L[273][7] = l_cell_wire[290];							inform_L[401][7] = l_cell_wire[291];							inform_L[274][7] = l_cell_wire[292];							inform_L[402][7] = l_cell_wire[293];							inform_L[275][7] = l_cell_wire[294];							inform_L[403][7] = l_cell_wire[295];							inform_L[276][7] = l_cell_wire[296];							inform_L[404][7] = l_cell_wire[297];							inform_L[277][7] = l_cell_wire[298];							inform_L[405][7] = l_cell_wire[299];							inform_L[278][7] = l_cell_wire[300];							inform_L[406][7] = l_cell_wire[301];							inform_L[279][7] = l_cell_wire[302];							inform_L[407][7] = l_cell_wire[303];							inform_L[280][7] = l_cell_wire[304];							inform_L[408][7] = l_cell_wire[305];							inform_L[281][7] = l_cell_wire[306];							inform_L[409][7] = l_cell_wire[307];							inform_L[282][7] = l_cell_wire[308];							inform_L[410][7] = l_cell_wire[309];							inform_L[283][7] = l_cell_wire[310];							inform_L[411][7] = l_cell_wire[311];							inform_L[284][7] = l_cell_wire[312];							inform_L[412][7] = l_cell_wire[313];							inform_L[285][7] = l_cell_wire[314];							inform_L[413][7] = l_cell_wire[315];							inform_L[286][7] = l_cell_wire[316];							inform_L[414][7] = l_cell_wire[317];							inform_L[287][7] = l_cell_wire[318];							inform_L[415][7] = l_cell_wire[319];							inform_L[288][7] = l_cell_wire[320];							inform_L[416][7] = l_cell_wire[321];							inform_L[289][7] = l_cell_wire[322];							inform_L[417][7] = l_cell_wire[323];							inform_L[290][7] = l_cell_wire[324];							inform_L[418][7] = l_cell_wire[325];							inform_L[291][7] = l_cell_wire[326];							inform_L[419][7] = l_cell_wire[327];							inform_L[292][7] = l_cell_wire[328];							inform_L[420][7] = l_cell_wire[329];							inform_L[293][7] = l_cell_wire[330];							inform_L[421][7] = l_cell_wire[331];							inform_L[294][7] = l_cell_wire[332];							inform_L[422][7] = l_cell_wire[333];							inform_L[295][7] = l_cell_wire[334];							inform_L[423][7] = l_cell_wire[335];							inform_L[296][7] = l_cell_wire[336];							inform_L[424][7] = l_cell_wire[337];							inform_L[297][7] = l_cell_wire[338];							inform_L[425][7] = l_cell_wire[339];							inform_L[298][7] = l_cell_wire[340];							inform_L[426][7] = l_cell_wire[341];							inform_L[299][7] = l_cell_wire[342];							inform_L[427][7] = l_cell_wire[343];							inform_L[300][7] = l_cell_wire[344];							inform_L[428][7] = l_cell_wire[345];							inform_L[301][7] = l_cell_wire[346];							inform_L[429][7] = l_cell_wire[347];							inform_L[302][7] = l_cell_wire[348];							inform_L[430][7] = l_cell_wire[349];							inform_L[303][7] = l_cell_wire[350];							inform_L[431][7] = l_cell_wire[351];							inform_L[304][7] = l_cell_wire[352];							inform_L[432][7] = l_cell_wire[353];							inform_L[305][7] = l_cell_wire[354];							inform_L[433][7] = l_cell_wire[355];							inform_L[306][7] = l_cell_wire[356];							inform_L[434][7] = l_cell_wire[357];							inform_L[307][7] = l_cell_wire[358];							inform_L[435][7] = l_cell_wire[359];							inform_L[308][7] = l_cell_wire[360];							inform_L[436][7] = l_cell_wire[361];							inform_L[309][7] = l_cell_wire[362];							inform_L[437][7] = l_cell_wire[363];							inform_L[310][7] = l_cell_wire[364];							inform_L[438][7] = l_cell_wire[365];							inform_L[311][7] = l_cell_wire[366];							inform_L[439][7] = l_cell_wire[367];							inform_L[312][7] = l_cell_wire[368];							inform_L[440][7] = l_cell_wire[369];							inform_L[313][7] = l_cell_wire[370];							inform_L[441][7] = l_cell_wire[371];							inform_L[314][7] = l_cell_wire[372];							inform_L[442][7] = l_cell_wire[373];							inform_L[315][7] = l_cell_wire[374];							inform_L[443][7] = l_cell_wire[375];							inform_L[316][7] = l_cell_wire[376];							inform_L[444][7] = l_cell_wire[377];							inform_L[317][7] = l_cell_wire[378];							inform_L[445][7] = l_cell_wire[379];							inform_L[318][7] = l_cell_wire[380];							inform_L[446][7] = l_cell_wire[381];							inform_L[319][7] = l_cell_wire[382];							inform_L[447][7] = l_cell_wire[383];							inform_L[320][7] = l_cell_wire[384];							inform_L[448][7] = l_cell_wire[385];							inform_L[321][7] = l_cell_wire[386];							inform_L[449][7] = l_cell_wire[387];							inform_L[322][7] = l_cell_wire[388];							inform_L[450][7] = l_cell_wire[389];							inform_L[323][7] = l_cell_wire[390];							inform_L[451][7] = l_cell_wire[391];							inform_L[324][7] = l_cell_wire[392];							inform_L[452][7] = l_cell_wire[393];							inform_L[325][7] = l_cell_wire[394];							inform_L[453][7] = l_cell_wire[395];							inform_L[326][7] = l_cell_wire[396];							inform_L[454][7] = l_cell_wire[397];							inform_L[327][7] = l_cell_wire[398];							inform_L[455][7] = l_cell_wire[399];							inform_L[328][7] = l_cell_wire[400];							inform_L[456][7] = l_cell_wire[401];							inform_L[329][7] = l_cell_wire[402];							inform_L[457][7] = l_cell_wire[403];							inform_L[330][7] = l_cell_wire[404];							inform_L[458][7] = l_cell_wire[405];							inform_L[331][7] = l_cell_wire[406];							inform_L[459][7] = l_cell_wire[407];							inform_L[332][7] = l_cell_wire[408];							inform_L[460][7] = l_cell_wire[409];							inform_L[333][7] = l_cell_wire[410];							inform_L[461][7] = l_cell_wire[411];							inform_L[334][7] = l_cell_wire[412];							inform_L[462][7] = l_cell_wire[413];							inform_L[335][7] = l_cell_wire[414];							inform_L[463][7] = l_cell_wire[415];							inform_L[336][7] = l_cell_wire[416];							inform_L[464][7] = l_cell_wire[417];							inform_L[337][7] = l_cell_wire[418];							inform_L[465][7] = l_cell_wire[419];							inform_L[338][7] = l_cell_wire[420];							inform_L[466][7] = l_cell_wire[421];							inform_L[339][7] = l_cell_wire[422];							inform_L[467][7] = l_cell_wire[423];							inform_L[340][7] = l_cell_wire[424];							inform_L[468][7] = l_cell_wire[425];							inform_L[341][7] = l_cell_wire[426];							inform_L[469][7] = l_cell_wire[427];							inform_L[342][7] = l_cell_wire[428];							inform_L[470][7] = l_cell_wire[429];							inform_L[343][7] = l_cell_wire[430];							inform_L[471][7] = l_cell_wire[431];							inform_L[344][7] = l_cell_wire[432];							inform_L[472][7] = l_cell_wire[433];							inform_L[345][7] = l_cell_wire[434];							inform_L[473][7] = l_cell_wire[435];							inform_L[346][7] = l_cell_wire[436];							inform_L[474][7] = l_cell_wire[437];							inform_L[347][7] = l_cell_wire[438];							inform_L[475][7] = l_cell_wire[439];							inform_L[348][7] = l_cell_wire[440];							inform_L[476][7] = l_cell_wire[441];							inform_L[349][7] = l_cell_wire[442];							inform_L[477][7] = l_cell_wire[443];							inform_L[350][7] = l_cell_wire[444];							inform_L[478][7] = l_cell_wire[445];							inform_L[351][7] = l_cell_wire[446];							inform_L[479][7] = l_cell_wire[447];							inform_L[352][7] = l_cell_wire[448];							inform_L[480][7] = l_cell_wire[449];							inform_L[353][7] = l_cell_wire[450];							inform_L[481][7] = l_cell_wire[451];							inform_L[354][7] = l_cell_wire[452];							inform_L[482][7] = l_cell_wire[453];							inform_L[355][7] = l_cell_wire[454];							inform_L[483][7] = l_cell_wire[455];							inform_L[356][7] = l_cell_wire[456];							inform_L[484][7] = l_cell_wire[457];							inform_L[357][7] = l_cell_wire[458];							inform_L[485][7] = l_cell_wire[459];							inform_L[358][7] = l_cell_wire[460];							inform_L[486][7] = l_cell_wire[461];							inform_L[359][7] = l_cell_wire[462];							inform_L[487][7] = l_cell_wire[463];							inform_L[360][7] = l_cell_wire[464];							inform_L[488][7] = l_cell_wire[465];							inform_L[361][7] = l_cell_wire[466];							inform_L[489][7] = l_cell_wire[467];							inform_L[362][7] = l_cell_wire[468];							inform_L[490][7] = l_cell_wire[469];							inform_L[363][7] = l_cell_wire[470];							inform_L[491][7] = l_cell_wire[471];							inform_L[364][7] = l_cell_wire[472];							inform_L[492][7] = l_cell_wire[473];							inform_L[365][7] = l_cell_wire[474];							inform_L[493][7] = l_cell_wire[475];							inform_L[366][7] = l_cell_wire[476];							inform_L[494][7] = l_cell_wire[477];							inform_L[367][7] = l_cell_wire[478];							inform_L[495][7] = l_cell_wire[479];							inform_L[368][7] = l_cell_wire[480];							inform_L[496][7] = l_cell_wire[481];							inform_L[369][7] = l_cell_wire[482];							inform_L[497][7] = l_cell_wire[483];							inform_L[370][7] = l_cell_wire[484];							inform_L[498][7] = l_cell_wire[485];							inform_L[371][7] = l_cell_wire[486];							inform_L[499][7] = l_cell_wire[487];							inform_L[372][7] = l_cell_wire[488];							inform_L[500][7] = l_cell_wire[489];							inform_L[373][7] = l_cell_wire[490];							inform_L[501][7] = l_cell_wire[491];							inform_L[374][7] = l_cell_wire[492];							inform_L[502][7] = l_cell_wire[493];							inform_L[375][7] = l_cell_wire[494];							inform_L[503][7] = l_cell_wire[495];							inform_L[376][7] = l_cell_wire[496];							inform_L[504][7] = l_cell_wire[497];							inform_L[377][7] = l_cell_wire[498];							inform_L[505][7] = l_cell_wire[499];							inform_L[378][7] = l_cell_wire[500];							inform_L[506][7] = l_cell_wire[501];							inform_L[379][7] = l_cell_wire[502];							inform_L[507][7] = l_cell_wire[503];							inform_L[380][7] = l_cell_wire[504];							inform_L[508][7] = l_cell_wire[505];							inform_L[381][7] = l_cell_wire[506];							inform_L[509][7] = l_cell_wire[507];							inform_L[382][7] = l_cell_wire[508];							inform_L[510][7] = l_cell_wire[509];							inform_L[383][7] = l_cell_wire[510];							inform_L[511][7] = l_cell_wire[511];							inform_L[512][7] = l_cell_wire[512];							inform_L[640][7] = l_cell_wire[513];							inform_L[513][7] = l_cell_wire[514];							inform_L[641][7] = l_cell_wire[515];							inform_L[514][7] = l_cell_wire[516];							inform_L[642][7] = l_cell_wire[517];							inform_L[515][7] = l_cell_wire[518];							inform_L[643][7] = l_cell_wire[519];							inform_L[516][7] = l_cell_wire[520];							inform_L[644][7] = l_cell_wire[521];							inform_L[517][7] = l_cell_wire[522];							inform_L[645][7] = l_cell_wire[523];							inform_L[518][7] = l_cell_wire[524];							inform_L[646][7] = l_cell_wire[525];							inform_L[519][7] = l_cell_wire[526];							inform_L[647][7] = l_cell_wire[527];							inform_L[520][7] = l_cell_wire[528];							inform_L[648][7] = l_cell_wire[529];							inform_L[521][7] = l_cell_wire[530];							inform_L[649][7] = l_cell_wire[531];							inform_L[522][7] = l_cell_wire[532];							inform_L[650][7] = l_cell_wire[533];							inform_L[523][7] = l_cell_wire[534];							inform_L[651][7] = l_cell_wire[535];							inform_L[524][7] = l_cell_wire[536];							inform_L[652][7] = l_cell_wire[537];							inform_L[525][7] = l_cell_wire[538];							inform_L[653][7] = l_cell_wire[539];							inform_L[526][7] = l_cell_wire[540];							inform_L[654][7] = l_cell_wire[541];							inform_L[527][7] = l_cell_wire[542];							inform_L[655][7] = l_cell_wire[543];							inform_L[528][7] = l_cell_wire[544];							inform_L[656][7] = l_cell_wire[545];							inform_L[529][7] = l_cell_wire[546];							inform_L[657][7] = l_cell_wire[547];							inform_L[530][7] = l_cell_wire[548];							inform_L[658][7] = l_cell_wire[549];							inform_L[531][7] = l_cell_wire[550];							inform_L[659][7] = l_cell_wire[551];							inform_L[532][7] = l_cell_wire[552];							inform_L[660][7] = l_cell_wire[553];							inform_L[533][7] = l_cell_wire[554];							inform_L[661][7] = l_cell_wire[555];							inform_L[534][7] = l_cell_wire[556];							inform_L[662][7] = l_cell_wire[557];							inform_L[535][7] = l_cell_wire[558];							inform_L[663][7] = l_cell_wire[559];							inform_L[536][7] = l_cell_wire[560];							inform_L[664][7] = l_cell_wire[561];							inform_L[537][7] = l_cell_wire[562];							inform_L[665][7] = l_cell_wire[563];							inform_L[538][7] = l_cell_wire[564];							inform_L[666][7] = l_cell_wire[565];							inform_L[539][7] = l_cell_wire[566];							inform_L[667][7] = l_cell_wire[567];							inform_L[540][7] = l_cell_wire[568];							inform_L[668][7] = l_cell_wire[569];							inform_L[541][7] = l_cell_wire[570];							inform_L[669][7] = l_cell_wire[571];							inform_L[542][7] = l_cell_wire[572];							inform_L[670][7] = l_cell_wire[573];							inform_L[543][7] = l_cell_wire[574];							inform_L[671][7] = l_cell_wire[575];							inform_L[544][7] = l_cell_wire[576];							inform_L[672][7] = l_cell_wire[577];							inform_L[545][7] = l_cell_wire[578];							inform_L[673][7] = l_cell_wire[579];							inform_L[546][7] = l_cell_wire[580];							inform_L[674][7] = l_cell_wire[581];							inform_L[547][7] = l_cell_wire[582];							inform_L[675][7] = l_cell_wire[583];							inform_L[548][7] = l_cell_wire[584];							inform_L[676][7] = l_cell_wire[585];							inform_L[549][7] = l_cell_wire[586];							inform_L[677][7] = l_cell_wire[587];							inform_L[550][7] = l_cell_wire[588];							inform_L[678][7] = l_cell_wire[589];							inform_L[551][7] = l_cell_wire[590];							inform_L[679][7] = l_cell_wire[591];							inform_L[552][7] = l_cell_wire[592];							inform_L[680][7] = l_cell_wire[593];							inform_L[553][7] = l_cell_wire[594];							inform_L[681][7] = l_cell_wire[595];							inform_L[554][7] = l_cell_wire[596];							inform_L[682][7] = l_cell_wire[597];							inform_L[555][7] = l_cell_wire[598];							inform_L[683][7] = l_cell_wire[599];							inform_L[556][7] = l_cell_wire[600];							inform_L[684][7] = l_cell_wire[601];							inform_L[557][7] = l_cell_wire[602];							inform_L[685][7] = l_cell_wire[603];							inform_L[558][7] = l_cell_wire[604];							inform_L[686][7] = l_cell_wire[605];							inform_L[559][7] = l_cell_wire[606];							inform_L[687][7] = l_cell_wire[607];							inform_L[560][7] = l_cell_wire[608];							inform_L[688][7] = l_cell_wire[609];							inform_L[561][7] = l_cell_wire[610];							inform_L[689][7] = l_cell_wire[611];							inform_L[562][7] = l_cell_wire[612];							inform_L[690][7] = l_cell_wire[613];							inform_L[563][7] = l_cell_wire[614];							inform_L[691][7] = l_cell_wire[615];							inform_L[564][7] = l_cell_wire[616];							inform_L[692][7] = l_cell_wire[617];							inform_L[565][7] = l_cell_wire[618];							inform_L[693][7] = l_cell_wire[619];							inform_L[566][7] = l_cell_wire[620];							inform_L[694][7] = l_cell_wire[621];							inform_L[567][7] = l_cell_wire[622];							inform_L[695][7] = l_cell_wire[623];							inform_L[568][7] = l_cell_wire[624];							inform_L[696][7] = l_cell_wire[625];							inform_L[569][7] = l_cell_wire[626];							inform_L[697][7] = l_cell_wire[627];							inform_L[570][7] = l_cell_wire[628];							inform_L[698][7] = l_cell_wire[629];							inform_L[571][7] = l_cell_wire[630];							inform_L[699][7] = l_cell_wire[631];							inform_L[572][7] = l_cell_wire[632];							inform_L[700][7] = l_cell_wire[633];							inform_L[573][7] = l_cell_wire[634];							inform_L[701][7] = l_cell_wire[635];							inform_L[574][7] = l_cell_wire[636];							inform_L[702][7] = l_cell_wire[637];							inform_L[575][7] = l_cell_wire[638];							inform_L[703][7] = l_cell_wire[639];							inform_L[576][7] = l_cell_wire[640];							inform_L[704][7] = l_cell_wire[641];							inform_L[577][7] = l_cell_wire[642];							inform_L[705][7] = l_cell_wire[643];							inform_L[578][7] = l_cell_wire[644];							inform_L[706][7] = l_cell_wire[645];							inform_L[579][7] = l_cell_wire[646];							inform_L[707][7] = l_cell_wire[647];							inform_L[580][7] = l_cell_wire[648];							inform_L[708][7] = l_cell_wire[649];							inform_L[581][7] = l_cell_wire[650];							inform_L[709][7] = l_cell_wire[651];							inform_L[582][7] = l_cell_wire[652];							inform_L[710][7] = l_cell_wire[653];							inform_L[583][7] = l_cell_wire[654];							inform_L[711][7] = l_cell_wire[655];							inform_L[584][7] = l_cell_wire[656];							inform_L[712][7] = l_cell_wire[657];							inform_L[585][7] = l_cell_wire[658];							inform_L[713][7] = l_cell_wire[659];							inform_L[586][7] = l_cell_wire[660];							inform_L[714][7] = l_cell_wire[661];							inform_L[587][7] = l_cell_wire[662];							inform_L[715][7] = l_cell_wire[663];							inform_L[588][7] = l_cell_wire[664];							inform_L[716][7] = l_cell_wire[665];							inform_L[589][7] = l_cell_wire[666];							inform_L[717][7] = l_cell_wire[667];							inform_L[590][7] = l_cell_wire[668];							inform_L[718][7] = l_cell_wire[669];							inform_L[591][7] = l_cell_wire[670];							inform_L[719][7] = l_cell_wire[671];							inform_L[592][7] = l_cell_wire[672];							inform_L[720][7] = l_cell_wire[673];							inform_L[593][7] = l_cell_wire[674];							inform_L[721][7] = l_cell_wire[675];							inform_L[594][7] = l_cell_wire[676];							inform_L[722][7] = l_cell_wire[677];							inform_L[595][7] = l_cell_wire[678];							inform_L[723][7] = l_cell_wire[679];							inform_L[596][7] = l_cell_wire[680];							inform_L[724][7] = l_cell_wire[681];							inform_L[597][7] = l_cell_wire[682];							inform_L[725][7] = l_cell_wire[683];							inform_L[598][7] = l_cell_wire[684];							inform_L[726][7] = l_cell_wire[685];							inform_L[599][7] = l_cell_wire[686];							inform_L[727][7] = l_cell_wire[687];							inform_L[600][7] = l_cell_wire[688];							inform_L[728][7] = l_cell_wire[689];							inform_L[601][7] = l_cell_wire[690];							inform_L[729][7] = l_cell_wire[691];							inform_L[602][7] = l_cell_wire[692];							inform_L[730][7] = l_cell_wire[693];							inform_L[603][7] = l_cell_wire[694];							inform_L[731][7] = l_cell_wire[695];							inform_L[604][7] = l_cell_wire[696];							inform_L[732][7] = l_cell_wire[697];							inform_L[605][7] = l_cell_wire[698];							inform_L[733][7] = l_cell_wire[699];							inform_L[606][7] = l_cell_wire[700];							inform_L[734][7] = l_cell_wire[701];							inform_L[607][7] = l_cell_wire[702];							inform_L[735][7] = l_cell_wire[703];							inform_L[608][7] = l_cell_wire[704];							inform_L[736][7] = l_cell_wire[705];							inform_L[609][7] = l_cell_wire[706];							inform_L[737][7] = l_cell_wire[707];							inform_L[610][7] = l_cell_wire[708];							inform_L[738][7] = l_cell_wire[709];							inform_L[611][7] = l_cell_wire[710];							inform_L[739][7] = l_cell_wire[711];							inform_L[612][7] = l_cell_wire[712];							inform_L[740][7] = l_cell_wire[713];							inform_L[613][7] = l_cell_wire[714];							inform_L[741][7] = l_cell_wire[715];							inform_L[614][7] = l_cell_wire[716];							inform_L[742][7] = l_cell_wire[717];							inform_L[615][7] = l_cell_wire[718];							inform_L[743][7] = l_cell_wire[719];							inform_L[616][7] = l_cell_wire[720];							inform_L[744][7] = l_cell_wire[721];							inform_L[617][7] = l_cell_wire[722];							inform_L[745][7] = l_cell_wire[723];							inform_L[618][7] = l_cell_wire[724];							inform_L[746][7] = l_cell_wire[725];							inform_L[619][7] = l_cell_wire[726];							inform_L[747][7] = l_cell_wire[727];							inform_L[620][7] = l_cell_wire[728];							inform_L[748][7] = l_cell_wire[729];							inform_L[621][7] = l_cell_wire[730];							inform_L[749][7] = l_cell_wire[731];							inform_L[622][7] = l_cell_wire[732];							inform_L[750][7] = l_cell_wire[733];							inform_L[623][7] = l_cell_wire[734];							inform_L[751][7] = l_cell_wire[735];							inform_L[624][7] = l_cell_wire[736];							inform_L[752][7] = l_cell_wire[737];							inform_L[625][7] = l_cell_wire[738];							inform_L[753][7] = l_cell_wire[739];							inform_L[626][7] = l_cell_wire[740];							inform_L[754][7] = l_cell_wire[741];							inform_L[627][7] = l_cell_wire[742];							inform_L[755][7] = l_cell_wire[743];							inform_L[628][7] = l_cell_wire[744];							inform_L[756][7] = l_cell_wire[745];							inform_L[629][7] = l_cell_wire[746];							inform_L[757][7] = l_cell_wire[747];							inform_L[630][7] = l_cell_wire[748];							inform_L[758][7] = l_cell_wire[749];							inform_L[631][7] = l_cell_wire[750];							inform_L[759][7] = l_cell_wire[751];							inform_L[632][7] = l_cell_wire[752];							inform_L[760][7] = l_cell_wire[753];							inform_L[633][7] = l_cell_wire[754];							inform_L[761][7] = l_cell_wire[755];							inform_L[634][7] = l_cell_wire[756];							inform_L[762][7] = l_cell_wire[757];							inform_L[635][7] = l_cell_wire[758];							inform_L[763][7] = l_cell_wire[759];							inform_L[636][7] = l_cell_wire[760];							inform_L[764][7] = l_cell_wire[761];							inform_L[637][7] = l_cell_wire[762];							inform_L[765][7] = l_cell_wire[763];							inform_L[638][7] = l_cell_wire[764];							inform_L[766][7] = l_cell_wire[765];							inform_L[639][7] = l_cell_wire[766];							inform_L[767][7] = l_cell_wire[767];							inform_L[768][7] = l_cell_wire[768];							inform_L[896][7] = l_cell_wire[769];							inform_L[769][7] = l_cell_wire[770];							inform_L[897][7] = l_cell_wire[771];							inform_L[770][7] = l_cell_wire[772];							inform_L[898][7] = l_cell_wire[773];							inform_L[771][7] = l_cell_wire[774];							inform_L[899][7] = l_cell_wire[775];							inform_L[772][7] = l_cell_wire[776];							inform_L[900][7] = l_cell_wire[777];							inform_L[773][7] = l_cell_wire[778];							inform_L[901][7] = l_cell_wire[779];							inform_L[774][7] = l_cell_wire[780];							inform_L[902][7] = l_cell_wire[781];							inform_L[775][7] = l_cell_wire[782];							inform_L[903][7] = l_cell_wire[783];							inform_L[776][7] = l_cell_wire[784];							inform_L[904][7] = l_cell_wire[785];							inform_L[777][7] = l_cell_wire[786];							inform_L[905][7] = l_cell_wire[787];							inform_L[778][7] = l_cell_wire[788];							inform_L[906][7] = l_cell_wire[789];							inform_L[779][7] = l_cell_wire[790];							inform_L[907][7] = l_cell_wire[791];							inform_L[780][7] = l_cell_wire[792];							inform_L[908][7] = l_cell_wire[793];							inform_L[781][7] = l_cell_wire[794];							inform_L[909][7] = l_cell_wire[795];							inform_L[782][7] = l_cell_wire[796];							inform_L[910][7] = l_cell_wire[797];							inform_L[783][7] = l_cell_wire[798];							inform_L[911][7] = l_cell_wire[799];							inform_L[784][7] = l_cell_wire[800];							inform_L[912][7] = l_cell_wire[801];							inform_L[785][7] = l_cell_wire[802];							inform_L[913][7] = l_cell_wire[803];							inform_L[786][7] = l_cell_wire[804];							inform_L[914][7] = l_cell_wire[805];							inform_L[787][7] = l_cell_wire[806];							inform_L[915][7] = l_cell_wire[807];							inform_L[788][7] = l_cell_wire[808];							inform_L[916][7] = l_cell_wire[809];							inform_L[789][7] = l_cell_wire[810];							inform_L[917][7] = l_cell_wire[811];							inform_L[790][7] = l_cell_wire[812];							inform_L[918][7] = l_cell_wire[813];							inform_L[791][7] = l_cell_wire[814];							inform_L[919][7] = l_cell_wire[815];							inform_L[792][7] = l_cell_wire[816];							inform_L[920][7] = l_cell_wire[817];							inform_L[793][7] = l_cell_wire[818];							inform_L[921][7] = l_cell_wire[819];							inform_L[794][7] = l_cell_wire[820];							inform_L[922][7] = l_cell_wire[821];							inform_L[795][7] = l_cell_wire[822];							inform_L[923][7] = l_cell_wire[823];							inform_L[796][7] = l_cell_wire[824];							inform_L[924][7] = l_cell_wire[825];							inform_L[797][7] = l_cell_wire[826];							inform_L[925][7] = l_cell_wire[827];							inform_L[798][7] = l_cell_wire[828];							inform_L[926][7] = l_cell_wire[829];							inform_L[799][7] = l_cell_wire[830];							inform_L[927][7] = l_cell_wire[831];							inform_L[800][7] = l_cell_wire[832];							inform_L[928][7] = l_cell_wire[833];							inform_L[801][7] = l_cell_wire[834];							inform_L[929][7] = l_cell_wire[835];							inform_L[802][7] = l_cell_wire[836];							inform_L[930][7] = l_cell_wire[837];							inform_L[803][7] = l_cell_wire[838];							inform_L[931][7] = l_cell_wire[839];							inform_L[804][7] = l_cell_wire[840];							inform_L[932][7] = l_cell_wire[841];							inform_L[805][7] = l_cell_wire[842];							inform_L[933][7] = l_cell_wire[843];							inform_L[806][7] = l_cell_wire[844];							inform_L[934][7] = l_cell_wire[845];							inform_L[807][7] = l_cell_wire[846];							inform_L[935][7] = l_cell_wire[847];							inform_L[808][7] = l_cell_wire[848];							inform_L[936][7] = l_cell_wire[849];							inform_L[809][7] = l_cell_wire[850];							inform_L[937][7] = l_cell_wire[851];							inform_L[810][7] = l_cell_wire[852];							inform_L[938][7] = l_cell_wire[853];							inform_L[811][7] = l_cell_wire[854];							inform_L[939][7] = l_cell_wire[855];							inform_L[812][7] = l_cell_wire[856];							inform_L[940][7] = l_cell_wire[857];							inform_L[813][7] = l_cell_wire[858];							inform_L[941][7] = l_cell_wire[859];							inform_L[814][7] = l_cell_wire[860];							inform_L[942][7] = l_cell_wire[861];							inform_L[815][7] = l_cell_wire[862];							inform_L[943][7] = l_cell_wire[863];							inform_L[816][7] = l_cell_wire[864];							inform_L[944][7] = l_cell_wire[865];							inform_L[817][7] = l_cell_wire[866];							inform_L[945][7] = l_cell_wire[867];							inform_L[818][7] = l_cell_wire[868];							inform_L[946][7] = l_cell_wire[869];							inform_L[819][7] = l_cell_wire[870];							inform_L[947][7] = l_cell_wire[871];							inform_L[820][7] = l_cell_wire[872];							inform_L[948][7] = l_cell_wire[873];							inform_L[821][7] = l_cell_wire[874];							inform_L[949][7] = l_cell_wire[875];							inform_L[822][7] = l_cell_wire[876];							inform_L[950][7] = l_cell_wire[877];							inform_L[823][7] = l_cell_wire[878];							inform_L[951][7] = l_cell_wire[879];							inform_L[824][7] = l_cell_wire[880];							inform_L[952][7] = l_cell_wire[881];							inform_L[825][7] = l_cell_wire[882];							inform_L[953][7] = l_cell_wire[883];							inform_L[826][7] = l_cell_wire[884];							inform_L[954][7] = l_cell_wire[885];							inform_L[827][7] = l_cell_wire[886];							inform_L[955][7] = l_cell_wire[887];							inform_L[828][7] = l_cell_wire[888];							inform_L[956][7] = l_cell_wire[889];							inform_L[829][7] = l_cell_wire[890];							inform_L[957][7] = l_cell_wire[891];							inform_L[830][7] = l_cell_wire[892];							inform_L[958][7] = l_cell_wire[893];							inform_L[831][7] = l_cell_wire[894];							inform_L[959][7] = l_cell_wire[895];							inform_L[832][7] = l_cell_wire[896];							inform_L[960][7] = l_cell_wire[897];							inform_L[833][7] = l_cell_wire[898];							inform_L[961][7] = l_cell_wire[899];							inform_L[834][7] = l_cell_wire[900];							inform_L[962][7] = l_cell_wire[901];							inform_L[835][7] = l_cell_wire[902];							inform_L[963][7] = l_cell_wire[903];							inform_L[836][7] = l_cell_wire[904];							inform_L[964][7] = l_cell_wire[905];							inform_L[837][7] = l_cell_wire[906];							inform_L[965][7] = l_cell_wire[907];							inform_L[838][7] = l_cell_wire[908];							inform_L[966][7] = l_cell_wire[909];							inform_L[839][7] = l_cell_wire[910];							inform_L[967][7] = l_cell_wire[911];							inform_L[840][7] = l_cell_wire[912];							inform_L[968][7] = l_cell_wire[913];							inform_L[841][7] = l_cell_wire[914];							inform_L[969][7] = l_cell_wire[915];							inform_L[842][7] = l_cell_wire[916];							inform_L[970][7] = l_cell_wire[917];							inform_L[843][7] = l_cell_wire[918];							inform_L[971][7] = l_cell_wire[919];							inform_L[844][7] = l_cell_wire[920];							inform_L[972][7] = l_cell_wire[921];							inform_L[845][7] = l_cell_wire[922];							inform_L[973][7] = l_cell_wire[923];							inform_L[846][7] = l_cell_wire[924];							inform_L[974][7] = l_cell_wire[925];							inform_L[847][7] = l_cell_wire[926];							inform_L[975][7] = l_cell_wire[927];							inform_L[848][7] = l_cell_wire[928];							inform_L[976][7] = l_cell_wire[929];							inform_L[849][7] = l_cell_wire[930];							inform_L[977][7] = l_cell_wire[931];							inform_L[850][7] = l_cell_wire[932];							inform_L[978][7] = l_cell_wire[933];							inform_L[851][7] = l_cell_wire[934];							inform_L[979][7] = l_cell_wire[935];							inform_L[852][7] = l_cell_wire[936];							inform_L[980][7] = l_cell_wire[937];							inform_L[853][7] = l_cell_wire[938];							inform_L[981][7] = l_cell_wire[939];							inform_L[854][7] = l_cell_wire[940];							inform_L[982][7] = l_cell_wire[941];							inform_L[855][7] = l_cell_wire[942];							inform_L[983][7] = l_cell_wire[943];							inform_L[856][7] = l_cell_wire[944];							inform_L[984][7] = l_cell_wire[945];							inform_L[857][7] = l_cell_wire[946];							inform_L[985][7] = l_cell_wire[947];							inform_L[858][7] = l_cell_wire[948];							inform_L[986][7] = l_cell_wire[949];							inform_L[859][7] = l_cell_wire[950];							inform_L[987][7] = l_cell_wire[951];							inform_L[860][7] = l_cell_wire[952];							inform_L[988][7] = l_cell_wire[953];							inform_L[861][7] = l_cell_wire[954];							inform_L[989][7] = l_cell_wire[955];							inform_L[862][7] = l_cell_wire[956];							inform_L[990][7] = l_cell_wire[957];							inform_L[863][7] = l_cell_wire[958];							inform_L[991][7] = l_cell_wire[959];							inform_L[864][7] = l_cell_wire[960];							inform_L[992][7] = l_cell_wire[961];							inform_L[865][7] = l_cell_wire[962];							inform_L[993][7] = l_cell_wire[963];							inform_L[866][7] = l_cell_wire[964];							inform_L[994][7] = l_cell_wire[965];							inform_L[867][7] = l_cell_wire[966];							inform_L[995][7] = l_cell_wire[967];							inform_L[868][7] = l_cell_wire[968];							inform_L[996][7] = l_cell_wire[969];							inform_L[869][7] = l_cell_wire[970];							inform_L[997][7] = l_cell_wire[971];							inform_L[870][7] = l_cell_wire[972];							inform_L[998][7] = l_cell_wire[973];							inform_L[871][7] = l_cell_wire[974];							inform_L[999][7] = l_cell_wire[975];							inform_L[872][7] = l_cell_wire[976];							inform_L[1000][7] = l_cell_wire[977];							inform_L[873][7] = l_cell_wire[978];							inform_L[1001][7] = l_cell_wire[979];							inform_L[874][7] = l_cell_wire[980];							inform_L[1002][7] = l_cell_wire[981];							inform_L[875][7] = l_cell_wire[982];							inform_L[1003][7] = l_cell_wire[983];							inform_L[876][7] = l_cell_wire[984];							inform_L[1004][7] = l_cell_wire[985];							inform_L[877][7] = l_cell_wire[986];							inform_L[1005][7] = l_cell_wire[987];							inform_L[878][7] = l_cell_wire[988];							inform_L[1006][7] = l_cell_wire[989];							inform_L[879][7] = l_cell_wire[990];							inform_L[1007][7] = l_cell_wire[991];							inform_L[880][7] = l_cell_wire[992];							inform_L[1008][7] = l_cell_wire[993];							inform_L[881][7] = l_cell_wire[994];							inform_L[1009][7] = l_cell_wire[995];							inform_L[882][7] = l_cell_wire[996];							inform_L[1010][7] = l_cell_wire[997];							inform_L[883][7] = l_cell_wire[998];							inform_L[1011][7] = l_cell_wire[999];							inform_L[884][7] = l_cell_wire[1000];							inform_L[1012][7] = l_cell_wire[1001];							inform_L[885][7] = l_cell_wire[1002];							inform_L[1013][7] = l_cell_wire[1003];							inform_L[886][7] = l_cell_wire[1004];							inform_L[1014][7] = l_cell_wire[1005];							inform_L[887][7] = l_cell_wire[1006];							inform_L[1015][7] = l_cell_wire[1007];							inform_L[888][7] = l_cell_wire[1008];							inform_L[1016][7] = l_cell_wire[1009];							inform_L[889][7] = l_cell_wire[1010];							inform_L[1017][7] = l_cell_wire[1011];							inform_L[890][7] = l_cell_wire[1012];							inform_L[1018][7] = l_cell_wire[1013];							inform_L[891][7] = l_cell_wire[1014];							inform_L[1019][7] = l_cell_wire[1015];							inform_L[892][7] = l_cell_wire[1016];							inform_L[1020][7] = l_cell_wire[1017];							inform_L[893][7] = l_cell_wire[1018];							inform_L[1021][7] = l_cell_wire[1019];							inform_L[894][7] = l_cell_wire[1020];							inform_L[1022][7] = l_cell_wire[1021];							inform_L[895][7] = l_cell_wire[1022];							inform_L[1023][7] = l_cell_wire[1023];						end
						9:						begin							inform_R[0][9] = r_cell_wire[0];							inform_R[256][9] = r_cell_wire[1];							inform_R[1][9] = r_cell_wire[2];							inform_R[257][9] = r_cell_wire[3];							inform_R[2][9] = r_cell_wire[4];							inform_R[258][9] = r_cell_wire[5];							inform_R[3][9] = r_cell_wire[6];							inform_R[259][9] = r_cell_wire[7];							inform_R[4][9] = r_cell_wire[8];							inform_R[260][9] = r_cell_wire[9];							inform_R[5][9] = r_cell_wire[10];							inform_R[261][9] = r_cell_wire[11];							inform_R[6][9] = r_cell_wire[12];							inform_R[262][9] = r_cell_wire[13];							inform_R[7][9] = r_cell_wire[14];							inform_R[263][9] = r_cell_wire[15];							inform_R[8][9] = r_cell_wire[16];							inform_R[264][9] = r_cell_wire[17];							inform_R[9][9] = r_cell_wire[18];							inform_R[265][9] = r_cell_wire[19];							inform_R[10][9] = r_cell_wire[20];							inform_R[266][9] = r_cell_wire[21];							inform_R[11][9] = r_cell_wire[22];							inform_R[267][9] = r_cell_wire[23];							inform_R[12][9] = r_cell_wire[24];							inform_R[268][9] = r_cell_wire[25];							inform_R[13][9] = r_cell_wire[26];							inform_R[269][9] = r_cell_wire[27];							inform_R[14][9] = r_cell_wire[28];							inform_R[270][9] = r_cell_wire[29];							inform_R[15][9] = r_cell_wire[30];							inform_R[271][9] = r_cell_wire[31];							inform_R[16][9] = r_cell_wire[32];							inform_R[272][9] = r_cell_wire[33];							inform_R[17][9] = r_cell_wire[34];							inform_R[273][9] = r_cell_wire[35];							inform_R[18][9] = r_cell_wire[36];							inform_R[274][9] = r_cell_wire[37];							inform_R[19][9] = r_cell_wire[38];							inform_R[275][9] = r_cell_wire[39];							inform_R[20][9] = r_cell_wire[40];							inform_R[276][9] = r_cell_wire[41];							inform_R[21][9] = r_cell_wire[42];							inform_R[277][9] = r_cell_wire[43];							inform_R[22][9] = r_cell_wire[44];							inform_R[278][9] = r_cell_wire[45];							inform_R[23][9] = r_cell_wire[46];							inform_R[279][9] = r_cell_wire[47];							inform_R[24][9] = r_cell_wire[48];							inform_R[280][9] = r_cell_wire[49];							inform_R[25][9] = r_cell_wire[50];							inform_R[281][9] = r_cell_wire[51];							inform_R[26][9] = r_cell_wire[52];							inform_R[282][9] = r_cell_wire[53];							inform_R[27][9] = r_cell_wire[54];							inform_R[283][9] = r_cell_wire[55];							inform_R[28][9] = r_cell_wire[56];							inform_R[284][9] = r_cell_wire[57];							inform_R[29][9] = r_cell_wire[58];							inform_R[285][9] = r_cell_wire[59];							inform_R[30][9] = r_cell_wire[60];							inform_R[286][9] = r_cell_wire[61];							inform_R[31][9] = r_cell_wire[62];							inform_R[287][9] = r_cell_wire[63];							inform_R[32][9] = r_cell_wire[64];							inform_R[288][9] = r_cell_wire[65];							inform_R[33][9] = r_cell_wire[66];							inform_R[289][9] = r_cell_wire[67];							inform_R[34][9] = r_cell_wire[68];							inform_R[290][9] = r_cell_wire[69];							inform_R[35][9] = r_cell_wire[70];							inform_R[291][9] = r_cell_wire[71];							inform_R[36][9] = r_cell_wire[72];							inform_R[292][9] = r_cell_wire[73];							inform_R[37][9] = r_cell_wire[74];							inform_R[293][9] = r_cell_wire[75];							inform_R[38][9] = r_cell_wire[76];							inform_R[294][9] = r_cell_wire[77];							inform_R[39][9] = r_cell_wire[78];							inform_R[295][9] = r_cell_wire[79];							inform_R[40][9] = r_cell_wire[80];							inform_R[296][9] = r_cell_wire[81];							inform_R[41][9] = r_cell_wire[82];							inform_R[297][9] = r_cell_wire[83];							inform_R[42][9] = r_cell_wire[84];							inform_R[298][9] = r_cell_wire[85];							inform_R[43][9] = r_cell_wire[86];							inform_R[299][9] = r_cell_wire[87];							inform_R[44][9] = r_cell_wire[88];							inform_R[300][9] = r_cell_wire[89];							inform_R[45][9] = r_cell_wire[90];							inform_R[301][9] = r_cell_wire[91];							inform_R[46][9] = r_cell_wire[92];							inform_R[302][9] = r_cell_wire[93];							inform_R[47][9] = r_cell_wire[94];							inform_R[303][9] = r_cell_wire[95];							inform_R[48][9] = r_cell_wire[96];							inform_R[304][9] = r_cell_wire[97];							inform_R[49][9] = r_cell_wire[98];							inform_R[305][9] = r_cell_wire[99];							inform_R[50][9] = r_cell_wire[100];							inform_R[306][9] = r_cell_wire[101];							inform_R[51][9] = r_cell_wire[102];							inform_R[307][9] = r_cell_wire[103];							inform_R[52][9] = r_cell_wire[104];							inform_R[308][9] = r_cell_wire[105];							inform_R[53][9] = r_cell_wire[106];							inform_R[309][9] = r_cell_wire[107];							inform_R[54][9] = r_cell_wire[108];							inform_R[310][9] = r_cell_wire[109];							inform_R[55][9] = r_cell_wire[110];							inform_R[311][9] = r_cell_wire[111];							inform_R[56][9] = r_cell_wire[112];							inform_R[312][9] = r_cell_wire[113];							inform_R[57][9] = r_cell_wire[114];							inform_R[313][9] = r_cell_wire[115];							inform_R[58][9] = r_cell_wire[116];							inform_R[314][9] = r_cell_wire[117];							inform_R[59][9] = r_cell_wire[118];							inform_R[315][9] = r_cell_wire[119];							inform_R[60][9] = r_cell_wire[120];							inform_R[316][9] = r_cell_wire[121];							inform_R[61][9] = r_cell_wire[122];							inform_R[317][9] = r_cell_wire[123];							inform_R[62][9] = r_cell_wire[124];							inform_R[318][9] = r_cell_wire[125];							inform_R[63][9] = r_cell_wire[126];							inform_R[319][9] = r_cell_wire[127];							inform_R[64][9] = r_cell_wire[128];							inform_R[320][9] = r_cell_wire[129];							inform_R[65][9] = r_cell_wire[130];							inform_R[321][9] = r_cell_wire[131];							inform_R[66][9] = r_cell_wire[132];							inform_R[322][9] = r_cell_wire[133];							inform_R[67][9] = r_cell_wire[134];							inform_R[323][9] = r_cell_wire[135];							inform_R[68][9] = r_cell_wire[136];							inform_R[324][9] = r_cell_wire[137];							inform_R[69][9] = r_cell_wire[138];							inform_R[325][9] = r_cell_wire[139];							inform_R[70][9] = r_cell_wire[140];							inform_R[326][9] = r_cell_wire[141];							inform_R[71][9] = r_cell_wire[142];							inform_R[327][9] = r_cell_wire[143];							inform_R[72][9] = r_cell_wire[144];							inform_R[328][9] = r_cell_wire[145];							inform_R[73][9] = r_cell_wire[146];							inform_R[329][9] = r_cell_wire[147];							inform_R[74][9] = r_cell_wire[148];							inform_R[330][9] = r_cell_wire[149];							inform_R[75][9] = r_cell_wire[150];							inform_R[331][9] = r_cell_wire[151];							inform_R[76][9] = r_cell_wire[152];							inform_R[332][9] = r_cell_wire[153];							inform_R[77][9] = r_cell_wire[154];							inform_R[333][9] = r_cell_wire[155];							inform_R[78][9] = r_cell_wire[156];							inform_R[334][9] = r_cell_wire[157];							inform_R[79][9] = r_cell_wire[158];							inform_R[335][9] = r_cell_wire[159];							inform_R[80][9] = r_cell_wire[160];							inform_R[336][9] = r_cell_wire[161];							inform_R[81][9] = r_cell_wire[162];							inform_R[337][9] = r_cell_wire[163];							inform_R[82][9] = r_cell_wire[164];							inform_R[338][9] = r_cell_wire[165];							inform_R[83][9] = r_cell_wire[166];							inform_R[339][9] = r_cell_wire[167];							inform_R[84][9] = r_cell_wire[168];							inform_R[340][9] = r_cell_wire[169];							inform_R[85][9] = r_cell_wire[170];							inform_R[341][9] = r_cell_wire[171];							inform_R[86][9] = r_cell_wire[172];							inform_R[342][9] = r_cell_wire[173];							inform_R[87][9] = r_cell_wire[174];							inform_R[343][9] = r_cell_wire[175];							inform_R[88][9] = r_cell_wire[176];							inform_R[344][9] = r_cell_wire[177];							inform_R[89][9] = r_cell_wire[178];							inform_R[345][9] = r_cell_wire[179];							inform_R[90][9] = r_cell_wire[180];							inform_R[346][9] = r_cell_wire[181];							inform_R[91][9] = r_cell_wire[182];							inform_R[347][9] = r_cell_wire[183];							inform_R[92][9] = r_cell_wire[184];							inform_R[348][9] = r_cell_wire[185];							inform_R[93][9] = r_cell_wire[186];							inform_R[349][9] = r_cell_wire[187];							inform_R[94][9] = r_cell_wire[188];							inform_R[350][9] = r_cell_wire[189];							inform_R[95][9] = r_cell_wire[190];							inform_R[351][9] = r_cell_wire[191];							inform_R[96][9] = r_cell_wire[192];							inform_R[352][9] = r_cell_wire[193];							inform_R[97][9] = r_cell_wire[194];							inform_R[353][9] = r_cell_wire[195];							inform_R[98][9] = r_cell_wire[196];							inform_R[354][9] = r_cell_wire[197];							inform_R[99][9] = r_cell_wire[198];							inform_R[355][9] = r_cell_wire[199];							inform_R[100][9] = r_cell_wire[200];							inform_R[356][9] = r_cell_wire[201];							inform_R[101][9] = r_cell_wire[202];							inform_R[357][9] = r_cell_wire[203];							inform_R[102][9] = r_cell_wire[204];							inform_R[358][9] = r_cell_wire[205];							inform_R[103][9] = r_cell_wire[206];							inform_R[359][9] = r_cell_wire[207];							inform_R[104][9] = r_cell_wire[208];							inform_R[360][9] = r_cell_wire[209];							inform_R[105][9] = r_cell_wire[210];							inform_R[361][9] = r_cell_wire[211];							inform_R[106][9] = r_cell_wire[212];							inform_R[362][9] = r_cell_wire[213];							inform_R[107][9] = r_cell_wire[214];							inform_R[363][9] = r_cell_wire[215];							inform_R[108][9] = r_cell_wire[216];							inform_R[364][9] = r_cell_wire[217];							inform_R[109][9] = r_cell_wire[218];							inform_R[365][9] = r_cell_wire[219];							inform_R[110][9] = r_cell_wire[220];							inform_R[366][9] = r_cell_wire[221];							inform_R[111][9] = r_cell_wire[222];							inform_R[367][9] = r_cell_wire[223];							inform_R[112][9] = r_cell_wire[224];							inform_R[368][9] = r_cell_wire[225];							inform_R[113][9] = r_cell_wire[226];							inform_R[369][9] = r_cell_wire[227];							inform_R[114][9] = r_cell_wire[228];							inform_R[370][9] = r_cell_wire[229];							inform_R[115][9] = r_cell_wire[230];							inform_R[371][9] = r_cell_wire[231];							inform_R[116][9] = r_cell_wire[232];							inform_R[372][9] = r_cell_wire[233];							inform_R[117][9] = r_cell_wire[234];							inform_R[373][9] = r_cell_wire[235];							inform_R[118][9] = r_cell_wire[236];							inform_R[374][9] = r_cell_wire[237];							inform_R[119][9] = r_cell_wire[238];							inform_R[375][9] = r_cell_wire[239];							inform_R[120][9] = r_cell_wire[240];							inform_R[376][9] = r_cell_wire[241];							inform_R[121][9] = r_cell_wire[242];							inform_R[377][9] = r_cell_wire[243];							inform_R[122][9] = r_cell_wire[244];							inform_R[378][9] = r_cell_wire[245];							inform_R[123][9] = r_cell_wire[246];							inform_R[379][9] = r_cell_wire[247];							inform_R[124][9] = r_cell_wire[248];							inform_R[380][9] = r_cell_wire[249];							inform_R[125][9] = r_cell_wire[250];							inform_R[381][9] = r_cell_wire[251];							inform_R[126][9] = r_cell_wire[252];							inform_R[382][9] = r_cell_wire[253];							inform_R[127][9] = r_cell_wire[254];							inform_R[383][9] = r_cell_wire[255];							inform_R[128][9] = r_cell_wire[256];							inform_R[384][9] = r_cell_wire[257];							inform_R[129][9] = r_cell_wire[258];							inform_R[385][9] = r_cell_wire[259];							inform_R[130][9] = r_cell_wire[260];							inform_R[386][9] = r_cell_wire[261];							inform_R[131][9] = r_cell_wire[262];							inform_R[387][9] = r_cell_wire[263];							inform_R[132][9] = r_cell_wire[264];							inform_R[388][9] = r_cell_wire[265];							inform_R[133][9] = r_cell_wire[266];							inform_R[389][9] = r_cell_wire[267];							inform_R[134][9] = r_cell_wire[268];							inform_R[390][9] = r_cell_wire[269];							inform_R[135][9] = r_cell_wire[270];							inform_R[391][9] = r_cell_wire[271];							inform_R[136][9] = r_cell_wire[272];							inform_R[392][9] = r_cell_wire[273];							inform_R[137][9] = r_cell_wire[274];							inform_R[393][9] = r_cell_wire[275];							inform_R[138][9] = r_cell_wire[276];							inform_R[394][9] = r_cell_wire[277];							inform_R[139][9] = r_cell_wire[278];							inform_R[395][9] = r_cell_wire[279];							inform_R[140][9] = r_cell_wire[280];							inform_R[396][9] = r_cell_wire[281];							inform_R[141][9] = r_cell_wire[282];							inform_R[397][9] = r_cell_wire[283];							inform_R[142][9] = r_cell_wire[284];							inform_R[398][9] = r_cell_wire[285];							inform_R[143][9] = r_cell_wire[286];							inform_R[399][9] = r_cell_wire[287];							inform_R[144][9] = r_cell_wire[288];							inform_R[400][9] = r_cell_wire[289];							inform_R[145][9] = r_cell_wire[290];							inform_R[401][9] = r_cell_wire[291];							inform_R[146][9] = r_cell_wire[292];							inform_R[402][9] = r_cell_wire[293];							inform_R[147][9] = r_cell_wire[294];							inform_R[403][9] = r_cell_wire[295];							inform_R[148][9] = r_cell_wire[296];							inform_R[404][9] = r_cell_wire[297];							inform_R[149][9] = r_cell_wire[298];							inform_R[405][9] = r_cell_wire[299];							inform_R[150][9] = r_cell_wire[300];							inform_R[406][9] = r_cell_wire[301];							inform_R[151][9] = r_cell_wire[302];							inform_R[407][9] = r_cell_wire[303];							inform_R[152][9] = r_cell_wire[304];							inform_R[408][9] = r_cell_wire[305];							inform_R[153][9] = r_cell_wire[306];							inform_R[409][9] = r_cell_wire[307];							inform_R[154][9] = r_cell_wire[308];							inform_R[410][9] = r_cell_wire[309];							inform_R[155][9] = r_cell_wire[310];							inform_R[411][9] = r_cell_wire[311];							inform_R[156][9] = r_cell_wire[312];							inform_R[412][9] = r_cell_wire[313];							inform_R[157][9] = r_cell_wire[314];							inform_R[413][9] = r_cell_wire[315];							inform_R[158][9] = r_cell_wire[316];							inform_R[414][9] = r_cell_wire[317];							inform_R[159][9] = r_cell_wire[318];							inform_R[415][9] = r_cell_wire[319];							inform_R[160][9] = r_cell_wire[320];							inform_R[416][9] = r_cell_wire[321];							inform_R[161][9] = r_cell_wire[322];							inform_R[417][9] = r_cell_wire[323];							inform_R[162][9] = r_cell_wire[324];							inform_R[418][9] = r_cell_wire[325];							inform_R[163][9] = r_cell_wire[326];							inform_R[419][9] = r_cell_wire[327];							inform_R[164][9] = r_cell_wire[328];							inform_R[420][9] = r_cell_wire[329];							inform_R[165][9] = r_cell_wire[330];							inform_R[421][9] = r_cell_wire[331];							inform_R[166][9] = r_cell_wire[332];							inform_R[422][9] = r_cell_wire[333];							inform_R[167][9] = r_cell_wire[334];							inform_R[423][9] = r_cell_wire[335];							inform_R[168][9] = r_cell_wire[336];							inform_R[424][9] = r_cell_wire[337];							inform_R[169][9] = r_cell_wire[338];							inform_R[425][9] = r_cell_wire[339];							inform_R[170][9] = r_cell_wire[340];							inform_R[426][9] = r_cell_wire[341];							inform_R[171][9] = r_cell_wire[342];							inform_R[427][9] = r_cell_wire[343];							inform_R[172][9] = r_cell_wire[344];							inform_R[428][9] = r_cell_wire[345];							inform_R[173][9] = r_cell_wire[346];							inform_R[429][9] = r_cell_wire[347];							inform_R[174][9] = r_cell_wire[348];							inform_R[430][9] = r_cell_wire[349];							inform_R[175][9] = r_cell_wire[350];							inform_R[431][9] = r_cell_wire[351];							inform_R[176][9] = r_cell_wire[352];							inform_R[432][9] = r_cell_wire[353];							inform_R[177][9] = r_cell_wire[354];							inform_R[433][9] = r_cell_wire[355];							inform_R[178][9] = r_cell_wire[356];							inform_R[434][9] = r_cell_wire[357];							inform_R[179][9] = r_cell_wire[358];							inform_R[435][9] = r_cell_wire[359];							inform_R[180][9] = r_cell_wire[360];							inform_R[436][9] = r_cell_wire[361];							inform_R[181][9] = r_cell_wire[362];							inform_R[437][9] = r_cell_wire[363];							inform_R[182][9] = r_cell_wire[364];							inform_R[438][9] = r_cell_wire[365];							inform_R[183][9] = r_cell_wire[366];							inform_R[439][9] = r_cell_wire[367];							inform_R[184][9] = r_cell_wire[368];							inform_R[440][9] = r_cell_wire[369];							inform_R[185][9] = r_cell_wire[370];							inform_R[441][9] = r_cell_wire[371];							inform_R[186][9] = r_cell_wire[372];							inform_R[442][9] = r_cell_wire[373];							inform_R[187][9] = r_cell_wire[374];							inform_R[443][9] = r_cell_wire[375];							inform_R[188][9] = r_cell_wire[376];							inform_R[444][9] = r_cell_wire[377];							inform_R[189][9] = r_cell_wire[378];							inform_R[445][9] = r_cell_wire[379];							inform_R[190][9] = r_cell_wire[380];							inform_R[446][9] = r_cell_wire[381];							inform_R[191][9] = r_cell_wire[382];							inform_R[447][9] = r_cell_wire[383];							inform_R[192][9] = r_cell_wire[384];							inform_R[448][9] = r_cell_wire[385];							inform_R[193][9] = r_cell_wire[386];							inform_R[449][9] = r_cell_wire[387];							inform_R[194][9] = r_cell_wire[388];							inform_R[450][9] = r_cell_wire[389];							inform_R[195][9] = r_cell_wire[390];							inform_R[451][9] = r_cell_wire[391];							inform_R[196][9] = r_cell_wire[392];							inform_R[452][9] = r_cell_wire[393];							inform_R[197][9] = r_cell_wire[394];							inform_R[453][9] = r_cell_wire[395];							inform_R[198][9] = r_cell_wire[396];							inform_R[454][9] = r_cell_wire[397];							inform_R[199][9] = r_cell_wire[398];							inform_R[455][9] = r_cell_wire[399];							inform_R[200][9] = r_cell_wire[400];							inform_R[456][9] = r_cell_wire[401];							inform_R[201][9] = r_cell_wire[402];							inform_R[457][9] = r_cell_wire[403];							inform_R[202][9] = r_cell_wire[404];							inform_R[458][9] = r_cell_wire[405];							inform_R[203][9] = r_cell_wire[406];							inform_R[459][9] = r_cell_wire[407];							inform_R[204][9] = r_cell_wire[408];							inform_R[460][9] = r_cell_wire[409];							inform_R[205][9] = r_cell_wire[410];							inform_R[461][9] = r_cell_wire[411];							inform_R[206][9] = r_cell_wire[412];							inform_R[462][9] = r_cell_wire[413];							inform_R[207][9] = r_cell_wire[414];							inform_R[463][9] = r_cell_wire[415];							inform_R[208][9] = r_cell_wire[416];							inform_R[464][9] = r_cell_wire[417];							inform_R[209][9] = r_cell_wire[418];							inform_R[465][9] = r_cell_wire[419];							inform_R[210][9] = r_cell_wire[420];							inform_R[466][9] = r_cell_wire[421];							inform_R[211][9] = r_cell_wire[422];							inform_R[467][9] = r_cell_wire[423];							inform_R[212][9] = r_cell_wire[424];							inform_R[468][9] = r_cell_wire[425];							inform_R[213][9] = r_cell_wire[426];							inform_R[469][9] = r_cell_wire[427];							inform_R[214][9] = r_cell_wire[428];							inform_R[470][9] = r_cell_wire[429];							inform_R[215][9] = r_cell_wire[430];							inform_R[471][9] = r_cell_wire[431];							inform_R[216][9] = r_cell_wire[432];							inform_R[472][9] = r_cell_wire[433];							inform_R[217][9] = r_cell_wire[434];							inform_R[473][9] = r_cell_wire[435];							inform_R[218][9] = r_cell_wire[436];							inform_R[474][9] = r_cell_wire[437];							inform_R[219][9] = r_cell_wire[438];							inform_R[475][9] = r_cell_wire[439];							inform_R[220][9] = r_cell_wire[440];							inform_R[476][9] = r_cell_wire[441];							inform_R[221][9] = r_cell_wire[442];							inform_R[477][9] = r_cell_wire[443];							inform_R[222][9] = r_cell_wire[444];							inform_R[478][9] = r_cell_wire[445];							inform_R[223][9] = r_cell_wire[446];							inform_R[479][9] = r_cell_wire[447];							inform_R[224][9] = r_cell_wire[448];							inform_R[480][9] = r_cell_wire[449];							inform_R[225][9] = r_cell_wire[450];							inform_R[481][9] = r_cell_wire[451];							inform_R[226][9] = r_cell_wire[452];							inform_R[482][9] = r_cell_wire[453];							inform_R[227][9] = r_cell_wire[454];							inform_R[483][9] = r_cell_wire[455];							inform_R[228][9] = r_cell_wire[456];							inform_R[484][9] = r_cell_wire[457];							inform_R[229][9] = r_cell_wire[458];							inform_R[485][9] = r_cell_wire[459];							inform_R[230][9] = r_cell_wire[460];							inform_R[486][9] = r_cell_wire[461];							inform_R[231][9] = r_cell_wire[462];							inform_R[487][9] = r_cell_wire[463];							inform_R[232][9] = r_cell_wire[464];							inform_R[488][9] = r_cell_wire[465];							inform_R[233][9] = r_cell_wire[466];							inform_R[489][9] = r_cell_wire[467];							inform_R[234][9] = r_cell_wire[468];							inform_R[490][9] = r_cell_wire[469];							inform_R[235][9] = r_cell_wire[470];							inform_R[491][9] = r_cell_wire[471];							inform_R[236][9] = r_cell_wire[472];							inform_R[492][9] = r_cell_wire[473];							inform_R[237][9] = r_cell_wire[474];							inform_R[493][9] = r_cell_wire[475];							inform_R[238][9] = r_cell_wire[476];							inform_R[494][9] = r_cell_wire[477];							inform_R[239][9] = r_cell_wire[478];							inform_R[495][9] = r_cell_wire[479];							inform_R[240][9] = r_cell_wire[480];							inform_R[496][9] = r_cell_wire[481];							inform_R[241][9] = r_cell_wire[482];							inform_R[497][9] = r_cell_wire[483];							inform_R[242][9] = r_cell_wire[484];							inform_R[498][9] = r_cell_wire[485];							inform_R[243][9] = r_cell_wire[486];							inform_R[499][9] = r_cell_wire[487];							inform_R[244][9] = r_cell_wire[488];							inform_R[500][9] = r_cell_wire[489];							inform_R[245][9] = r_cell_wire[490];							inform_R[501][9] = r_cell_wire[491];							inform_R[246][9] = r_cell_wire[492];							inform_R[502][9] = r_cell_wire[493];							inform_R[247][9] = r_cell_wire[494];							inform_R[503][9] = r_cell_wire[495];							inform_R[248][9] = r_cell_wire[496];							inform_R[504][9] = r_cell_wire[497];							inform_R[249][9] = r_cell_wire[498];							inform_R[505][9] = r_cell_wire[499];							inform_R[250][9] = r_cell_wire[500];							inform_R[506][9] = r_cell_wire[501];							inform_R[251][9] = r_cell_wire[502];							inform_R[507][9] = r_cell_wire[503];							inform_R[252][9] = r_cell_wire[504];							inform_R[508][9] = r_cell_wire[505];							inform_R[253][9] = r_cell_wire[506];							inform_R[509][9] = r_cell_wire[507];							inform_R[254][9] = r_cell_wire[508];							inform_R[510][9] = r_cell_wire[509];							inform_R[255][9] = r_cell_wire[510];							inform_R[511][9] = r_cell_wire[511];							inform_R[512][9] = r_cell_wire[512];							inform_R[768][9] = r_cell_wire[513];							inform_R[513][9] = r_cell_wire[514];							inform_R[769][9] = r_cell_wire[515];							inform_R[514][9] = r_cell_wire[516];							inform_R[770][9] = r_cell_wire[517];							inform_R[515][9] = r_cell_wire[518];							inform_R[771][9] = r_cell_wire[519];							inform_R[516][9] = r_cell_wire[520];							inform_R[772][9] = r_cell_wire[521];							inform_R[517][9] = r_cell_wire[522];							inform_R[773][9] = r_cell_wire[523];							inform_R[518][9] = r_cell_wire[524];							inform_R[774][9] = r_cell_wire[525];							inform_R[519][9] = r_cell_wire[526];							inform_R[775][9] = r_cell_wire[527];							inform_R[520][9] = r_cell_wire[528];							inform_R[776][9] = r_cell_wire[529];							inform_R[521][9] = r_cell_wire[530];							inform_R[777][9] = r_cell_wire[531];							inform_R[522][9] = r_cell_wire[532];							inform_R[778][9] = r_cell_wire[533];							inform_R[523][9] = r_cell_wire[534];							inform_R[779][9] = r_cell_wire[535];							inform_R[524][9] = r_cell_wire[536];							inform_R[780][9] = r_cell_wire[537];							inform_R[525][9] = r_cell_wire[538];							inform_R[781][9] = r_cell_wire[539];							inform_R[526][9] = r_cell_wire[540];							inform_R[782][9] = r_cell_wire[541];							inform_R[527][9] = r_cell_wire[542];							inform_R[783][9] = r_cell_wire[543];							inform_R[528][9] = r_cell_wire[544];							inform_R[784][9] = r_cell_wire[545];							inform_R[529][9] = r_cell_wire[546];							inform_R[785][9] = r_cell_wire[547];							inform_R[530][9] = r_cell_wire[548];							inform_R[786][9] = r_cell_wire[549];							inform_R[531][9] = r_cell_wire[550];							inform_R[787][9] = r_cell_wire[551];							inform_R[532][9] = r_cell_wire[552];							inform_R[788][9] = r_cell_wire[553];							inform_R[533][9] = r_cell_wire[554];							inform_R[789][9] = r_cell_wire[555];							inform_R[534][9] = r_cell_wire[556];							inform_R[790][9] = r_cell_wire[557];							inform_R[535][9] = r_cell_wire[558];							inform_R[791][9] = r_cell_wire[559];							inform_R[536][9] = r_cell_wire[560];							inform_R[792][9] = r_cell_wire[561];							inform_R[537][9] = r_cell_wire[562];							inform_R[793][9] = r_cell_wire[563];							inform_R[538][9] = r_cell_wire[564];							inform_R[794][9] = r_cell_wire[565];							inform_R[539][9] = r_cell_wire[566];							inform_R[795][9] = r_cell_wire[567];							inform_R[540][9] = r_cell_wire[568];							inform_R[796][9] = r_cell_wire[569];							inform_R[541][9] = r_cell_wire[570];							inform_R[797][9] = r_cell_wire[571];							inform_R[542][9] = r_cell_wire[572];							inform_R[798][9] = r_cell_wire[573];							inform_R[543][9] = r_cell_wire[574];							inform_R[799][9] = r_cell_wire[575];							inform_R[544][9] = r_cell_wire[576];							inform_R[800][9] = r_cell_wire[577];							inform_R[545][9] = r_cell_wire[578];							inform_R[801][9] = r_cell_wire[579];							inform_R[546][9] = r_cell_wire[580];							inform_R[802][9] = r_cell_wire[581];							inform_R[547][9] = r_cell_wire[582];							inform_R[803][9] = r_cell_wire[583];							inform_R[548][9] = r_cell_wire[584];							inform_R[804][9] = r_cell_wire[585];							inform_R[549][9] = r_cell_wire[586];							inform_R[805][9] = r_cell_wire[587];							inform_R[550][9] = r_cell_wire[588];							inform_R[806][9] = r_cell_wire[589];							inform_R[551][9] = r_cell_wire[590];							inform_R[807][9] = r_cell_wire[591];							inform_R[552][9] = r_cell_wire[592];							inform_R[808][9] = r_cell_wire[593];							inform_R[553][9] = r_cell_wire[594];							inform_R[809][9] = r_cell_wire[595];							inform_R[554][9] = r_cell_wire[596];							inform_R[810][9] = r_cell_wire[597];							inform_R[555][9] = r_cell_wire[598];							inform_R[811][9] = r_cell_wire[599];							inform_R[556][9] = r_cell_wire[600];							inform_R[812][9] = r_cell_wire[601];							inform_R[557][9] = r_cell_wire[602];							inform_R[813][9] = r_cell_wire[603];							inform_R[558][9] = r_cell_wire[604];							inform_R[814][9] = r_cell_wire[605];							inform_R[559][9] = r_cell_wire[606];							inform_R[815][9] = r_cell_wire[607];							inform_R[560][9] = r_cell_wire[608];							inform_R[816][9] = r_cell_wire[609];							inform_R[561][9] = r_cell_wire[610];							inform_R[817][9] = r_cell_wire[611];							inform_R[562][9] = r_cell_wire[612];							inform_R[818][9] = r_cell_wire[613];							inform_R[563][9] = r_cell_wire[614];							inform_R[819][9] = r_cell_wire[615];							inform_R[564][9] = r_cell_wire[616];							inform_R[820][9] = r_cell_wire[617];							inform_R[565][9] = r_cell_wire[618];							inform_R[821][9] = r_cell_wire[619];							inform_R[566][9] = r_cell_wire[620];							inform_R[822][9] = r_cell_wire[621];							inform_R[567][9] = r_cell_wire[622];							inform_R[823][9] = r_cell_wire[623];							inform_R[568][9] = r_cell_wire[624];							inform_R[824][9] = r_cell_wire[625];							inform_R[569][9] = r_cell_wire[626];							inform_R[825][9] = r_cell_wire[627];							inform_R[570][9] = r_cell_wire[628];							inform_R[826][9] = r_cell_wire[629];							inform_R[571][9] = r_cell_wire[630];							inform_R[827][9] = r_cell_wire[631];							inform_R[572][9] = r_cell_wire[632];							inform_R[828][9] = r_cell_wire[633];							inform_R[573][9] = r_cell_wire[634];							inform_R[829][9] = r_cell_wire[635];							inform_R[574][9] = r_cell_wire[636];							inform_R[830][9] = r_cell_wire[637];							inform_R[575][9] = r_cell_wire[638];							inform_R[831][9] = r_cell_wire[639];							inform_R[576][9] = r_cell_wire[640];							inform_R[832][9] = r_cell_wire[641];							inform_R[577][9] = r_cell_wire[642];							inform_R[833][9] = r_cell_wire[643];							inform_R[578][9] = r_cell_wire[644];							inform_R[834][9] = r_cell_wire[645];							inform_R[579][9] = r_cell_wire[646];							inform_R[835][9] = r_cell_wire[647];							inform_R[580][9] = r_cell_wire[648];							inform_R[836][9] = r_cell_wire[649];							inform_R[581][9] = r_cell_wire[650];							inform_R[837][9] = r_cell_wire[651];							inform_R[582][9] = r_cell_wire[652];							inform_R[838][9] = r_cell_wire[653];							inform_R[583][9] = r_cell_wire[654];							inform_R[839][9] = r_cell_wire[655];							inform_R[584][9] = r_cell_wire[656];							inform_R[840][9] = r_cell_wire[657];							inform_R[585][9] = r_cell_wire[658];							inform_R[841][9] = r_cell_wire[659];							inform_R[586][9] = r_cell_wire[660];							inform_R[842][9] = r_cell_wire[661];							inform_R[587][9] = r_cell_wire[662];							inform_R[843][9] = r_cell_wire[663];							inform_R[588][9] = r_cell_wire[664];							inform_R[844][9] = r_cell_wire[665];							inform_R[589][9] = r_cell_wire[666];							inform_R[845][9] = r_cell_wire[667];							inform_R[590][9] = r_cell_wire[668];							inform_R[846][9] = r_cell_wire[669];							inform_R[591][9] = r_cell_wire[670];							inform_R[847][9] = r_cell_wire[671];							inform_R[592][9] = r_cell_wire[672];							inform_R[848][9] = r_cell_wire[673];							inform_R[593][9] = r_cell_wire[674];							inform_R[849][9] = r_cell_wire[675];							inform_R[594][9] = r_cell_wire[676];							inform_R[850][9] = r_cell_wire[677];							inform_R[595][9] = r_cell_wire[678];							inform_R[851][9] = r_cell_wire[679];							inform_R[596][9] = r_cell_wire[680];							inform_R[852][9] = r_cell_wire[681];							inform_R[597][9] = r_cell_wire[682];							inform_R[853][9] = r_cell_wire[683];							inform_R[598][9] = r_cell_wire[684];							inform_R[854][9] = r_cell_wire[685];							inform_R[599][9] = r_cell_wire[686];							inform_R[855][9] = r_cell_wire[687];							inform_R[600][9] = r_cell_wire[688];							inform_R[856][9] = r_cell_wire[689];							inform_R[601][9] = r_cell_wire[690];							inform_R[857][9] = r_cell_wire[691];							inform_R[602][9] = r_cell_wire[692];							inform_R[858][9] = r_cell_wire[693];							inform_R[603][9] = r_cell_wire[694];							inform_R[859][9] = r_cell_wire[695];							inform_R[604][9] = r_cell_wire[696];							inform_R[860][9] = r_cell_wire[697];							inform_R[605][9] = r_cell_wire[698];							inform_R[861][9] = r_cell_wire[699];							inform_R[606][9] = r_cell_wire[700];							inform_R[862][9] = r_cell_wire[701];							inform_R[607][9] = r_cell_wire[702];							inform_R[863][9] = r_cell_wire[703];							inform_R[608][9] = r_cell_wire[704];							inform_R[864][9] = r_cell_wire[705];							inform_R[609][9] = r_cell_wire[706];							inform_R[865][9] = r_cell_wire[707];							inform_R[610][9] = r_cell_wire[708];							inform_R[866][9] = r_cell_wire[709];							inform_R[611][9] = r_cell_wire[710];							inform_R[867][9] = r_cell_wire[711];							inform_R[612][9] = r_cell_wire[712];							inform_R[868][9] = r_cell_wire[713];							inform_R[613][9] = r_cell_wire[714];							inform_R[869][9] = r_cell_wire[715];							inform_R[614][9] = r_cell_wire[716];							inform_R[870][9] = r_cell_wire[717];							inform_R[615][9] = r_cell_wire[718];							inform_R[871][9] = r_cell_wire[719];							inform_R[616][9] = r_cell_wire[720];							inform_R[872][9] = r_cell_wire[721];							inform_R[617][9] = r_cell_wire[722];							inform_R[873][9] = r_cell_wire[723];							inform_R[618][9] = r_cell_wire[724];							inform_R[874][9] = r_cell_wire[725];							inform_R[619][9] = r_cell_wire[726];							inform_R[875][9] = r_cell_wire[727];							inform_R[620][9] = r_cell_wire[728];							inform_R[876][9] = r_cell_wire[729];							inform_R[621][9] = r_cell_wire[730];							inform_R[877][9] = r_cell_wire[731];							inform_R[622][9] = r_cell_wire[732];							inform_R[878][9] = r_cell_wire[733];							inform_R[623][9] = r_cell_wire[734];							inform_R[879][9] = r_cell_wire[735];							inform_R[624][9] = r_cell_wire[736];							inform_R[880][9] = r_cell_wire[737];							inform_R[625][9] = r_cell_wire[738];							inform_R[881][9] = r_cell_wire[739];							inform_R[626][9] = r_cell_wire[740];							inform_R[882][9] = r_cell_wire[741];							inform_R[627][9] = r_cell_wire[742];							inform_R[883][9] = r_cell_wire[743];							inform_R[628][9] = r_cell_wire[744];							inform_R[884][9] = r_cell_wire[745];							inform_R[629][9] = r_cell_wire[746];							inform_R[885][9] = r_cell_wire[747];							inform_R[630][9] = r_cell_wire[748];							inform_R[886][9] = r_cell_wire[749];							inform_R[631][9] = r_cell_wire[750];							inform_R[887][9] = r_cell_wire[751];							inform_R[632][9] = r_cell_wire[752];							inform_R[888][9] = r_cell_wire[753];							inform_R[633][9] = r_cell_wire[754];							inform_R[889][9] = r_cell_wire[755];							inform_R[634][9] = r_cell_wire[756];							inform_R[890][9] = r_cell_wire[757];							inform_R[635][9] = r_cell_wire[758];							inform_R[891][9] = r_cell_wire[759];							inform_R[636][9] = r_cell_wire[760];							inform_R[892][9] = r_cell_wire[761];							inform_R[637][9] = r_cell_wire[762];							inform_R[893][9] = r_cell_wire[763];							inform_R[638][9] = r_cell_wire[764];							inform_R[894][9] = r_cell_wire[765];							inform_R[639][9] = r_cell_wire[766];							inform_R[895][9] = r_cell_wire[767];							inform_R[640][9] = r_cell_wire[768];							inform_R[896][9] = r_cell_wire[769];							inform_R[641][9] = r_cell_wire[770];							inform_R[897][9] = r_cell_wire[771];							inform_R[642][9] = r_cell_wire[772];							inform_R[898][9] = r_cell_wire[773];							inform_R[643][9] = r_cell_wire[774];							inform_R[899][9] = r_cell_wire[775];							inform_R[644][9] = r_cell_wire[776];							inform_R[900][9] = r_cell_wire[777];							inform_R[645][9] = r_cell_wire[778];							inform_R[901][9] = r_cell_wire[779];							inform_R[646][9] = r_cell_wire[780];							inform_R[902][9] = r_cell_wire[781];							inform_R[647][9] = r_cell_wire[782];							inform_R[903][9] = r_cell_wire[783];							inform_R[648][9] = r_cell_wire[784];							inform_R[904][9] = r_cell_wire[785];							inform_R[649][9] = r_cell_wire[786];							inform_R[905][9] = r_cell_wire[787];							inform_R[650][9] = r_cell_wire[788];							inform_R[906][9] = r_cell_wire[789];							inform_R[651][9] = r_cell_wire[790];							inform_R[907][9] = r_cell_wire[791];							inform_R[652][9] = r_cell_wire[792];							inform_R[908][9] = r_cell_wire[793];							inform_R[653][9] = r_cell_wire[794];							inform_R[909][9] = r_cell_wire[795];							inform_R[654][9] = r_cell_wire[796];							inform_R[910][9] = r_cell_wire[797];							inform_R[655][9] = r_cell_wire[798];							inform_R[911][9] = r_cell_wire[799];							inform_R[656][9] = r_cell_wire[800];							inform_R[912][9] = r_cell_wire[801];							inform_R[657][9] = r_cell_wire[802];							inform_R[913][9] = r_cell_wire[803];							inform_R[658][9] = r_cell_wire[804];							inform_R[914][9] = r_cell_wire[805];							inform_R[659][9] = r_cell_wire[806];							inform_R[915][9] = r_cell_wire[807];							inform_R[660][9] = r_cell_wire[808];							inform_R[916][9] = r_cell_wire[809];							inform_R[661][9] = r_cell_wire[810];							inform_R[917][9] = r_cell_wire[811];							inform_R[662][9] = r_cell_wire[812];							inform_R[918][9] = r_cell_wire[813];							inform_R[663][9] = r_cell_wire[814];							inform_R[919][9] = r_cell_wire[815];							inform_R[664][9] = r_cell_wire[816];							inform_R[920][9] = r_cell_wire[817];							inform_R[665][9] = r_cell_wire[818];							inform_R[921][9] = r_cell_wire[819];							inform_R[666][9] = r_cell_wire[820];							inform_R[922][9] = r_cell_wire[821];							inform_R[667][9] = r_cell_wire[822];							inform_R[923][9] = r_cell_wire[823];							inform_R[668][9] = r_cell_wire[824];							inform_R[924][9] = r_cell_wire[825];							inform_R[669][9] = r_cell_wire[826];							inform_R[925][9] = r_cell_wire[827];							inform_R[670][9] = r_cell_wire[828];							inform_R[926][9] = r_cell_wire[829];							inform_R[671][9] = r_cell_wire[830];							inform_R[927][9] = r_cell_wire[831];							inform_R[672][9] = r_cell_wire[832];							inform_R[928][9] = r_cell_wire[833];							inform_R[673][9] = r_cell_wire[834];							inform_R[929][9] = r_cell_wire[835];							inform_R[674][9] = r_cell_wire[836];							inform_R[930][9] = r_cell_wire[837];							inform_R[675][9] = r_cell_wire[838];							inform_R[931][9] = r_cell_wire[839];							inform_R[676][9] = r_cell_wire[840];							inform_R[932][9] = r_cell_wire[841];							inform_R[677][9] = r_cell_wire[842];							inform_R[933][9] = r_cell_wire[843];							inform_R[678][9] = r_cell_wire[844];							inform_R[934][9] = r_cell_wire[845];							inform_R[679][9] = r_cell_wire[846];							inform_R[935][9] = r_cell_wire[847];							inform_R[680][9] = r_cell_wire[848];							inform_R[936][9] = r_cell_wire[849];							inform_R[681][9] = r_cell_wire[850];							inform_R[937][9] = r_cell_wire[851];							inform_R[682][9] = r_cell_wire[852];							inform_R[938][9] = r_cell_wire[853];							inform_R[683][9] = r_cell_wire[854];							inform_R[939][9] = r_cell_wire[855];							inform_R[684][9] = r_cell_wire[856];							inform_R[940][9] = r_cell_wire[857];							inform_R[685][9] = r_cell_wire[858];							inform_R[941][9] = r_cell_wire[859];							inform_R[686][9] = r_cell_wire[860];							inform_R[942][9] = r_cell_wire[861];							inform_R[687][9] = r_cell_wire[862];							inform_R[943][9] = r_cell_wire[863];							inform_R[688][9] = r_cell_wire[864];							inform_R[944][9] = r_cell_wire[865];							inform_R[689][9] = r_cell_wire[866];							inform_R[945][9] = r_cell_wire[867];							inform_R[690][9] = r_cell_wire[868];							inform_R[946][9] = r_cell_wire[869];							inform_R[691][9] = r_cell_wire[870];							inform_R[947][9] = r_cell_wire[871];							inform_R[692][9] = r_cell_wire[872];							inform_R[948][9] = r_cell_wire[873];							inform_R[693][9] = r_cell_wire[874];							inform_R[949][9] = r_cell_wire[875];							inform_R[694][9] = r_cell_wire[876];							inform_R[950][9] = r_cell_wire[877];							inform_R[695][9] = r_cell_wire[878];							inform_R[951][9] = r_cell_wire[879];							inform_R[696][9] = r_cell_wire[880];							inform_R[952][9] = r_cell_wire[881];							inform_R[697][9] = r_cell_wire[882];							inform_R[953][9] = r_cell_wire[883];							inform_R[698][9] = r_cell_wire[884];							inform_R[954][9] = r_cell_wire[885];							inform_R[699][9] = r_cell_wire[886];							inform_R[955][9] = r_cell_wire[887];							inform_R[700][9] = r_cell_wire[888];							inform_R[956][9] = r_cell_wire[889];							inform_R[701][9] = r_cell_wire[890];							inform_R[957][9] = r_cell_wire[891];							inform_R[702][9] = r_cell_wire[892];							inform_R[958][9] = r_cell_wire[893];							inform_R[703][9] = r_cell_wire[894];							inform_R[959][9] = r_cell_wire[895];							inform_R[704][9] = r_cell_wire[896];							inform_R[960][9] = r_cell_wire[897];							inform_R[705][9] = r_cell_wire[898];							inform_R[961][9] = r_cell_wire[899];							inform_R[706][9] = r_cell_wire[900];							inform_R[962][9] = r_cell_wire[901];							inform_R[707][9] = r_cell_wire[902];							inform_R[963][9] = r_cell_wire[903];							inform_R[708][9] = r_cell_wire[904];							inform_R[964][9] = r_cell_wire[905];							inform_R[709][9] = r_cell_wire[906];							inform_R[965][9] = r_cell_wire[907];							inform_R[710][9] = r_cell_wire[908];							inform_R[966][9] = r_cell_wire[909];							inform_R[711][9] = r_cell_wire[910];							inform_R[967][9] = r_cell_wire[911];							inform_R[712][9] = r_cell_wire[912];							inform_R[968][9] = r_cell_wire[913];							inform_R[713][9] = r_cell_wire[914];							inform_R[969][9] = r_cell_wire[915];							inform_R[714][9] = r_cell_wire[916];							inform_R[970][9] = r_cell_wire[917];							inform_R[715][9] = r_cell_wire[918];							inform_R[971][9] = r_cell_wire[919];							inform_R[716][9] = r_cell_wire[920];							inform_R[972][9] = r_cell_wire[921];							inform_R[717][9] = r_cell_wire[922];							inform_R[973][9] = r_cell_wire[923];							inform_R[718][9] = r_cell_wire[924];							inform_R[974][9] = r_cell_wire[925];							inform_R[719][9] = r_cell_wire[926];							inform_R[975][9] = r_cell_wire[927];							inform_R[720][9] = r_cell_wire[928];							inform_R[976][9] = r_cell_wire[929];							inform_R[721][9] = r_cell_wire[930];							inform_R[977][9] = r_cell_wire[931];							inform_R[722][9] = r_cell_wire[932];							inform_R[978][9] = r_cell_wire[933];							inform_R[723][9] = r_cell_wire[934];							inform_R[979][9] = r_cell_wire[935];							inform_R[724][9] = r_cell_wire[936];							inform_R[980][9] = r_cell_wire[937];							inform_R[725][9] = r_cell_wire[938];							inform_R[981][9] = r_cell_wire[939];							inform_R[726][9] = r_cell_wire[940];							inform_R[982][9] = r_cell_wire[941];							inform_R[727][9] = r_cell_wire[942];							inform_R[983][9] = r_cell_wire[943];							inform_R[728][9] = r_cell_wire[944];							inform_R[984][9] = r_cell_wire[945];							inform_R[729][9] = r_cell_wire[946];							inform_R[985][9] = r_cell_wire[947];							inform_R[730][9] = r_cell_wire[948];							inform_R[986][9] = r_cell_wire[949];							inform_R[731][9] = r_cell_wire[950];							inform_R[987][9] = r_cell_wire[951];							inform_R[732][9] = r_cell_wire[952];							inform_R[988][9] = r_cell_wire[953];							inform_R[733][9] = r_cell_wire[954];							inform_R[989][9] = r_cell_wire[955];							inform_R[734][9] = r_cell_wire[956];							inform_R[990][9] = r_cell_wire[957];							inform_R[735][9] = r_cell_wire[958];							inform_R[991][9] = r_cell_wire[959];							inform_R[736][9] = r_cell_wire[960];							inform_R[992][9] = r_cell_wire[961];							inform_R[737][9] = r_cell_wire[962];							inform_R[993][9] = r_cell_wire[963];							inform_R[738][9] = r_cell_wire[964];							inform_R[994][9] = r_cell_wire[965];							inform_R[739][9] = r_cell_wire[966];							inform_R[995][9] = r_cell_wire[967];							inform_R[740][9] = r_cell_wire[968];							inform_R[996][9] = r_cell_wire[969];							inform_R[741][9] = r_cell_wire[970];							inform_R[997][9] = r_cell_wire[971];							inform_R[742][9] = r_cell_wire[972];							inform_R[998][9] = r_cell_wire[973];							inform_R[743][9] = r_cell_wire[974];							inform_R[999][9] = r_cell_wire[975];							inform_R[744][9] = r_cell_wire[976];							inform_R[1000][9] = r_cell_wire[977];							inform_R[745][9] = r_cell_wire[978];							inform_R[1001][9] = r_cell_wire[979];							inform_R[746][9] = r_cell_wire[980];							inform_R[1002][9] = r_cell_wire[981];							inform_R[747][9] = r_cell_wire[982];							inform_R[1003][9] = r_cell_wire[983];							inform_R[748][9] = r_cell_wire[984];							inform_R[1004][9] = r_cell_wire[985];							inform_R[749][9] = r_cell_wire[986];							inform_R[1005][9] = r_cell_wire[987];							inform_R[750][9] = r_cell_wire[988];							inform_R[1006][9] = r_cell_wire[989];							inform_R[751][9] = r_cell_wire[990];							inform_R[1007][9] = r_cell_wire[991];							inform_R[752][9] = r_cell_wire[992];							inform_R[1008][9] = r_cell_wire[993];							inform_R[753][9] = r_cell_wire[994];							inform_R[1009][9] = r_cell_wire[995];							inform_R[754][9] = r_cell_wire[996];							inform_R[1010][9] = r_cell_wire[997];							inform_R[755][9] = r_cell_wire[998];							inform_R[1011][9] = r_cell_wire[999];							inform_R[756][9] = r_cell_wire[1000];							inform_R[1012][9] = r_cell_wire[1001];							inform_R[757][9] = r_cell_wire[1002];							inform_R[1013][9] = r_cell_wire[1003];							inform_R[758][9] = r_cell_wire[1004];							inform_R[1014][9] = r_cell_wire[1005];							inform_R[759][9] = r_cell_wire[1006];							inform_R[1015][9] = r_cell_wire[1007];							inform_R[760][9] = r_cell_wire[1008];							inform_R[1016][9] = r_cell_wire[1009];							inform_R[761][9] = r_cell_wire[1010];							inform_R[1017][9] = r_cell_wire[1011];							inform_R[762][9] = r_cell_wire[1012];							inform_R[1018][9] = r_cell_wire[1013];							inform_R[763][9] = r_cell_wire[1014];							inform_R[1019][9] = r_cell_wire[1015];							inform_R[764][9] = r_cell_wire[1016];							inform_R[1020][9] = r_cell_wire[1017];							inform_R[765][9] = r_cell_wire[1018];							inform_R[1021][9] = r_cell_wire[1019];							inform_R[766][9] = r_cell_wire[1020];							inform_R[1022][9] = r_cell_wire[1021];							inform_R[767][9] = r_cell_wire[1022];							inform_R[1023][9] = r_cell_wire[1023];							inform_L[0][8] = l_cell_wire[0];							inform_L[256][8] = l_cell_wire[1];							inform_L[1][8] = l_cell_wire[2];							inform_L[257][8] = l_cell_wire[3];							inform_L[2][8] = l_cell_wire[4];							inform_L[258][8] = l_cell_wire[5];							inform_L[3][8] = l_cell_wire[6];							inform_L[259][8] = l_cell_wire[7];							inform_L[4][8] = l_cell_wire[8];							inform_L[260][8] = l_cell_wire[9];							inform_L[5][8] = l_cell_wire[10];							inform_L[261][8] = l_cell_wire[11];							inform_L[6][8] = l_cell_wire[12];							inform_L[262][8] = l_cell_wire[13];							inform_L[7][8] = l_cell_wire[14];							inform_L[263][8] = l_cell_wire[15];							inform_L[8][8] = l_cell_wire[16];							inform_L[264][8] = l_cell_wire[17];							inform_L[9][8] = l_cell_wire[18];							inform_L[265][8] = l_cell_wire[19];							inform_L[10][8] = l_cell_wire[20];							inform_L[266][8] = l_cell_wire[21];							inform_L[11][8] = l_cell_wire[22];							inform_L[267][8] = l_cell_wire[23];							inform_L[12][8] = l_cell_wire[24];							inform_L[268][8] = l_cell_wire[25];							inform_L[13][8] = l_cell_wire[26];							inform_L[269][8] = l_cell_wire[27];							inform_L[14][8] = l_cell_wire[28];							inform_L[270][8] = l_cell_wire[29];							inform_L[15][8] = l_cell_wire[30];							inform_L[271][8] = l_cell_wire[31];							inform_L[16][8] = l_cell_wire[32];							inform_L[272][8] = l_cell_wire[33];							inform_L[17][8] = l_cell_wire[34];							inform_L[273][8] = l_cell_wire[35];							inform_L[18][8] = l_cell_wire[36];							inform_L[274][8] = l_cell_wire[37];							inform_L[19][8] = l_cell_wire[38];							inform_L[275][8] = l_cell_wire[39];							inform_L[20][8] = l_cell_wire[40];							inform_L[276][8] = l_cell_wire[41];							inform_L[21][8] = l_cell_wire[42];							inform_L[277][8] = l_cell_wire[43];							inform_L[22][8] = l_cell_wire[44];							inform_L[278][8] = l_cell_wire[45];							inform_L[23][8] = l_cell_wire[46];							inform_L[279][8] = l_cell_wire[47];							inform_L[24][8] = l_cell_wire[48];							inform_L[280][8] = l_cell_wire[49];							inform_L[25][8] = l_cell_wire[50];							inform_L[281][8] = l_cell_wire[51];							inform_L[26][8] = l_cell_wire[52];							inform_L[282][8] = l_cell_wire[53];							inform_L[27][8] = l_cell_wire[54];							inform_L[283][8] = l_cell_wire[55];							inform_L[28][8] = l_cell_wire[56];							inform_L[284][8] = l_cell_wire[57];							inform_L[29][8] = l_cell_wire[58];							inform_L[285][8] = l_cell_wire[59];							inform_L[30][8] = l_cell_wire[60];							inform_L[286][8] = l_cell_wire[61];							inform_L[31][8] = l_cell_wire[62];							inform_L[287][8] = l_cell_wire[63];							inform_L[32][8] = l_cell_wire[64];							inform_L[288][8] = l_cell_wire[65];							inform_L[33][8] = l_cell_wire[66];							inform_L[289][8] = l_cell_wire[67];							inform_L[34][8] = l_cell_wire[68];							inform_L[290][8] = l_cell_wire[69];							inform_L[35][8] = l_cell_wire[70];							inform_L[291][8] = l_cell_wire[71];							inform_L[36][8] = l_cell_wire[72];							inform_L[292][8] = l_cell_wire[73];							inform_L[37][8] = l_cell_wire[74];							inform_L[293][8] = l_cell_wire[75];							inform_L[38][8] = l_cell_wire[76];							inform_L[294][8] = l_cell_wire[77];							inform_L[39][8] = l_cell_wire[78];							inform_L[295][8] = l_cell_wire[79];							inform_L[40][8] = l_cell_wire[80];							inform_L[296][8] = l_cell_wire[81];							inform_L[41][8] = l_cell_wire[82];							inform_L[297][8] = l_cell_wire[83];							inform_L[42][8] = l_cell_wire[84];							inform_L[298][8] = l_cell_wire[85];							inform_L[43][8] = l_cell_wire[86];							inform_L[299][8] = l_cell_wire[87];							inform_L[44][8] = l_cell_wire[88];							inform_L[300][8] = l_cell_wire[89];							inform_L[45][8] = l_cell_wire[90];							inform_L[301][8] = l_cell_wire[91];							inform_L[46][8] = l_cell_wire[92];							inform_L[302][8] = l_cell_wire[93];							inform_L[47][8] = l_cell_wire[94];							inform_L[303][8] = l_cell_wire[95];							inform_L[48][8] = l_cell_wire[96];							inform_L[304][8] = l_cell_wire[97];							inform_L[49][8] = l_cell_wire[98];							inform_L[305][8] = l_cell_wire[99];							inform_L[50][8] = l_cell_wire[100];							inform_L[306][8] = l_cell_wire[101];							inform_L[51][8] = l_cell_wire[102];							inform_L[307][8] = l_cell_wire[103];							inform_L[52][8] = l_cell_wire[104];							inform_L[308][8] = l_cell_wire[105];							inform_L[53][8] = l_cell_wire[106];							inform_L[309][8] = l_cell_wire[107];							inform_L[54][8] = l_cell_wire[108];							inform_L[310][8] = l_cell_wire[109];							inform_L[55][8] = l_cell_wire[110];							inform_L[311][8] = l_cell_wire[111];							inform_L[56][8] = l_cell_wire[112];							inform_L[312][8] = l_cell_wire[113];							inform_L[57][8] = l_cell_wire[114];							inform_L[313][8] = l_cell_wire[115];							inform_L[58][8] = l_cell_wire[116];							inform_L[314][8] = l_cell_wire[117];							inform_L[59][8] = l_cell_wire[118];							inform_L[315][8] = l_cell_wire[119];							inform_L[60][8] = l_cell_wire[120];							inform_L[316][8] = l_cell_wire[121];							inform_L[61][8] = l_cell_wire[122];							inform_L[317][8] = l_cell_wire[123];							inform_L[62][8] = l_cell_wire[124];							inform_L[318][8] = l_cell_wire[125];							inform_L[63][8] = l_cell_wire[126];							inform_L[319][8] = l_cell_wire[127];							inform_L[64][8] = l_cell_wire[128];							inform_L[320][8] = l_cell_wire[129];							inform_L[65][8] = l_cell_wire[130];							inform_L[321][8] = l_cell_wire[131];							inform_L[66][8] = l_cell_wire[132];							inform_L[322][8] = l_cell_wire[133];							inform_L[67][8] = l_cell_wire[134];							inform_L[323][8] = l_cell_wire[135];							inform_L[68][8] = l_cell_wire[136];							inform_L[324][8] = l_cell_wire[137];							inform_L[69][8] = l_cell_wire[138];							inform_L[325][8] = l_cell_wire[139];							inform_L[70][8] = l_cell_wire[140];							inform_L[326][8] = l_cell_wire[141];							inform_L[71][8] = l_cell_wire[142];							inform_L[327][8] = l_cell_wire[143];							inform_L[72][8] = l_cell_wire[144];							inform_L[328][8] = l_cell_wire[145];							inform_L[73][8] = l_cell_wire[146];							inform_L[329][8] = l_cell_wire[147];							inform_L[74][8] = l_cell_wire[148];							inform_L[330][8] = l_cell_wire[149];							inform_L[75][8] = l_cell_wire[150];							inform_L[331][8] = l_cell_wire[151];							inform_L[76][8] = l_cell_wire[152];							inform_L[332][8] = l_cell_wire[153];							inform_L[77][8] = l_cell_wire[154];							inform_L[333][8] = l_cell_wire[155];							inform_L[78][8] = l_cell_wire[156];							inform_L[334][8] = l_cell_wire[157];							inform_L[79][8] = l_cell_wire[158];							inform_L[335][8] = l_cell_wire[159];							inform_L[80][8] = l_cell_wire[160];							inform_L[336][8] = l_cell_wire[161];							inform_L[81][8] = l_cell_wire[162];							inform_L[337][8] = l_cell_wire[163];							inform_L[82][8] = l_cell_wire[164];							inform_L[338][8] = l_cell_wire[165];							inform_L[83][8] = l_cell_wire[166];							inform_L[339][8] = l_cell_wire[167];							inform_L[84][8] = l_cell_wire[168];							inform_L[340][8] = l_cell_wire[169];							inform_L[85][8] = l_cell_wire[170];							inform_L[341][8] = l_cell_wire[171];							inform_L[86][8] = l_cell_wire[172];							inform_L[342][8] = l_cell_wire[173];							inform_L[87][8] = l_cell_wire[174];							inform_L[343][8] = l_cell_wire[175];							inform_L[88][8] = l_cell_wire[176];							inform_L[344][8] = l_cell_wire[177];							inform_L[89][8] = l_cell_wire[178];							inform_L[345][8] = l_cell_wire[179];							inform_L[90][8] = l_cell_wire[180];							inform_L[346][8] = l_cell_wire[181];							inform_L[91][8] = l_cell_wire[182];							inform_L[347][8] = l_cell_wire[183];							inform_L[92][8] = l_cell_wire[184];							inform_L[348][8] = l_cell_wire[185];							inform_L[93][8] = l_cell_wire[186];							inform_L[349][8] = l_cell_wire[187];							inform_L[94][8] = l_cell_wire[188];							inform_L[350][8] = l_cell_wire[189];							inform_L[95][8] = l_cell_wire[190];							inform_L[351][8] = l_cell_wire[191];							inform_L[96][8] = l_cell_wire[192];							inform_L[352][8] = l_cell_wire[193];							inform_L[97][8] = l_cell_wire[194];							inform_L[353][8] = l_cell_wire[195];							inform_L[98][8] = l_cell_wire[196];							inform_L[354][8] = l_cell_wire[197];							inform_L[99][8] = l_cell_wire[198];							inform_L[355][8] = l_cell_wire[199];							inform_L[100][8] = l_cell_wire[200];							inform_L[356][8] = l_cell_wire[201];							inform_L[101][8] = l_cell_wire[202];							inform_L[357][8] = l_cell_wire[203];							inform_L[102][8] = l_cell_wire[204];							inform_L[358][8] = l_cell_wire[205];							inform_L[103][8] = l_cell_wire[206];							inform_L[359][8] = l_cell_wire[207];							inform_L[104][8] = l_cell_wire[208];							inform_L[360][8] = l_cell_wire[209];							inform_L[105][8] = l_cell_wire[210];							inform_L[361][8] = l_cell_wire[211];							inform_L[106][8] = l_cell_wire[212];							inform_L[362][8] = l_cell_wire[213];							inform_L[107][8] = l_cell_wire[214];							inform_L[363][8] = l_cell_wire[215];							inform_L[108][8] = l_cell_wire[216];							inform_L[364][8] = l_cell_wire[217];							inform_L[109][8] = l_cell_wire[218];							inform_L[365][8] = l_cell_wire[219];							inform_L[110][8] = l_cell_wire[220];							inform_L[366][8] = l_cell_wire[221];							inform_L[111][8] = l_cell_wire[222];							inform_L[367][8] = l_cell_wire[223];							inform_L[112][8] = l_cell_wire[224];							inform_L[368][8] = l_cell_wire[225];							inform_L[113][8] = l_cell_wire[226];							inform_L[369][8] = l_cell_wire[227];							inform_L[114][8] = l_cell_wire[228];							inform_L[370][8] = l_cell_wire[229];							inform_L[115][8] = l_cell_wire[230];							inform_L[371][8] = l_cell_wire[231];							inform_L[116][8] = l_cell_wire[232];							inform_L[372][8] = l_cell_wire[233];							inform_L[117][8] = l_cell_wire[234];							inform_L[373][8] = l_cell_wire[235];							inform_L[118][8] = l_cell_wire[236];							inform_L[374][8] = l_cell_wire[237];							inform_L[119][8] = l_cell_wire[238];							inform_L[375][8] = l_cell_wire[239];							inform_L[120][8] = l_cell_wire[240];							inform_L[376][8] = l_cell_wire[241];							inform_L[121][8] = l_cell_wire[242];							inform_L[377][8] = l_cell_wire[243];							inform_L[122][8] = l_cell_wire[244];							inform_L[378][8] = l_cell_wire[245];							inform_L[123][8] = l_cell_wire[246];							inform_L[379][8] = l_cell_wire[247];							inform_L[124][8] = l_cell_wire[248];							inform_L[380][8] = l_cell_wire[249];							inform_L[125][8] = l_cell_wire[250];							inform_L[381][8] = l_cell_wire[251];							inform_L[126][8] = l_cell_wire[252];							inform_L[382][8] = l_cell_wire[253];							inform_L[127][8] = l_cell_wire[254];							inform_L[383][8] = l_cell_wire[255];							inform_L[128][8] = l_cell_wire[256];							inform_L[384][8] = l_cell_wire[257];							inform_L[129][8] = l_cell_wire[258];							inform_L[385][8] = l_cell_wire[259];							inform_L[130][8] = l_cell_wire[260];							inform_L[386][8] = l_cell_wire[261];							inform_L[131][8] = l_cell_wire[262];							inform_L[387][8] = l_cell_wire[263];							inform_L[132][8] = l_cell_wire[264];							inform_L[388][8] = l_cell_wire[265];							inform_L[133][8] = l_cell_wire[266];							inform_L[389][8] = l_cell_wire[267];							inform_L[134][8] = l_cell_wire[268];							inform_L[390][8] = l_cell_wire[269];							inform_L[135][8] = l_cell_wire[270];							inform_L[391][8] = l_cell_wire[271];							inform_L[136][8] = l_cell_wire[272];							inform_L[392][8] = l_cell_wire[273];							inform_L[137][8] = l_cell_wire[274];							inform_L[393][8] = l_cell_wire[275];							inform_L[138][8] = l_cell_wire[276];							inform_L[394][8] = l_cell_wire[277];							inform_L[139][8] = l_cell_wire[278];							inform_L[395][8] = l_cell_wire[279];							inform_L[140][8] = l_cell_wire[280];							inform_L[396][8] = l_cell_wire[281];							inform_L[141][8] = l_cell_wire[282];							inform_L[397][8] = l_cell_wire[283];							inform_L[142][8] = l_cell_wire[284];							inform_L[398][8] = l_cell_wire[285];							inform_L[143][8] = l_cell_wire[286];							inform_L[399][8] = l_cell_wire[287];							inform_L[144][8] = l_cell_wire[288];							inform_L[400][8] = l_cell_wire[289];							inform_L[145][8] = l_cell_wire[290];							inform_L[401][8] = l_cell_wire[291];							inform_L[146][8] = l_cell_wire[292];							inform_L[402][8] = l_cell_wire[293];							inform_L[147][8] = l_cell_wire[294];							inform_L[403][8] = l_cell_wire[295];							inform_L[148][8] = l_cell_wire[296];							inform_L[404][8] = l_cell_wire[297];							inform_L[149][8] = l_cell_wire[298];							inform_L[405][8] = l_cell_wire[299];							inform_L[150][8] = l_cell_wire[300];							inform_L[406][8] = l_cell_wire[301];							inform_L[151][8] = l_cell_wire[302];							inform_L[407][8] = l_cell_wire[303];							inform_L[152][8] = l_cell_wire[304];							inform_L[408][8] = l_cell_wire[305];							inform_L[153][8] = l_cell_wire[306];							inform_L[409][8] = l_cell_wire[307];							inform_L[154][8] = l_cell_wire[308];							inform_L[410][8] = l_cell_wire[309];							inform_L[155][8] = l_cell_wire[310];							inform_L[411][8] = l_cell_wire[311];							inform_L[156][8] = l_cell_wire[312];							inform_L[412][8] = l_cell_wire[313];							inform_L[157][8] = l_cell_wire[314];							inform_L[413][8] = l_cell_wire[315];							inform_L[158][8] = l_cell_wire[316];							inform_L[414][8] = l_cell_wire[317];							inform_L[159][8] = l_cell_wire[318];							inform_L[415][8] = l_cell_wire[319];							inform_L[160][8] = l_cell_wire[320];							inform_L[416][8] = l_cell_wire[321];							inform_L[161][8] = l_cell_wire[322];							inform_L[417][8] = l_cell_wire[323];							inform_L[162][8] = l_cell_wire[324];							inform_L[418][8] = l_cell_wire[325];							inform_L[163][8] = l_cell_wire[326];							inform_L[419][8] = l_cell_wire[327];							inform_L[164][8] = l_cell_wire[328];							inform_L[420][8] = l_cell_wire[329];							inform_L[165][8] = l_cell_wire[330];							inform_L[421][8] = l_cell_wire[331];							inform_L[166][8] = l_cell_wire[332];							inform_L[422][8] = l_cell_wire[333];							inform_L[167][8] = l_cell_wire[334];							inform_L[423][8] = l_cell_wire[335];							inform_L[168][8] = l_cell_wire[336];							inform_L[424][8] = l_cell_wire[337];							inform_L[169][8] = l_cell_wire[338];							inform_L[425][8] = l_cell_wire[339];							inform_L[170][8] = l_cell_wire[340];							inform_L[426][8] = l_cell_wire[341];							inform_L[171][8] = l_cell_wire[342];							inform_L[427][8] = l_cell_wire[343];							inform_L[172][8] = l_cell_wire[344];							inform_L[428][8] = l_cell_wire[345];							inform_L[173][8] = l_cell_wire[346];							inform_L[429][8] = l_cell_wire[347];							inform_L[174][8] = l_cell_wire[348];							inform_L[430][8] = l_cell_wire[349];							inform_L[175][8] = l_cell_wire[350];							inform_L[431][8] = l_cell_wire[351];							inform_L[176][8] = l_cell_wire[352];							inform_L[432][8] = l_cell_wire[353];							inform_L[177][8] = l_cell_wire[354];							inform_L[433][8] = l_cell_wire[355];							inform_L[178][8] = l_cell_wire[356];							inform_L[434][8] = l_cell_wire[357];							inform_L[179][8] = l_cell_wire[358];							inform_L[435][8] = l_cell_wire[359];							inform_L[180][8] = l_cell_wire[360];							inform_L[436][8] = l_cell_wire[361];							inform_L[181][8] = l_cell_wire[362];							inform_L[437][8] = l_cell_wire[363];							inform_L[182][8] = l_cell_wire[364];							inform_L[438][8] = l_cell_wire[365];							inform_L[183][8] = l_cell_wire[366];							inform_L[439][8] = l_cell_wire[367];							inform_L[184][8] = l_cell_wire[368];							inform_L[440][8] = l_cell_wire[369];							inform_L[185][8] = l_cell_wire[370];							inform_L[441][8] = l_cell_wire[371];							inform_L[186][8] = l_cell_wire[372];							inform_L[442][8] = l_cell_wire[373];							inform_L[187][8] = l_cell_wire[374];							inform_L[443][8] = l_cell_wire[375];							inform_L[188][8] = l_cell_wire[376];							inform_L[444][8] = l_cell_wire[377];							inform_L[189][8] = l_cell_wire[378];							inform_L[445][8] = l_cell_wire[379];							inform_L[190][8] = l_cell_wire[380];							inform_L[446][8] = l_cell_wire[381];							inform_L[191][8] = l_cell_wire[382];							inform_L[447][8] = l_cell_wire[383];							inform_L[192][8] = l_cell_wire[384];							inform_L[448][8] = l_cell_wire[385];							inform_L[193][8] = l_cell_wire[386];							inform_L[449][8] = l_cell_wire[387];							inform_L[194][8] = l_cell_wire[388];							inform_L[450][8] = l_cell_wire[389];							inform_L[195][8] = l_cell_wire[390];							inform_L[451][8] = l_cell_wire[391];							inform_L[196][8] = l_cell_wire[392];							inform_L[452][8] = l_cell_wire[393];							inform_L[197][8] = l_cell_wire[394];							inform_L[453][8] = l_cell_wire[395];							inform_L[198][8] = l_cell_wire[396];							inform_L[454][8] = l_cell_wire[397];							inform_L[199][8] = l_cell_wire[398];							inform_L[455][8] = l_cell_wire[399];							inform_L[200][8] = l_cell_wire[400];							inform_L[456][8] = l_cell_wire[401];							inform_L[201][8] = l_cell_wire[402];							inform_L[457][8] = l_cell_wire[403];							inform_L[202][8] = l_cell_wire[404];							inform_L[458][8] = l_cell_wire[405];							inform_L[203][8] = l_cell_wire[406];							inform_L[459][8] = l_cell_wire[407];							inform_L[204][8] = l_cell_wire[408];							inform_L[460][8] = l_cell_wire[409];							inform_L[205][8] = l_cell_wire[410];							inform_L[461][8] = l_cell_wire[411];							inform_L[206][8] = l_cell_wire[412];							inform_L[462][8] = l_cell_wire[413];							inform_L[207][8] = l_cell_wire[414];							inform_L[463][8] = l_cell_wire[415];							inform_L[208][8] = l_cell_wire[416];							inform_L[464][8] = l_cell_wire[417];							inform_L[209][8] = l_cell_wire[418];							inform_L[465][8] = l_cell_wire[419];							inform_L[210][8] = l_cell_wire[420];							inform_L[466][8] = l_cell_wire[421];							inform_L[211][8] = l_cell_wire[422];							inform_L[467][8] = l_cell_wire[423];							inform_L[212][8] = l_cell_wire[424];							inform_L[468][8] = l_cell_wire[425];							inform_L[213][8] = l_cell_wire[426];							inform_L[469][8] = l_cell_wire[427];							inform_L[214][8] = l_cell_wire[428];							inform_L[470][8] = l_cell_wire[429];							inform_L[215][8] = l_cell_wire[430];							inform_L[471][8] = l_cell_wire[431];							inform_L[216][8] = l_cell_wire[432];							inform_L[472][8] = l_cell_wire[433];							inform_L[217][8] = l_cell_wire[434];							inform_L[473][8] = l_cell_wire[435];							inform_L[218][8] = l_cell_wire[436];							inform_L[474][8] = l_cell_wire[437];							inform_L[219][8] = l_cell_wire[438];							inform_L[475][8] = l_cell_wire[439];							inform_L[220][8] = l_cell_wire[440];							inform_L[476][8] = l_cell_wire[441];							inform_L[221][8] = l_cell_wire[442];							inform_L[477][8] = l_cell_wire[443];							inform_L[222][8] = l_cell_wire[444];							inform_L[478][8] = l_cell_wire[445];							inform_L[223][8] = l_cell_wire[446];							inform_L[479][8] = l_cell_wire[447];							inform_L[224][8] = l_cell_wire[448];							inform_L[480][8] = l_cell_wire[449];							inform_L[225][8] = l_cell_wire[450];							inform_L[481][8] = l_cell_wire[451];							inform_L[226][8] = l_cell_wire[452];							inform_L[482][8] = l_cell_wire[453];							inform_L[227][8] = l_cell_wire[454];							inform_L[483][8] = l_cell_wire[455];							inform_L[228][8] = l_cell_wire[456];							inform_L[484][8] = l_cell_wire[457];							inform_L[229][8] = l_cell_wire[458];							inform_L[485][8] = l_cell_wire[459];							inform_L[230][8] = l_cell_wire[460];							inform_L[486][8] = l_cell_wire[461];							inform_L[231][8] = l_cell_wire[462];							inform_L[487][8] = l_cell_wire[463];							inform_L[232][8] = l_cell_wire[464];							inform_L[488][8] = l_cell_wire[465];							inform_L[233][8] = l_cell_wire[466];							inform_L[489][8] = l_cell_wire[467];							inform_L[234][8] = l_cell_wire[468];							inform_L[490][8] = l_cell_wire[469];							inform_L[235][8] = l_cell_wire[470];							inform_L[491][8] = l_cell_wire[471];							inform_L[236][8] = l_cell_wire[472];							inform_L[492][8] = l_cell_wire[473];							inform_L[237][8] = l_cell_wire[474];							inform_L[493][8] = l_cell_wire[475];							inform_L[238][8] = l_cell_wire[476];							inform_L[494][8] = l_cell_wire[477];							inform_L[239][8] = l_cell_wire[478];							inform_L[495][8] = l_cell_wire[479];							inform_L[240][8] = l_cell_wire[480];							inform_L[496][8] = l_cell_wire[481];							inform_L[241][8] = l_cell_wire[482];							inform_L[497][8] = l_cell_wire[483];							inform_L[242][8] = l_cell_wire[484];							inform_L[498][8] = l_cell_wire[485];							inform_L[243][8] = l_cell_wire[486];							inform_L[499][8] = l_cell_wire[487];							inform_L[244][8] = l_cell_wire[488];							inform_L[500][8] = l_cell_wire[489];							inform_L[245][8] = l_cell_wire[490];							inform_L[501][8] = l_cell_wire[491];							inform_L[246][8] = l_cell_wire[492];							inform_L[502][8] = l_cell_wire[493];							inform_L[247][8] = l_cell_wire[494];							inform_L[503][8] = l_cell_wire[495];							inform_L[248][8] = l_cell_wire[496];							inform_L[504][8] = l_cell_wire[497];							inform_L[249][8] = l_cell_wire[498];							inform_L[505][8] = l_cell_wire[499];							inform_L[250][8] = l_cell_wire[500];							inform_L[506][8] = l_cell_wire[501];							inform_L[251][8] = l_cell_wire[502];							inform_L[507][8] = l_cell_wire[503];							inform_L[252][8] = l_cell_wire[504];							inform_L[508][8] = l_cell_wire[505];							inform_L[253][8] = l_cell_wire[506];							inform_L[509][8] = l_cell_wire[507];							inform_L[254][8] = l_cell_wire[508];							inform_L[510][8] = l_cell_wire[509];							inform_L[255][8] = l_cell_wire[510];							inform_L[511][8] = l_cell_wire[511];							inform_L[512][8] = l_cell_wire[512];							inform_L[768][8] = l_cell_wire[513];							inform_L[513][8] = l_cell_wire[514];							inform_L[769][8] = l_cell_wire[515];							inform_L[514][8] = l_cell_wire[516];							inform_L[770][8] = l_cell_wire[517];							inform_L[515][8] = l_cell_wire[518];							inform_L[771][8] = l_cell_wire[519];							inform_L[516][8] = l_cell_wire[520];							inform_L[772][8] = l_cell_wire[521];							inform_L[517][8] = l_cell_wire[522];							inform_L[773][8] = l_cell_wire[523];							inform_L[518][8] = l_cell_wire[524];							inform_L[774][8] = l_cell_wire[525];							inform_L[519][8] = l_cell_wire[526];							inform_L[775][8] = l_cell_wire[527];							inform_L[520][8] = l_cell_wire[528];							inform_L[776][8] = l_cell_wire[529];							inform_L[521][8] = l_cell_wire[530];							inform_L[777][8] = l_cell_wire[531];							inform_L[522][8] = l_cell_wire[532];							inform_L[778][8] = l_cell_wire[533];							inform_L[523][8] = l_cell_wire[534];							inform_L[779][8] = l_cell_wire[535];							inform_L[524][8] = l_cell_wire[536];							inform_L[780][8] = l_cell_wire[537];							inform_L[525][8] = l_cell_wire[538];							inform_L[781][8] = l_cell_wire[539];							inform_L[526][8] = l_cell_wire[540];							inform_L[782][8] = l_cell_wire[541];							inform_L[527][8] = l_cell_wire[542];							inform_L[783][8] = l_cell_wire[543];							inform_L[528][8] = l_cell_wire[544];							inform_L[784][8] = l_cell_wire[545];							inform_L[529][8] = l_cell_wire[546];							inform_L[785][8] = l_cell_wire[547];							inform_L[530][8] = l_cell_wire[548];							inform_L[786][8] = l_cell_wire[549];							inform_L[531][8] = l_cell_wire[550];							inform_L[787][8] = l_cell_wire[551];							inform_L[532][8] = l_cell_wire[552];							inform_L[788][8] = l_cell_wire[553];							inform_L[533][8] = l_cell_wire[554];							inform_L[789][8] = l_cell_wire[555];							inform_L[534][8] = l_cell_wire[556];							inform_L[790][8] = l_cell_wire[557];							inform_L[535][8] = l_cell_wire[558];							inform_L[791][8] = l_cell_wire[559];							inform_L[536][8] = l_cell_wire[560];							inform_L[792][8] = l_cell_wire[561];							inform_L[537][8] = l_cell_wire[562];							inform_L[793][8] = l_cell_wire[563];							inform_L[538][8] = l_cell_wire[564];							inform_L[794][8] = l_cell_wire[565];							inform_L[539][8] = l_cell_wire[566];							inform_L[795][8] = l_cell_wire[567];							inform_L[540][8] = l_cell_wire[568];							inform_L[796][8] = l_cell_wire[569];							inform_L[541][8] = l_cell_wire[570];							inform_L[797][8] = l_cell_wire[571];							inform_L[542][8] = l_cell_wire[572];							inform_L[798][8] = l_cell_wire[573];							inform_L[543][8] = l_cell_wire[574];							inform_L[799][8] = l_cell_wire[575];							inform_L[544][8] = l_cell_wire[576];							inform_L[800][8] = l_cell_wire[577];							inform_L[545][8] = l_cell_wire[578];							inform_L[801][8] = l_cell_wire[579];							inform_L[546][8] = l_cell_wire[580];							inform_L[802][8] = l_cell_wire[581];							inform_L[547][8] = l_cell_wire[582];							inform_L[803][8] = l_cell_wire[583];							inform_L[548][8] = l_cell_wire[584];							inform_L[804][8] = l_cell_wire[585];							inform_L[549][8] = l_cell_wire[586];							inform_L[805][8] = l_cell_wire[587];							inform_L[550][8] = l_cell_wire[588];							inform_L[806][8] = l_cell_wire[589];							inform_L[551][8] = l_cell_wire[590];							inform_L[807][8] = l_cell_wire[591];							inform_L[552][8] = l_cell_wire[592];							inform_L[808][8] = l_cell_wire[593];							inform_L[553][8] = l_cell_wire[594];							inform_L[809][8] = l_cell_wire[595];							inform_L[554][8] = l_cell_wire[596];							inform_L[810][8] = l_cell_wire[597];							inform_L[555][8] = l_cell_wire[598];							inform_L[811][8] = l_cell_wire[599];							inform_L[556][8] = l_cell_wire[600];							inform_L[812][8] = l_cell_wire[601];							inform_L[557][8] = l_cell_wire[602];							inform_L[813][8] = l_cell_wire[603];							inform_L[558][8] = l_cell_wire[604];							inform_L[814][8] = l_cell_wire[605];							inform_L[559][8] = l_cell_wire[606];							inform_L[815][8] = l_cell_wire[607];							inform_L[560][8] = l_cell_wire[608];							inform_L[816][8] = l_cell_wire[609];							inform_L[561][8] = l_cell_wire[610];							inform_L[817][8] = l_cell_wire[611];							inform_L[562][8] = l_cell_wire[612];							inform_L[818][8] = l_cell_wire[613];							inform_L[563][8] = l_cell_wire[614];							inform_L[819][8] = l_cell_wire[615];							inform_L[564][8] = l_cell_wire[616];							inform_L[820][8] = l_cell_wire[617];							inform_L[565][8] = l_cell_wire[618];							inform_L[821][8] = l_cell_wire[619];							inform_L[566][8] = l_cell_wire[620];							inform_L[822][8] = l_cell_wire[621];							inform_L[567][8] = l_cell_wire[622];							inform_L[823][8] = l_cell_wire[623];							inform_L[568][8] = l_cell_wire[624];							inform_L[824][8] = l_cell_wire[625];							inform_L[569][8] = l_cell_wire[626];							inform_L[825][8] = l_cell_wire[627];							inform_L[570][8] = l_cell_wire[628];							inform_L[826][8] = l_cell_wire[629];							inform_L[571][8] = l_cell_wire[630];							inform_L[827][8] = l_cell_wire[631];							inform_L[572][8] = l_cell_wire[632];							inform_L[828][8] = l_cell_wire[633];							inform_L[573][8] = l_cell_wire[634];							inform_L[829][8] = l_cell_wire[635];							inform_L[574][8] = l_cell_wire[636];							inform_L[830][8] = l_cell_wire[637];							inform_L[575][8] = l_cell_wire[638];							inform_L[831][8] = l_cell_wire[639];							inform_L[576][8] = l_cell_wire[640];							inform_L[832][8] = l_cell_wire[641];							inform_L[577][8] = l_cell_wire[642];							inform_L[833][8] = l_cell_wire[643];							inform_L[578][8] = l_cell_wire[644];							inform_L[834][8] = l_cell_wire[645];							inform_L[579][8] = l_cell_wire[646];							inform_L[835][8] = l_cell_wire[647];							inform_L[580][8] = l_cell_wire[648];							inform_L[836][8] = l_cell_wire[649];							inform_L[581][8] = l_cell_wire[650];							inform_L[837][8] = l_cell_wire[651];							inform_L[582][8] = l_cell_wire[652];							inform_L[838][8] = l_cell_wire[653];							inform_L[583][8] = l_cell_wire[654];							inform_L[839][8] = l_cell_wire[655];							inform_L[584][8] = l_cell_wire[656];							inform_L[840][8] = l_cell_wire[657];							inform_L[585][8] = l_cell_wire[658];							inform_L[841][8] = l_cell_wire[659];							inform_L[586][8] = l_cell_wire[660];							inform_L[842][8] = l_cell_wire[661];							inform_L[587][8] = l_cell_wire[662];							inform_L[843][8] = l_cell_wire[663];							inform_L[588][8] = l_cell_wire[664];							inform_L[844][8] = l_cell_wire[665];							inform_L[589][8] = l_cell_wire[666];							inform_L[845][8] = l_cell_wire[667];							inform_L[590][8] = l_cell_wire[668];							inform_L[846][8] = l_cell_wire[669];							inform_L[591][8] = l_cell_wire[670];							inform_L[847][8] = l_cell_wire[671];							inform_L[592][8] = l_cell_wire[672];							inform_L[848][8] = l_cell_wire[673];							inform_L[593][8] = l_cell_wire[674];							inform_L[849][8] = l_cell_wire[675];							inform_L[594][8] = l_cell_wire[676];							inform_L[850][8] = l_cell_wire[677];							inform_L[595][8] = l_cell_wire[678];							inform_L[851][8] = l_cell_wire[679];							inform_L[596][8] = l_cell_wire[680];							inform_L[852][8] = l_cell_wire[681];							inform_L[597][8] = l_cell_wire[682];							inform_L[853][8] = l_cell_wire[683];							inform_L[598][8] = l_cell_wire[684];							inform_L[854][8] = l_cell_wire[685];							inform_L[599][8] = l_cell_wire[686];							inform_L[855][8] = l_cell_wire[687];							inform_L[600][8] = l_cell_wire[688];							inform_L[856][8] = l_cell_wire[689];							inform_L[601][8] = l_cell_wire[690];							inform_L[857][8] = l_cell_wire[691];							inform_L[602][8] = l_cell_wire[692];							inform_L[858][8] = l_cell_wire[693];							inform_L[603][8] = l_cell_wire[694];							inform_L[859][8] = l_cell_wire[695];							inform_L[604][8] = l_cell_wire[696];							inform_L[860][8] = l_cell_wire[697];							inform_L[605][8] = l_cell_wire[698];							inform_L[861][8] = l_cell_wire[699];							inform_L[606][8] = l_cell_wire[700];							inform_L[862][8] = l_cell_wire[701];							inform_L[607][8] = l_cell_wire[702];							inform_L[863][8] = l_cell_wire[703];							inform_L[608][8] = l_cell_wire[704];							inform_L[864][8] = l_cell_wire[705];							inform_L[609][8] = l_cell_wire[706];							inform_L[865][8] = l_cell_wire[707];							inform_L[610][8] = l_cell_wire[708];							inform_L[866][8] = l_cell_wire[709];							inform_L[611][8] = l_cell_wire[710];							inform_L[867][8] = l_cell_wire[711];							inform_L[612][8] = l_cell_wire[712];							inform_L[868][8] = l_cell_wire[713];							inform_L[613][8] = l_cell_wire[714];							inform_L[869][8] = l_cell_wire[715];							inform_L[614][8] = l_cell_wire[716];							inform_L[870][8] = l_cell_wire[717];							inform_L[615][8] = l_cell_wire[718];							inform_L[871][8] = l_cell_wire[719];							inform_L[616][8] = l_cell_wire[720];							inform_L[872][8] = l_cell_wire[721];							inform_L[617][8] = l_cell_wire[722];							inform_L[873][8] = l_cell_wire[723];							inform_L[618][8] = l_cell_wire[724];							inform_L[874][8] = l_cell_wire[725];							inform_L[619][8] = l_cell_wire[726];							inform_L[875][8] = l_cell_wire[727];							inform_L[620][8] = l_cell_wire[728];							inform_L[876][8] = l_cell_wire[729];							inform_L[621][8] = l_cell_wire[730];							inform_L[877][8] = l_cell_wire[731];							inform_L[622][8] = l_cell_wire[732];							inform_L[878][8] = l_cell_wire[733];							inform_L[623][8] = l_cell_wire[734];							inform_L[879][8] = l_cell_wire[735];							inform_L[624][8] = l_cell_wire[736];							inform_L[880][8] = l_cell_wire[737];							inform_L[625][8] = l_cell_wire[738];							inform_L[881][8] = l_cell_wire[739];							inform_L[626][8] = l_cell_wire[740];							inform_L[882][8] = l_cell_wire[741];							inform_L[627][8] = l_cell_wire[742];							inform_L[883][8] = l_cell_wire[743];							inform_L[628][8] = l_cell_wire[744];							inform_L[884][8] = l_cell_wire[745];							inform_L[629][8] = l_cell_wire[746];							inform_L[885][8] = l_cell_wire[747];							inform_L[630][8] = l_cell_wire[748];							inform_L[886][8] = l_cell_wire[749];							inform_L[631][8] = l_cell_wire[750];							inform_L[887][8] = l_cell_wire[751];							inform_L[632][8] = l_cell_wire[752];							inform_L[888][8] = l_cell_wire[753];							inform_L[633][8] = l_cell_wire[754];							inform_L[889][8] = l_cell_wire[755];							inform_L[634][8] = l_cell_wire[756];							inform_L[890][8] = l_cell_wire[757];							inform_L[635][8] = l_cell_wire[758];							inform_L[891][8] = l_cell_wire[759];							inform_L[636][8] = l_cell_wire[760];							inform_L[892][8] = l_cell_wire[761];							inform_L[637][8] = l_cell_wire[762];							inform_L[893][8] = l_cell_wire[763];							inform_L[638][8] = l_cell_wire[764];							inform_L[894][8] = l_cell_wire[765];							inform_L[639][8] = l_cell_wire[766];							inform_L[895][8] = l_cell_wire[767];							inform_L[640][8] = l_cell_wire[768];							inform_L[896][8] = l_cell_wire[769];							inform_L[641][8] = l_cell_wire[770];							inform_L[897][8] = l_cell_wire[771];							inform_L[642][8] = l_cell_wire[772];							inform_L[898][8] = l_cell_wire[773];							inform_L[643][8] = l_cell_wire[774];							inform_L[899][8] = l_cell_wire[775];							inform_L[644][8] = l_cell_wire[776];							inform_L[900][8] = l_cell_wire[777];							inform_L[645][8] = l_cell_wire[778];							inform_L[901][8] = l_cell_wire[779];							inform_L[646][8] = l_cell_wire[780];							inform_L[902][8] = l_cell_wire[781];							inform_L[647][8] = l_cell_wire[782];							inform_L[903][8] = l_cell_wire[783];							inform_L[648][8] = l_cell_wire[784];							inform_L[904][8] = l_cell_wire[785];							inform_L[649][8] = l_cell_wire[786];							inform_L[905][8] = l_cell_wire[787];							inform_L[650][8] = l_cell_wire[788];							inform_L[906][8] = l_cell_wire[789];							inform_L[651][8] = l_cell_wire[790];							inform_L[907][8] = l_cell_wire[791];							inform_L[652][8] = l_cell_wire[792];							inform_L[908][8] = l_cell_wire[793];							inform_L[653][8] = l_cell_wire[794];							inform_L[909][8] = l_cell_wire[795];							inform_L[654][8] = l_cell_wire[796];							inform_L[910][8] = l_cell_wire[797];							inform_L[655][8] = l_cell_wire[798];							inform_L[911][8] = l_cell_wire[799];							inform_L[656][8] = l_cell_wire[800];							inform_L[912][8] = l_cell_wire[801];							inform_L[657][8] = l_cell_wire[802];							inform_L[913][8] = l_cell_wire[803];							inform_L[658][8] = l_cell_wire[804];							inform_L[914][8] = l_cell_wire[805];							inform_L[659][8] = l_cell_wire[806];							inform_L[915][8] = l_cell_wire[807];							inform_L[660][8] = l_cell_wire[808];							inform_L[916][8] = l_cell_wire[809];							inform_L[661][8] = l_cell_wire[810];							inform_L[917][8] = l_cell_wire[811];							inform_L[662][8] = l_cell_wire[812];							inform_L[918][8] = l_cell_wire[813];							inform_L[663][8] = l_cell_wire[814];							inform_L[919][8] = l_cell_wire[815];							inform_L[664][8] = l_cell_wire[816];							inform_L[920][8] = l_cell_wire[817];							inform_L[665][8] = l_cell_wire[818];							inform_L[921][8] = l_cell_wire[819];							inform_L[666][8] = l_cell_wire[820];							inform_L[922][8] = l_cell_wire[821];							inform_L[667][8] = l_cell_wire[822];							inform_L[923][8] = l_cell_wire[823];							inform_L[668][8] = l_cell_wire[824];							inform_L[924][8] = l_cell_wire[825];							inform_L[669][8] = l_cell_wire[826];							inform_L[925][8] = l_cell_wire[827];							inform_L[670][8] = l_cell_wire[828];							inform_L[926][8] = l_cell_wire[829];							inform_L[671][8] = l_cell_wire[830];							inform_L[927][8] = l_cell_wire[831];							inform_L[672][8] = l_cell_wire[832];							inform_L[928][8] = l_cell_wire[833];							inform_L[673][8] = l_cell_wire[834];							inform_L[929][8] = l_cell_wire[835];							inform_L[674][8] = l_cell_wire[836];							inform_L[930][8] = l_cell_wire[837];							inform_L[675][8] = l_cell_wire[838];							inform_L[931][8] = l_cell_wire[839];							inform_L[676][8] = l_cell_wire[840];							inform_L[932][8] = l_cell_wire[841];							inform_L[677][8] = l_cell_wire[842];							inform_L[933][8] = l_cell_wire[843];							inform_L[678][8] = l_cell_wire[844];							inform_L[934][8] = l_cell_wire[845];							inform_L[679][8] = l_cell_wire[846];							inform_L[935][8] = l_cell_wire[847];							inform_L[680][8] = l_cell_wire[848];							inform_L[936][8] = l_cell_wire[849];							inform_L[681][8] = l_cell_wire[850];							inform_L[937][8] = l_cell_wire[851];							inform_L[682][8] = l_cell_wire[852];							inform_L[938][8] = l_cell_wire[853];							inform_L[683][8] = l_cell_wire[854];							inform_L[939][8] = l_cell_wire[855];							inform_L[684][8] = l_cell_wire[856];							inform_L[940][8] = l_cell_wire[857];							inform_L[685][8] = l_cell_wire[858];							inform_L[941][8] = l_cell_wire[859];							inform_L[686][8] = l_cell_wire[860];							inform_L[942][8] = l_cell_wire[861];							inform_L[687][8] = l_cell_wire[862];							inform_L[943][8] = l_cell_wire[863];							inform_L[688][8] = l_cell_wire[864];							inform_L[944][8] = l_cell_wire[865];							inform_L[689][8] = l_cell_wire[866];							inform_L[945][8] = l_cell_wire[867];							inform_L[690][8] = l_cell_wire[868];							inform_L[946][8] = l_cell_wire[869];							inform_L[691][8] = l_cell_wire[870];							inform_L[947][8] = l_cell_wire[871];							inform_L[692][8] = l_cell_wire[872];							inform_L[948][8] = l_cell_wire[873];							inform_L[693][8] = l_cell_wire[874];							inform_L[949][8] = l_cell_wire[875];							inform_L[694][8] = l_cell_wire[876];							inform_L[950][8] = l_cell_wire[877];							inform_L[695][8] = l_cell_wire[878];							inform_L[951][8] = l_cell_wire[879];							inform_L[696][8] = l_cell_wire[880];							inform_L[952][8] = l_cell_wire[881];							inform_L[697][8] = l_cell_wire[882];							inform_L[953][8] = l_cell_wire[883];							inform_L[698][8] = l_cell_wire[884];							inform_L[954][8] = l_cell_wire[885];							inform_L[699][8] = l_cell_wire[886];							inform_L[955][8] = l_cell_wire[887];							inform_L[700][8] = l_cell_wire[888];							inform_L[956][8] = l_cell_wire[889];							inform_L[701][8] = l_cell_wire[890];							inform_L[957][8] = l_cell_wire[891];							inform_L[702][8] = l_cell_wire[892];							inform_L[958][8] = l_cell_wire[893];							inform_L[703][8] = l_cell_wire[894];							inform_L[959][8] = l_cell_wire[895];							inform_L[704][8] = l_cell_wire[896];							inform_L[960][8] = l_cell_wire[897];							inform_L[705][8] = l_cell_wire[898];							inform_L[961][8] = l_cell_wire[899];							inform_L[706][8] = l_cell_wire[900];							inform_L[962][8] = l_cell_wire[901];							inform_L[707][8] = l_cell_wire[902];							inform_L[963][8] = l_cell_wire[903];							inform_L[708][8] = l_cell_wire[904];							inform_L[964][8] = l_cell_wire[905];							inform_L[709][8] = l_cell_wire[906];							inform_L[965][8] = l_cell_wire[907];							inform_L[710][8] = l_cell_wire[908];							inform_L[966][8] = l_cell_wire[909];							inform_L[711][8] = l_cell_wire[910];							inform_L[967][8] = l_cell_wire[911];							inform_L[712][8] = l_cell_wire[912];							inform_L[968][8] = l_cell_wire[913];							inform_L[713][8] = l_cell_wire[914];							inform_L[969][8] = l_cell_wire[915];							inform_L[714][8] = l_cell_wire[916];							inform_L[970][8] = l_cell_wire[917];							inform_L[715][8] = l_cell_wire[918];							inform_L[971][8] = l_cell_wire[919];							inform_L[716][8] = l_cell_wire[920];							inform_L[972][8] = l_cell_wire[921];							inform_L[717][8] = l_cell_wire[922];							inform_L[973][8] = l_cell_wire[923];							inform_L[718][8] = l_cell_wire[924];							inform_L[974][8] = l_cell_wire[925];							inform_L[719][8] = l_cell_wire[926];							inform_L[975][8] = l_cell_wire[927];							inform_L[720][8] = l_cell_wire[928];							inform_L[976][8] = l_cell_wire[929];							inform_L[721][8] = l_cell_wire[930];							inform_L[977][8] = l_cell_wire[931];							inform_L[722][8] = l_cell_wire[932];							inform_L[978][8] = l_cell_wire[933];							inform_L[723][8] = l_cell_wire[934];							inform_L[979][8] = l_cell_wire[935];							inform_L[724][8] = l_cell_wire[936];							inform_L[980][8] = l_cell_wire[937];							inform_L[725][8] = l_cell_wire[938];							inform_L[981][8] = l_cell_wire[939];							inform_L[726][8] = l_cell_wire[940];							inform_L[982][8] = l_cell_wire[941];							inform_L[727][8] = l_cell_wire[942];							inform_L[983][8] = l_cell_wire[943];							inform_L[728][8] = l_cell_wire[944];							inform_L[984][8] = l_cell_wire[945];							inform_L[729][8] = l_cell_wire[946];							inform_L[985][8] = l_cell_wire[947];							inform_L[730][8] = l_cell_wire[948];							inform_L[986][8] = l_cell_wire[949];							inform_L[731][8] = l_cell_wire[950];							inform_L[987][8] = l_cell_wire[951];							inform_L[732][8] = l_cell_wire[952];							inform_L[988][8] = l_cell_wire[953];							inform_L[733][8] = l_cell_wire[954];							inform_L[989][8] = l_cell_wire[955];							inform_L[734][8] = l_cell_wire[956];							inform_L[990][8] = l_cell_wire[957];							inform_L[735][8] = l_cell_wire[958];							inform_L[991][8] = l_cell_wire[959];							inform_L[736][8] = l_cell_wire[960];							inform_L[992][8] = l_cell_wire[961];							inform_L[737][8] = l_cell_wire[962];							inform_L[993][8] = l_cell_wire[963];							inform_L[738][8] = l_cell_wire[964];							inform_L[994][8] = l_cell_wire[965];							inform_L[739][8] = l_cell_wire[966];							inform_L[995][8] = l_cell_wire[967];							inform_L[740][8] = l_cell_wire[968];							inform_L[996][8] = l_cell_wire[969];							inform_L[741][8] = l_cell_wire[970];							inform_L[997][8] = l_cell_wire[971];							inform_L[742][8] = l_cell_wire[972];							inform_L[998][8] = l_cell_wire[973];							inform_L[743][8] = l_cell_wire[974];							inform_L[999][8] = l_cell_wire[975];							inform_L[744][8] = l_cell_wire[976];							inform_L[1000][8] = l_cell_wire[977];							inform_L[745][8] = l_cell_wire[978];							inform_L[1001][8] = l_cell_wire[979];							inform_L[746][8] = l_cell_wire[980];							inform_L[1002][8] = l_cell_wire[981];							inform_L[747][8] = l_cell_wire[982];							inform_L[1003][8] = l_cell_wire[983];							inform_L[748][8] = l_cell_wire[984];							inform_L[1004][8] = l_cell_wire[985];							inform_L[749][8] = l_cell_wire[986];							inform_L[1005][8] = l_cell_wire[987];							inform_L[750][8] = l_cell_wire[988];							inform_L[1006][8] = l_cell_wire[989];							inform_L[751][8] = l_cell_wire[990];							inform_L[1007][8] = l_cell_wire[991];							inform_L[752][8] = l_cell_wire[992];							inform_L[1008][8] = l_cell_wire[993];							inform_L[753][8] = l_cell_wire[994];							inform_L[1009][8] = l_cell_wire[995];							inform_L[754][8] = l_cell_wire[996];							inform_L[1010][8] = l_cell_wire[997];							inform_L[755][8] = l_cell_wire[998];							inform_L[1011][8] = l_cell_wire[999];							inform_L[756][8] = l_cell_wire[1000];							inform_L[1012][8] = l_cell_wire[1001];							inform_L[757][8] = l_cell_wire[1002];							inform_L[1013][8] = l_cell_wire[1003];							inform_L[758][8] = l_cell_wire[1004];							inform_L[1014][8] = l_cell_wire[1005];							inform_L[759][8] = l_cell_wire[1006];							inform_L[1015][8] = l_cell_wire[1007];							inform_L[760][8] = l_cell_wire[1008];							inform_L[1016][8] = l_cell_wire[1009];							inform_L[761][8] = l_cell_wire[1010];							inform_L[1017][8] = l_cell_wire[1011];							inform_L[762][8] = l_cell_wire[1012];							inform_L[1018][8] = l_cell_wire[1013];							inform_L[763][8] = l_cell_wire[1014];							inform_L[1019][8] = l_cell_wire[1015];							inform_L[764][8] = l_cell_wire[1016];							inform_L[1020][8] = l_cell_wire[1017];							inform_L[765][8] = l_cell_wire[1018];							inform_L[1021][8] = l_cell_wire[1019];							inform_L[766][8] = l_cell_wire[1020];							inform_L[1022][8] = l_cell_wire[1021];							inform_L[767][8] = l_cell_wire[1022];							inform_L[1023][8] = l_cell_wire[1023];						end
						10:						begin							inform_R[0][10] = r_cell_wire[0];							inform_R[512][10] = r_cell_wire[1];							inform_R[1][10] = r_cell_wire[2];							inform_R[513][10] = r_cell_wire[3];							inform_R[2][10] = r_cell_wire[4];							inform_R[514][10] = r_cell_wire[5];							inform_R[3][10] = r_cell_wire[6];							inform_R[515][10] = r_cell_wire[7];							inform_R[4][10] = r_cell_wire[8];							inform_R[516][10] = r_cell_wire[9];							inform_R[5][10] = r_cell_wire[10];							inform_R[517][10] = r_cell_wire[11];							inform_R[6][10] = r_cell_wire[12];							inform_R[518][10] = r_cell_wire[13];							inform_R[7][10] = r_cell_wire[14];							inform_R[519][10] = r_cell_wire[15];							inform_R[8][10] = r_cell_wire[16];							inform_R[520][10] = r_cell_wire[17];							inform_R[9][10] = r_cell_wire[18];							inform_R[521][10] = r_cell_wire[19];							inform_R[10][10] = r_cell_wire[20];							inform_R[522][10] = r_cell_wire[21];							inform_R[11][10] = r_cell_wire[22];							inform_R[523][10] = r_cell_wire[23];							inform_R[12][10] = r_cell_wire[24];							inform_R[524][10] = r_cell_wire[25];							inform_R[13][10] = r_cell_wire[26];							inform_R[525][10] = r_cell_wire[27];							inform_R[14][10] = r_cell_wire[28];							inform_R[526][10] = r_cell_wire[29];							inform_R[15][10] = r_cell_wire[30];							inform_R[527][10] = r_cell_wire[31];							inform_R[16][10] = r_cell_wire[32];							inform_R[528][10] = r_cell_wire[33];							inform_R[17][10] = r_cell_wire[34];							inform_R[529][10] = r_cell_wire[35];							inform_R[18][10] = r_cell_wire[36];							inform_R[530][10] = r_cell_wire[37];							inform_R[19][10] = r_cell_wire[38];							inform_R[531][10] = r_cell_wire[39];							inform_R[20][10] = r_cell_wire[40];							inform_R[532][10] = r_cell_wire[41];							inform_R[21][10] = r_cell_wire[42];							inform_R[533][10] = r_cell_wire[43];							inform_R[22][10] = r_cell_wire[44];							inform_R[534][10] = r_cell_wire[45];							inform_R[23][10] = r_cell_wire[46];							inform_R[535][10] = r_cell_wire[47];							inform_R[24][10] = r_cell_wire[48];							inform_R[536][10] = r_cell_wire[49];							inform_R[25][10] = r_cell_wire[50];							inform_R[537][10] = r_cell_wire[51];							inform_R[26][10] = r_cell_wire[52];							inform_R[538][10] = r_cell_wire[53];							inform_R[27][10] = r_cell_wire[54];							inform_R[539][10] = r_cell_wire[55];							inform_R[28][10] = r_cell_wire[56];							inform_R[540][10] = r_cell_wire[57];							inform_R[29][10] = r_cell_wire[58];							inform_R[541][10] = r_cell_wire[59];							inform_R[30][10] = r_cell_wire[60];							inform_R[542][10] = r_cell_wire[61];							inform_R[31][10] = r_cell_wire[62];							inform_R[543][10] = r_cell_wire[63];							inform_R[32][10] = r_cell_wire[64];							inform_R[544][10] = r_cell_wire[65];							inform_R[33][10] = r_cell_wire[66];							inform_R[545][10] = r_cell_wire[67];							inform_R[34][10] = r_cell_wire[68];							inform_R[546][10] = r_cell_wire[69];							inform_R[35][10] = r_cell_wire[70];							inform_R[547][10] = r_cell_wire[71];							inform_R[36][10] = r_cell_wire[72];							inform_R[548][10] = r_cell_wire[73];							inform_R[37][10] = r_cell_wire[74];							inform_R[549][10] = r_cell_wire[75];							inform_R[38][10] = r_cell_wire[76];							inform_R[550][10] = r_cell_wire[77];							inform_R[39][10] = r_cell_wire[78];							inform_R[551][10] = r_cell_wire[79];							inform_R[40][10] = r_cell_wire[80];							inform_R[552][10] = r_cell_wire[81];							inform_R[41][10] = r_cell_wire[82];							inform_R[553][10] = r_cell_wire[83];							inform_R[42][10] = r_cell_wire[84];							inform_R[554][10] = r_cell_wire[85];							inform_R[43][10] = r_cell_wire[86];							inform_R[555][10] = r_cell_wire[87];							inform_R[44][10] = r_cell_wire[88];							inform_R[556][10] = r_cell_wire[89];							inform_R[45][10] = r_cell_wire[90];							inform_R[557][10] = r_cell_wire[91];							inform_R[46][10] = r_cell_wire[92];							inform_R[558][10] = r_cell_wire[93];							inform_R[47][10] = r_cell_wire[94];							inform_R[559][10] = r_cell_wire[95];							inform_R[48][10] = r_cell_wire[96];							inform_R[560][10] = r_cell_wire[97];							inform_R[49][10] = r_cell_wire[98];							inform_R[561][10] = r_cell_wire[99];							inform_R[50][10] = r_cell_wire[100];							inform_R[562][10] = r_cell_wire[101];							inform_R[51][10] = r_cell_wire[102];							inform_R[563][10] = r_cell_wire[103];							inform_R[52][10] = r_cell_wire[104];							inform_R[564][10] = r_cell_wire[105];							inform_R[53][10] = r_cell_wire[106];							inform_R[565][10] = r_cell_wire[107];							inform_R[54][10] = r_cell_wire[108];							inform_R[566][10] = r_cell_wire[109];							inform_R[55][10] = r_cell_wire[110];							inform_R[567][10] = r_cell_wire[111];							inform_R[56][10] = r_cell_wire[112];							inform_R[568][10] = r_cell_wire[113];							inform_R[57][10] = r_cell_wire[114];							inform_R[569][10] = r_cell_wire[115];							inform_R[58][10] = r_cell_wire[116];							inform_R[570][10] = r_cell_wire[117];							inform_R[59][10] = r_cell_wire[118];							inform_R[571][10] = r_cell_wire[119];							inform_R[60][10] = r_cell_wire[120];							inform_R[572][10] = r_cell_wire[121];							inform_R[61][10] = r_cell_wire[122];							inform_R[573][10] = r_cell_wire[123];							inform_R[62][10] = r_cell_wire[124];							inform_R[574][10] = r_cell_wire[125];							inform_R[63][10] = r_cell_wire[126];							inform_R[575][10] = r_cell_wire[127];							inform_R[64][10] = r_cell_wire[128];							inform_R[576][10] = r_cell_wire[129];							inform_R[65][10] = r_cell_wire[130];							inform_R[577][10] = r_cell_wire[131];							inform_R[66][10] = r_cell_wire[132];							inform_R[578][10] = r_cell_wire[133];							inform_R[67][10] = r_cell_wire[134];							inform_R[579][10] = r_cell_wire[135];							inform_R[68][10] = r_cell_wire[136];							inform_R[580][10] = r_cell_wire[137];							inform_R[69][10] = r_cell_wire[138];							inform_R[581][10] = r_cell_wire[139];							inform_R[70][10] = r_cell_wire[140];							inform_R[582][10] = r_cell_wire[141];							inform_R[71][10] = r_cell_wire[142];							inform_R[583][10] = r_cell_wire[143];							inform_R[72][10] = r_cell_wire[144];							inform_R[584][10] = r_cell_wire[145];							inform_R[73][10] = r_cell_wire[146];							inform_R[585][10] = r_cell_wire[147];							inform_R[74][10] = r_cell_wire[148];							inform_R[586][10] = r_cell_wire[149];							inform_R[75][10] = r_cell_wire[150];							inform_R[587][10] = r_cell_wire[151];							inform_R[76][10] = r_cell_wire[152];							inform_R[588][10] = r_cell_wire[153];							inform_R[77][10] = r_cell_wire[154];							inform_R[589][10] = r_cell_wire[155];							inform_R[78][10] = r_cell_wire[156];							inform_R[590][10] = r_cell_wire[157];							inform_R[79][10] = r_cell_wire[158];							inform_R[591][10] = r_cell_wire[159];							inform_R[80][10] = r_cell_wire[160];							inform_R[592][10] = r_cell_wire[161];							inform_R[81][10] = r_cell_wire[162];							inform_R[593][10] = r_cell_wire[163];							inform_R[82][10] = r_cell_wire[164];							inform_R[594][10] = r_cell_wire[165];							inform_R[83][10] = r_cell_wire[166];							inform_R[595][10] = r_cell_wire[167];							inform_R[84][10] = r_cell_wire[168];							inform_R[596][10] = r_cell_wire[169];							inform_R[85][10] = r_cell_wire[170];							inform_R[597][10] = r_cell_wire[171];							inform_R[86][10] = r_cell_wire[172];							inform_R[598][10] = r_cell_wire[173];							inform_R[87][10] = r_cell_wire[174];							inform_R[599][10] = r_cell_wire[175];							inform_R[88][10] = r_cell_wire[176];							inform_R[600][10] = r_cell_wire[177];							inform_R[89][10] = r_cell_wire[178];							inform_R[601][10] = r_cell_wire[179];							inform_R[90][10] = r_cell_wire[180];							inform_R[602][10] = r_cell_wire[181];							inform_R[91][10] = r_cell_wire[182];							inform_R[603][10] = r_cell_wire[183];							inform_R[92][10] = r_cell_wire[184];							inform_R[604][10] = r_cell_wire[185];							inform_R[93][10] = r_cell_wire[186];							inform_R[605][10] = r_cell_wire[187];							inform_R[94][10] = r_cell_wire[188];							inform_R[606][10] = r_cell_wire[189];							inform_R[95][10] = r_cell_wire[190];							inform_R[607][10] = r_cell_wire[191];							inform_R[96][10] = r_cell_wire[192];							inform_R[608][10] = r_cell_wire[193];							inform_R[97][10] = r_cell_wire[194];							inform_R[609][10] = r_cell_wire[195];							inform_R[98][10] = r_cell_wire[196];							inform_R[610][10] = r_cell_wire[197];							inform_R[99][10] = r_cell_wire[198];							inform_R[611][10] = r_cell_wire[199];							inform_R[100][10] = r_cell_wire[200];							inform_R[612][10] = r_cell_wire[201];							inform_R[101][10] = r_cell_wire[202];							inform_R[613][10] = r_cell_wire[203];							inform_R[102][10] = r_cell_wire[204];							inform_R[614][10] = r_cell_wire[205];							inform_R[103][10] = r_cell_wire[206];							inform_R[615][10] = r_cell_wire[207];							inform_R[104][10] = r_cell_wire[208];							inform_R[616][10] = r_cell_wire[209];							inform_R[105][10] = r_cell_wire[210];							inform_R[617][10] = r_cell_wire[211];							inform_R[106][10] = r_cell_wire[212];							inform_R[618][10] = r_cell_wire[213];							inform_R[107][10] = r_cell_wire[214];							inform_R[619][10] = r_cell_wire[215];							inform_R[108][10] = r_cell_wire[216];							inform_R[620][10] = r_cell_wire[217];							inform_R[109][10] = r_cell_wire[218];							inform_R[621][10] = r_cell_wire[219];							inform_R[110][10] = r_cell_wire[220];							inform_R[622][10] = r_cell_wire[221];							inform_R[111][10] = r_cell_wire[222];							inform_R[623][10] = r_cell_wire[223];							inform_R[112][10] = r_cell_wire[224];							inform_R[624][10] = r_cell_wire[225];							inform_R[113][10] = r_cell_wire[226];							inform_R[625][10] = r_cell_wire[227];							inform_R[114][10] = r_cell_wire[228];							inform_R[626][10] = r_cell_wire[229];							inform_R[115][10] = r_cell_wire[230];							inform_R[627][10] = r_cell_wire[231];							inform_R[116][10] = r_cell_wire[232];							inform_R[628][10] = r_cell_wire[233];							inform_R[117][10] = r_cell_wire[234];							inform_R[629][10] = r_cell_wire[235];							inform_R[118][10] = r_cell_wire[236];							inform_R[630][10] = r_cell_wire[237];							inform_R[119][10] = r_cell_wire[238];							inform_R[631][10] = r_cell_wire[239];							inform_R[120][10] = r_cell_wire[240];							inform_R[632][10] = r_cell_wire[241];							inform_R[121][10] = r_cell_wire[242];							inform_R[633][10] = r_cell_wire[243];							inform_R[122][10] = r_cell_wire[244];							inform_R[634][10] = r_cell_wire[245];							inform_R[123][10] = r_cell_wire[246];							inform_R[635][10] = r_cell_wire[247];							inform_R[124][10] = r_cell_wire[248];							inform_R[636][10] = r_cell_wire[249];							inform_R[125][10] = r_cell_wire[250];							inform_R[637][10] = r_cell_wire[251];							inform_R[126][10] = r_cell_wire[252];							inform_R[638][10] = r_cell_wire[253];							inform_R[127][10] = r_cell_wire[254];							inform_R[639][10] = r_cell_wire[255];							inform_R[128][10] = r_cell_wire[256];							inform_R[640][10] = r_cell_wire[257];							inform_R[129][10] = r_cell_wire[258];							inform_R[641][10] = r_cell_wire[259];							inform_R[130][10] = r_cell_wire[260];							inform_R[642][10] = r_cell_wire[261];							inform_R[131][10] = r_cell_wire[262];							inform_R[643][10] = r_cell_wire[263];							inform_R[132][10] = r_cell_wire[264];							inform_R[644][10] = r_cell_wire[265];							inform_R[133][10] = r_cell_wire[266];							inform_R[645][10] = r_cell_wire[267];							inform_R[134][10] = r_cell_wire[268];							inform_R[646][10] = r_cell_wire[269];							inform_R[135][10] = r_cell_wire[270];							inform_R[647][10] = r_cell_wire[271];							inform_R[136][10] = r_cell_wire[272];							inform_R[648][10] = r_cell_wire[273];							inform_R[137][10] = r_cell_wire[274];							inform_R[649][10] = r_cell_wire[275];							inform_R[138][10] = r_cell_wire[276];							inform_R[650][10] = r_cell_wire[277];							inform_R[139][10] = r_cell_wire[278];							inform_R[651][10] = r_cell_wire[279];							inform_R[140][10] = r_cell_wire[280];							inform_R[652][10] = r_cell_wire[281];							inform_R[141][10] = r_cell_wire[282];							inform_R[653][10] = r_cell_wire[283];							inform_R[142][10] = r_cell_wire[284];							inform_R[654][10] = r_cell_wire[285];							inform_R[143][10] = r_cell_wire[286];							inform_R[655][10] = r_cell_wire[287];							inform_R[144][10] = r_cell_wire[288];							inform_R[656][10] = r_cell_wire[289];							inform_R[145][10] = r_cell_wire[290];							inform_R[657][10] = r_cell_wire[291];							inform_R[146][10] = r_cell_wire[292];							inform_R[658][10] = r_cell_wire[293];							inform_R[147][10] = r_cell_wire[294];							inform_R[659][10] = r_cell_wire[295];							inform_R[148][10] = r_cell_wire[296];							inform_R[660][10] = r_cell_wire[297];							inform_R[149][10] = r_cell_wire[298];							inform_R[661][10] = r_cell_wire[299];							inform_R[150][10] = r_cell_wire[300];							inform_R[662][10] = r_cell_wire[301];							inform_R[151][10] = r_cell_wire[302];							inform_R[663][10] = r_cell_wire[303];							inform_R[152][10] = r_cell_wire[304];							inform_R[664][10] = r_cell_wire[305];							inform_R[153][10] = r_cell_wire[306];							inform_R[665][10] = r_cell_wire[307];							inform_R[154][10] = r_cell_wire[308];							inform_R[666][10] = r_cell_wire[309];							inform_R[155][10] = r_cell_wire[310];							inform_R[667][10] = r_cell_wire[311];							inform_R[156][10] = r_cell_wire[312];							inform_R[668][10] = r_cell_wire[313];							inform_R[157][10] = r_cell_wire[314];							inform_R[669][10] = r_cell_wire[315];							inform_R[158][10] = r_cell_wire[316];							inform_R[670][10] = r_cell_wire[317];							inform_R[159][10] = r_cell_wire[318];							inform_R[671][10] = r_cell_wire[319];							inform_R[160][10] = r_cell_wire[320];							inform_R[672][10] = r_cell_wire[321];							inform_R[161][10] = r_cell_wire[322];							inform_R[673][10] = r_cell_wire[323];							inform_R[162][10] = r_cell_wire[324];							inform_R[674][10] = r_cell_wire[325];							inform_R[163][10] = r_cell_wire[326];							inform_R[675][10] = r_cell_wire[327];							inform_R[164][10] = r_cell_wire[328];							inform_R[676][10] = r_cell_wire[329];							inform_R[165][10] = r_cell_wire[330];							inform_R[677][10] = r_cell_wire[331];							inform_R[166][10] = r_cell_wire[332];							inform_R[678][10] = r_cell_wire[333];							inform_R[167][10] = r_cell_wire[334];							inform_R[679][10] = r_cell_wire[335];							inform_R[168][10] = r_cell_wire[336];							inform_R[680][10] = r_cell_wire[337];							inform_R[169][10] = r_cell_wire[338];							inform_R[681][10] = r_cell_wire[339];							inform_R[170][10] = r_cell_wire[340];							inform_R[682][10] = r_cell_wire[341];							inform_R[171][10] = r_cell_wire[342];							inform_R[683][10] = r_cell_wire[343];							inform_R[172][10] = r_cell_wire[344];							inform_R[684][10] = r_cell_wire[345];							inform_R[173][10] = r_cell_wire[346];							inform_R[685][10] = r_cell_wire[347];							inform_R[174][10] = r_cell_wire[348];							inform_R[686][10] = r_cell_wire[349];							inform_R[175][10] = r_cell_wire[350];							inform_R[687][10] = r_cell_wire[351];							inform_R[176][10] = r_cell_wire[352];							inform_R[688][10] = r_cell_wire[353];							inform_R[177][10] = r_cell_wire[354];							inform_R[689][10] = r_cell_wire[355];							inform_R[178][10] = r_cell_wire[356];							inform_R[690][10] = r_cell_wire[357];							inform_R[179][10] = r_cell_wire[358];							inform_R[691][10] = r_cell_wire[359];							inform_R[180][10] = r_cell_wire[360];							inform_R[692][10] = r_cell_wire[361];							inform_R[181][10] = r_cell_wire[362];							inform_R[693][10] = r_cell_wire[363];							inform_R[182][10] = r_cell_wire[364];							inform_R[694][10] = r_cell_wire[365];							inform_R[183][10] = r_cell_wire[366];							inform_R[695][10] = r_cell_wire[367];							inform_R[184][10] = r_cell_wire[368];							inform_R[696][10] = r_cell_wire[369];							inform_R[185][10] = r_cell_wire[370];							inform_R[697][10] = r_cell_wire[371];							inform_R[186][10] = r_cell_wire[372];							inform_R[698][10] = r_cell_wire[373];							inform_R[187][10] = r_cell_wire[374];							inform_R[699][10] = r_cell_wire[375];							inform_R[188][10] = r_cell_wire[376];							inform_R[700][10] = r_cell_wire[377];							inform_R[189][10] = r_cell_wire[378];							inform_R[701][10] = r_cell_wire[379];							inform_R[190][10] = r_cell_wire[380];							inform_R[702][10] = r_cell_wire[381];							inform_R[191][10] = r_cell_wire[382];							inform_R[703][10] = r_cell_wire[383];							inform_R[192][10] = r_cell_wire[384];							inform_R[704][10] = r_cell_wire[385];							inform_R[193][10] = r_cell_wire[386];							inform_R[705][10] = r_cell_wire[387];							inform_R[194][10] = r_cell_wire[388];							inform_R[706][10] = r_cell_wire[389];							inform_R[195][10] = r_cell_wire[390];							inform_R[707][10] = r_cell_wire[391];							inform_R[196][10] = r_cell_wire[392];							inform_R[708][10] = r_cell_wire[393];							inform_R[197][10] = r_cell_wire[394];							inform_R[709][10] = r_cell_wire[395];							inform_R[198][10] = r_cell_wire[396];							inform_R[710][10] = r_cell_wire[397];							inform_R[199][10] = r_cell_wire[398];							inform_R[711][10] = r_cell_wire[399];							inform_R[200][10] = r_cell_wire[400];							inform_R[712][10] = r_cell_wire[401];							inform_R[201][10] = r_cell_wire[402];							inform_R[713][10] = r_cell_wire[403];							inform_R[202][10] = r_cell_wire[404];							inform_R[714][10] = r_cell_wire[405];							inform_R[203][10] = r_cell_wire[406];							inform_R[715][10] = r_cell_wire[407];							inform_R[204][10] = r_cell_wire[408];							inform_R[716][10] = r_cell_wire[409];							inform_R[205][10] = r_cell_wire[410];							inform_R[717][10] = r_cell_wire[411];							inform_R[206][10] = r_cell_wire[412];							inform_R[718][10] = r_cell_wire[413];							inform_R[207][10] = r_cell_wire[414];							inform_R[719][10] = r_cell_wire[415];							inform_R[208][10] = r_cell_wire[416];							inform_R[720][10] = r_cell_wire[417];							inform_R[209][10] = r_cell_wire[418];							inform_R[721][10] = r_cell_wire[419];							inform_R[210][10] = r_cell_wire[420];							inform_R[722][10] = r_cell_wire[421];							inform_R[211][10] = r_cell_wire[422];							inform_R[723][10] = r_cell_wire[423];							inform_R[212][10] = r_cell_wire[424];							inform_R[724][10] = r_cell_wire[425];							inform_R[213][10] = r_cell_wire[426];							inform_R[725][10] = r_cell_wire[427];							inform_R[214][10] = r_cell_wire[428];							inform_R[726][10] = r_cell_wire[429];							inform_R[215][10] = r_cell_wire[430];							inform_R[727][10] = r_cell_wire[431];							inform_R[216][10] = r_cell_wire[432];							inform_R[728][10] = r_cell_wire[433];							inform_R[217][10] = r_cell_wire[434];							inform_R[729][10] = r_cell_wire[435];							inform_R[218][10] = r_cell_wire[436];							inform_R[730][10] = r_cell_wire[437];							inform_R[219][10] = r_cell_wire[438];							inform_R[731][10] = r_cell_wire[439];							inform_R[220][10] = r_cell_wire[440];							inform_R[732][10] = r_cell_wire[441];							inform_R[221][10] = r_cell_wire[442];							inform_R[733][10] = r_cell_wire[443];							inform_R[222][10] = r_cell_wire[444];							inform_R[734][10] = r_cell_wire[445];							inform_R[223][10] = r_cell_wire[446];							inform_R[735][10] = r_cell_wire[447];							inform_R[224][10] = r_cell_wire[448];							inform_R[736][10] = r_cell_wire[449];							inform_R[225][10] = r_cell_wire[450];							inform_R[737][10] = r_cell_wire[451];							inform_R[226][10] = r_cell_wire[452];							inform_R[738][10] = r_cell_wire[453];							inform_R[227][10] = r_cell_wire[454];							inform_R[739][10] = r_cell_wire[455];							inform_R[228][10] = r_cell_wire[456];							inform_R[740][10] = r_cell_wire[457];							inform_R[229][10] = r_cell_wire[458];							inform_R[741][10] = r_cell_wire[459];							inform_R[230][10] = r_cell_wire[460];							inform_R[742][10] = r_cell_wire[461];							inform_R[231][10] = r_cell_wire[462];							inform_R[743][10] = r_cell_wire[463];							inform_R[232][10] = r_cell_wire[464];							inform_R[744][10] = r_cell_wire[465];							inform_R[233][10] = r_cell_wire[466];							inform_R[745][10] = r_cell_wire[467];							inform_R[234][10] = r_cell_wire[468];							inform_R[746][10] = r_cell_wire[469];							inform_R[235][10] = r_cell_wire[470];							inform_R[747][10] = r_cell_wire[471];							inform_R[236][10] = r_cell_wire[472];							inform_R[748][10] = r_cell_wire[473];							inform_R[237][10] = r_cell_wire[474];							inform_R[749][10] = r_cell_wire[475];							inform_R[238][10] = r_cell_wire[476];							inform_R[750][10] = r_cell_wire[477];							inform_R[239][10] = r_cell_wire[478];							inform_R[751][10] = r_cell_wire[479];							inform_R[240][10] = r_cell_wire[480];							inform_R[752][10] = r_cell_wire[481];							inform_R[241][10] = r_cell_wire[482];							inform_R[753][10] = r_cell_wire[483];							inform_R[242][10] = r_cell_wire[484];							inform_R[754][10] = r_cell_wire[485];							inform_R[243][10] = r_cell_wire[486];							inform_R[755][10] = r_cell_wire[487];							inform_R[244][10] = r_cell_wire[488];							inform_R[756][10] = r_cell_wire[489];							inform_R[245][10] = r_cell_wire[490];							inform_R[757][10] = r_cell_wire[491];							inform_R[246][10] = r_cell_wire[492];							inform_R[758][10] = r_cell_wire[493];							inform_R[247][10] = r_cell_wire[494];							inform_R[759][10] = r_cell_wire[495];							inform_R[248][10] = r_cell_wire[496];							inform_R[760][10] = r_cell_wire[497];							inform_R[249][10] = r_cell_wire[498];							inform_R[761][10] = r_cell_wire[499];							inform_R[250][10] = r_cell_wire[500];							inform_R[762][10] = r_cell_wire[501];							inform_R[251][10] = r_cell_wire[502];							inform_R[763][10] = r_cell_wire[503];							inform_R[252][10] = r_cell_wire[504];							inform_R[764][10] = r_cell_wire[505];							inform_R[253][10] = r_cell_wire[506];							inform_R[765][10] = r_cell_wire[507];							inform_R[254][10] = r_cell_wire[508];							inform_R[766][10] = r_cell_wire[509];							inform_R[255][10] = r_cell_wire[510];							inform_R[767][10] = r_cell_wire[511];							inform_R[256][10] = r_cell_wire[512];							inform_R[768][10] = r_cell_wire[513];							inform_R[257][10] = r_cell_wire[514];							inform_R[769][10] = r_cell_wire[515];							inform_R[258][10] = r_cell_wire[516];							inform_R[770][10] = r_cell_wire[517];							inform_R[259][10] = r_cell_wire[518];							inform_R[771][10] = r_cell_wire[519];							inform_R[260][10] = r_cell_wire[520];							inform_R[772][10] = r_cell_wire[521];							inform_R[261][10] = r_cell_wire[522];							inform_R[773][10] = r_cell_wire[523];							inform_R[262][10] = r_cell_wire[524];							inform_R[774][10] = r_cell_wire[525];							inform_R[263][10] = r_cell_wire[526];							inform_R[775][10] = r_cell_wire[527];							inform_R[264][10] = r_cell_wire[528];							inform_R[776][10] = r_cell_wire[529];							inform_R[265][10] = r_cell_wire[530];							inform_R[777][10] = r_cell_wire[531];							inform_R[266][10] = r_cell_wire[532];							inform_R[778][10] = r_cell_wire[533];							inform_R[267][10] = r_cell_wire[534];							inform_R[779][10] = r_cell_wire[535];							inform_R[268][10] = r_cell_wire[536];							inform_R[780][10] = r_cell_wire[537];							inform_R[269][10] = r_cell_wire[538];							inform_R[781][10] = r_cell_wire[539];							inform_R[270][10] = r_cell_wire[540];							inform_R[782][10] = r_cell_wire[541];							inform_R[271][10] = r_cell_wire[542];							inform_R[783][10] = r_cell_wire[543];							inform_R[272][10] = r_cell_wire[544];							inform_R[784][10] = r_cell_wire[545];							inform_R[273][10] = r_cell_wire[546];							inform_R[785][10] = r_cell_wire[547];							inform_R[274][10] = r_cell_wire[548];							inform_R[786][10] = r_cell_wire[549];							inform_R[275][10] = r_cell_wire[550];							inform_R[787][10] = r_cell_wire[551];							inform_R[276][10] = r_cell_wire[552];							inform_R[788][10] = r_cell_wire[553];							inform_R[277][10] = r_cell_wire[554];							inform_R[789][10] = r_cell_wire[555];							inform_R[278][10] = r_cell_wire[556];							inform_R[790][10] = r_cell_wire[557];							inform_R[279][10] = r_cell_wire[558];							inform_R[791][10] = r_cell_wire[559];							inform_R[280][10] = r_cell_wire[560];							inform_R[792][10] = r_cell_wire[561];							inform_R[281][10] = r_cell_wire[562];							inform_R[793][10] = r_cell_wire[563];							inform_R[282][10] = r_cell_wire[564];							inform_R[794][10] = r_cell_wire[565];							inform_R[283][10] = r_cell_wire[566];							inform_R[795][10] = r_cell_wire[567];							inform_R[284][10] = r_cell_wire[568];							inform_R[796][10] = r_cell_wire[569];							inform_R[285][10] = r_cell_wire[570];							inform_R[797][10] = r_cell_wire[571];							inform_R[286][10] = r_cell_wire[572];							inform_R[798][10] = r_cell_wire[573];							inform_R[287][10] = r_cell_wire[574];							inform_R[799][10] = r_cell_wire[575];							inform_R[288][10] = r_cell_wire[576];							inform_R[800][10] = r_cell_wire[577];							inform_R[289][10] = r_cell_wire[578];							inform_R[801][10] = r_cell_wire[579];							inform_R[290][10] = r_cell_wire[580];							inform_R[802][10] = r_cell_wire[581];							inform_R[291][10] = r_cell_wire[582];							inform_R[803][10] = r_cell_wire[583];							inform_R[292][10] = r_cell_wire[584];							inform_R[804][10] = r_cell_wire[585];							inform_R[293][10] = r_cell_wire[586];							inform_R[805][10] = r_cell_wire[587];							inform_R[294][10] = r_cell_wire[588];							inform_R[806][10] = r_cell_wire[589];							inform_R[295][10] = r_cell_wire[590];							inform_R[807][10] = r_cell_wire[591];							inform_R[296][10] = r_cell_wire[592];							inform_R[808][10] = r_cell_wire[593];							inform_R[297][10] = r_cell_wire[594];							inform_R[809][10] = r_cell_wire[595];							inform_R[298][10] = r_cell_wire[596];							inform_R[810][10] = r_cell_wire[597];							inform_R[299][10] = r_cell_wire[598];							inform_R[811][10] = r_cell_wire[599];							inform_R[300][10] = r_cell_wire[600];							inform_R[812][10] = r_cell_wire[601];							inform_R[301][10] = r_cell_wire[602];							inform_R[813][10] = r_cell_wire[603];							inform_R[302][10] = r_cell_wire[604];							inform_R[814][10] = r_cell_wire[605];							inform_R[303][10] = r_cell_wire[606];							inform_R[815][10] = r_cell_wire[607];							inform_R[304][10] = r_cell_wire[608];							inform_R[816][10] = r_cell_wire[609];							inform_R[305][10] = r_cell_wire[610];							inform_R[817][10] = r_cell_wire[611];							inform_R[306][10] = r_cell_wire[612];							inform_R[818][10] = r_cell_wire[613];							inform_R[307][10] = r_cell_wire[614];							inform_R[819][10] = r_cell_wire[615];							inform_R[308][10] = r_cell_wire[616];							inform_R[820][10] = r_cell_wire[617];							inform_R[309][10] = r_cell_wire[618];							inform_R[821][10] = r_cell_wire[619];							inform_R[310][10] = r_cell_wire[620];							inform_R[822][10] = r_cell_wire[621];							inform_R[311][10] = r_cell_wire[622];							inform_R[823][10] = r_cell_wire[623];							inform_R[312][10] = r_cell_wire[624];							inform_R[824][10] = r_cell_wire[625];							inform_R[313][10] = r_cell_wire[626];							inform_R[825][10] = r_cell_wire[627];							inform_R[314][10] = r_cell_wire[628];							inform_R[826][10] = r_cell_wire[629];							inform_R[315][10] = r_cell_wire[630];							inform_R[827][10] = r_cell_wire[631];							inform_R[316][10] = r_cell_wire[632];							inform_R[828][10] = r_cell_wire[633];							inform_R[317][10] = r_cell_wire[634];							inform_R[829][10] = r_cell_wire[635];							inform_R[318][10] = r_cell_wire[636];							inform_R[830][10] = r_cell_wire[637];							inform_R[319][10] = r_cell_wire[638];							inform_R[831][10] = r_cell_wire[639];							inform_R[320][10] = r_cell_wire[640];							inform_R[832][10] = r_cell_wire[641];							inform_R[321][10] = r_cell_wire[642];							inform_R[833][10] = r_cell_wire[643];							inform_R[322][10] = r_cell_wire[644];							inform_R[834][10] = r_cell_wire[645];							inform_R[323][10] = r_cell_wire[646];							inform_R[835][10] = r_cell_wire[647];							inform_R[324][10] = r_cell_wire[648];							inform_R[836][10] = r_cell_wire[649];							inform_R[325][10] = r_cell_wire[650];							inform_R[837][10] = r_cell_wire[651];							inform_R[326][10] = r_cell_wire[652];							inform_R[838][10] = r_cell_wire[653];							inform_R[327][10] = r_cell_wire[654];							inform_R[839][10] = r_cell_wire[655];							inform_R[328][10] = r_cell_wire[656];							inform_R[840][10] = r_cell_wire[657];							inform_R[329][10] = r_cell_wire[658];							inform_R[841][10] = r_cell_wire[659];							inform_R[330][10] = r_cell_wire[660];							inform_R[842][10] = r_cell_wire[661];							inform_R[331][10] = r_cell_wire[662];							inform_R[843][10] = r_cell_wire[663];							inform_R[332][10] = r_cell_wire[664];							inform_R[844][10] = r_cell_wire[665];							inform_R[333][10] = r_cell_wire[666];							inform_R[845][10] = r_cell_wire[667];							inform_R[334][10] = r_cell_wire[668];							inform_R[846][10] = r_cell_wire[669];							inform_R[335][10] = r_cell_wire[670];							inform_R[847][10] = r_cell_wire[671];							inform_R[336][10] = r_cell_wire[672];							inform_R[848][10] = r_cell_wire[673];							inform_R[337][10] = r_cell_wire[674];							inform_R[849][10] = r_cell_wire[675];							inform_R[338][10] = r_cell_wire[676];							inform_R[850][10] = r_cell_wire[677];							inform_R[339][10] = r_cell_wire[678];							inform_R[851][10] = r_cell_wire[679];							inform_R[340][10] = r_cell_wire[680];							inform_R[852][10] = r_cell_wire[681];							inform_R[341][10] = r_cell_wire[682];							inform_R[853][10] = r_cell_wire[683];							inform_R[342][10] = r_cell_wire[684];							inform_R[854][10] = r_cell_wire[685];							inform_R[343][10] = r_cell_wire[686];							inform_R[855][10] = r_cell_wire[687];							inform_R[344][10] = r_cell_wire[688];							inform_R[856][10] = r_cell_wire[689];							inform_R[345][10] = r_cell_wire[690];							inform_R[857][10] = r_cell_wire[691];							inform_R[346][10] = r_cell_wire[692];							inform_R[858][10] = r_cell_wire[693];							inform_R[347][10] = r_cell_wire[694];							inform_R[859][10] = r_cell_wire[695];							inform_R[348][10] = r_cell_wire[696];							inform_R[860][10] = r_cell_wire[697];							inform_R[349][10] = r_cell_wire[698];							inform_R[861][10] = r_cell_wire[699];							inform_R[350][10] = r_cell_wire[700];							inform_R[862][10] = r_cell_wire[701];							inform_R[351][10] = r_cell_wire[702];							inform_R[863][10] = r_cell_wire[703];							inform_R[352][10] = r_cell_wire[704];							inform_R[864][10] = r_cell_wire[705];							inform_R[353][10] = r_cell_wire[706];							inform_R[865][10] = r_cell_wire[707];							inform_R[354][10] = r_cell_wire[708];							inform_R[866][10] = r_cell_wire[709];							inform_R[355][10] = r_cell_wire[710];							inform_R[867][10] = r_cell_wire[711];							inform_R[356][10] = r_cell_wire[712];							inform_R[868][10] = r_cell_wire[713];							inform_R[357][10] = r_cell_wire[714];							inform_R[869][10] = r_cell_wire[715];							inform_R[358][10] = r_cell_wire[716];							inform_R[870][10] = r_cell_wire[717];							inform_R[359][10] = r_cell_wire[718];							inform_R[871][10] = r_cell_wire[719];							inform_R[360][10] = r_cell_wire[720];							inform_R[872][10] = r_cell_wire[721];							inform_R[361][10] = r_cell_wire[722];							inform_R[873][10] = r_cell_wire[723];							inform_R[362][10] = r_cell_wire[724];							inform_R[874][10] = r_cell_wire[725];							inform_R[363][10] = r_cell_wire[726];							inform_R[875][10] = r_cell_wire[727];							inform_R[364][10] = r_cell_wire[728];							inform_R[876][10] = r_cell_wire[729];							inform_R[365][10] = r_cell_wire[730];							inform_R[877][10] = r_cell_wire[731];							inform_R[366][10] = r_cell_wire[732];							inform_R[878][10] = r_cell_wire[733];							inform_R[367][10] = r_cell_wire[734];							inform_R[879][10] = r_cell_wire[735];							inform_R[368][10] = r_cell_wire[736];							inform_R[880][10] = r_cell_wire[737];							inform_R[369][10] = r_cell_wire[738];							inform_R[881][10] = r_cell_wire[739];							inform_R[370][10] = r_cell_wire[740];							inform_R[882][10] = r_cell_wire[741];							inform_R[371][10] = r_cell_wire[742];							inform_R[883][10] = r_cell_wire[743];							inform_R[372][10] = r_cell_wire[744];							inform_R[884][10] = r_cell_wire[745];							inform_R[373][10] = r_cell_wire[746];							inform_R[885][10] = r_cell_wire[747];							inform_R[374][10] = r_cell_wire[748];							inform_R[886][10] = r_cell_wire[749];							inform_R[375][10] = r_cell_wire[750];							inform_R[887][10] = r_cell_wire[751];							inform_R[376][10] = r_cell_wire[752];							inform_R[888][10] = r_cell_wire[753];							inform_R[377][10] = r_cell_wire[754];							inform_R[889][10] = r_cell_wire[755];							inform_R[378][10] = r_cell_wire[756];							inform_R[890][10] = r_cell_wire[757];							inform_R[379][10] = r_cell_wire[758];							inform_R[891][10] = r_cell_wire[759];							inform_R[380][10] = r_cell_wire[760];							inform_R[892][10] = r_cell_wire[761];							inform_R[381][10] = r_cell_wire[762];							inform_R[893][10] = r_cell_wire[763];							inform_R[382][10] = r_cell_wire[764];							inform_R[894][10] = r_cell_wire[765];							inform_R[383][10] = r_cell_wire[766];							inform_R[895][10] = r_cell_wire[767];							inform_R[384][10] = r_cell_wire[768];							inform_R[896][10] = r_cell_wire[769];							inform_R[385][10] = r_cell_wire[770];							inform_R[897][10] = r_cell_wire[771];							inform_R[386][10] = r_cell_wire[772];							inform_R[898][10] = r_cell_wire[773];							inform_R[387][10] = r_cell_wire[774];							inform_R[899][10] = r_cell_wire[775];							inform_R[388][10] = r_cell_wire[776];							inform_R[900][10] = r_cell_wire[777];							inform_R[389][10] = r_cell_wire[778];							inform_R[901][10] = r_cell_wire[779];							inform_R[390][10] = r_cell_wire[780];							inform_R[902][10] = r_cell_wire[781];							inform_R[391][10] = r_cell_wire[782];							inform_R[903][10] = r_cell_wire[783];							inform_R[392][10] = r_cell_wire[784];							inform_R[904][10] = r_cell_wire[785];							inform_R[393][10] = r_cell_wire[786];							inform_R[905][10] = r_cell_wire[787];							inform_R[394][10] = r_cell_wire[788];							inform_R[906][10] = r_cell_wire[789];							inform_R[395][10] = r_cell_wire[790];							inform_R[907][10] = r_cell_wire[791];							inform_R[396][10] = r_cell_wire[792];							inform_R[908][10] = r_cell_wire[793];							inform_R[397][10] = r_cell_wire[794];							inform_R[909][10] = r_cell_wire[795];							inform_R[398][10] = r_cell_wire[796];							inform_R[910][10] = r_cell_wire[797];							inform_R[399][10] = r_cell_wire[798];							inform_R[911][10] = r_cell_wire[799];							inform_R[400][10] = r_cell_wire[800];							inform_R[912][10] = r_cell_wire[801];							inform_R[401][10] = r_cell_wire[802];							inform_R[913][10] = r_cell_wire[803];							inform_R[402][10] = r_cell_wire[804];							inform_R[914][10] = r_cell_wire[805];							inform_R[403][10] = r_cell_wire[806];							inform_R[915][10] = r_cell_wire[807];							inform_R[404][10] = r_cell_wire[808];							inform_R[916][10] = r_cell_wire[809];							inform_R[405][10] = r_cell_wire[810];							inform_R[917][10] = r_cell_wire[811];							inform_R[406][10] = r_cell_wire[812];							inform_R[918][10] = r_cell_wire[813];							inform_R[407][10] = r_cell_wire[814];							inform_R[919][10] = r_cell_wire[815];							inform_R[408][10] = r_cell_wire[816];							inform_R[920][10] = r_cell_wire[817];							inform_R[409][10] = r_cell_wire[818];							inform_R[921][10] = r_cell_wire[819];							inform_R[410][10] = r_cell_wire[820];							inform_R[922][10] = r_cell_wire[821];							inform_R[411][10] = r_cell_wire[822];							inform_R[923][10] = r_cell_wire[823];							inform_R[412][10] = r_cell_wire[824];							inform_R[924][10] = r_cell_wire[825];							inform_R[413][10] = r_cell_wire[826];							inform_R[925][10] = r_cell_wire[827];							inform_R[414][10] = r_cell_wire[828];							inform_R[926][10] = r_cell_wire[829];							inform_R[415][10] = r_cell_wire[830];							inform_R[927][10] = r_cell_wire[831];							inform_R[416][10] = r_cell_wire[832];							inform_R[928][10] = r_cell_wire[833];							inform_R[417][10] = r_cell_wire[834];							inform_R[929][10] = r_cell_wire[835];							inform_R[418][10] = r_cell_wire[836];							inform_R[930][10] = r_cell_wire[837];							inform_R[419][10] = r_cell_wire[838];							inform_R[931][10] = r_cell_wire[839];							inform_R[420][10] = r_cell_wire[840];							inform_R[932][10] = r_cell_wire[841];							inform_R[421][10] = r_cell_wire[842];							inform_R[933][10] = r_cell_wire[843];							inform_R[422][10] = r_cell_wire[844];							inform_R[934][10] = r_cell_wire[845];							inform_R[423][10] = r_cell_wire[846];							inform_R[935][10] = r_cell_wire[847];							inform_R[424][10] = r_cell_wire[848];							inform_R[936][10] = r_cell_wire[849];							inform_R[425][10] = r_cell_wire[850];							inform_R[937][10] = r_cell_wire[851];							inform_R[426][10] = r_cell_wire[852];							inform_R[938][10] = r_cell_wire[853];							inform_R[427][10] = r_cell_wire[854];							inform_R[939][10] = r_cell_wire[855];							inform_R[428][10] = r_cell_wire[856];							inform_R[940][10] = r_cell_wire[857];							inform_R[429][10] = r_cell_wire[858];							inform_R[941][10] = r_cell_wire[859];							inform_R[430][10] = r_cell_wire[860];							inform_R[942][10] = r_cell_wire[861];							inform_R[431][10] = r_cell_wire[862];							inform_R[943][10] = r_cell_wire[863];							inform_R[432][10] = r_cell_wire[864];							inform_R[944][10] = r_cell_wire[865];							inform_R[433][10] = r_cell_wire[866];							inform_R[945][10] = r_cell_wire[867];							inform_R[434][10] = r_cell_wire[868];							inform_R[946][10] = r_cell_wire[869];							inform_R[435][10] = r_cell_wire[870];							inform_R[947][10] = r_cell_wire[871];							inform_R[436][10] = r_cell_wire[872];							inform_R[948][10] = r_cell_wire[873];							inform_R[437][10] = r_cell_wire[874];							inform_R[949][10] = r_cell_wire[875];							inform_R[438][10] = r_cell_wire[876];							inform_R[950][10] = r_cell_wire[877];							inform_R[439][10] = r_cell_wire[878];							inform_R[951][10] = r_cell_wire[879];							inform_R[440][10] = r_cell_wire[880];							inform_R[952][10] = r_cell_wire[881];							inform_R[441][10] = r_cell_wire[882];							inform_R[953][10] = r_cell_wire[883];							inform_R[442][10] = r_cell_wire[884];							inform_R[954][10] = r_cell_wire[885];							inform_R[443][10] = r_cell_wire[886];							inform_R[955][10] = r_cell_wire[887];							inform_R[444][10] = r_cell_wire[888];							inform_R[956][10] = r_cell_wire[889];							inform_R[445][10] = r_cell_wire[890];							inform_R[957][10] = r_cell_wire[891];							inform_R[446][10] = r_cell_wire[892];							inform_R[958][10] = r_cell_wire[893];							inform_R[447][10] = r_cell_wire[894];							inform_R[959][10] = r_cell_wire[895];							inform_R[448][10] = r_cell_wire[896];							inform_R[960][10] = r_cell_wire[897];							inform_R[449][10] = r_cell_wire[898];							inform_R[961][10] = r_cell_wire[899];							inform_R[450][10] = r_cell_wire[900];							inform_R[962][10] = r_cell_wire[901];							inform_R[451][10] = r_cell_wire[902];							inform_R[963][10] = r_cell_wire[903];							inform_R[452][10] = r_cell_wire[904];							inform_R[964][10] = r_cell_wire[905];							inform_R[453][10] = r_cell_wire[906];							inform_R[965][10] = r_cell_wire[907];							inform_R[454][10] = r_cell_wire[908];							inform_R[966][10] = r_cell_wire[909];							inform_R[455][10] = r_cell_wire[910];							inform_R[967][10] = r_cell_wire[911];							inform_R[456][10] = r_cell_wire[912];							inform_R[968][10] = r_cell_wire[913];							inform_R[457][10] = r_cell_wire[914];							inform_R[969][10] = r_cell_wire[915];							inform_R[458][10] = r_cell_wire[916];							inform_R[970][10] = r_cell_wire[917];							inform_R[459][10] = r_cell_wire[918];							inform_R[971][10] = r_cell_wire[919];							inform_R[460][10] = r_cell_wire[920];							inform_R[972][10] = r_cell_wire[921];							inform_R[461][10] = r_cell_wire[922];							inform_R[973][10] = r_cell_wire[923];							inform_R[462][10] = r_cell_wire[924];							inform_R[974][10] = r_cell_wire[925];							inform_R[463][10] = r_cell_wire[926];							inform_R[975][10] = r_cell_wire[927];							inform_R[464][10] = r_cell_wire[928];							inform_R[976][10] = r_cell_wire[929];							inform_R[465][10] = r_cell_wire[930];							inform_R[977][10] = r_cell_wire[931];							inform_R[466][10] = r_cell_wire[932];							inform_R[978][10] = r_cell_wire[933];							inform_R[467][10] = r_cell_wire[934];							inform_R[979][10] = r_cell_wire[935];							inform_R[468][10] = r_cell_wire[936];							inform_R[980][10] = r_cell_wire[937];							inform_R[469][10] = r_cell_wire[938];							inform_R[981][10] = r_cell_wire[939];							inform_R[470][10] = r_cell_wire[940];							inform_R[982][10] = r_cell_wire[941];							inform_R[471][10] = r_cell_wire[942];							inform_R[983][10] = r_cell_wire[943];							inform_R[472][10] = r_cell_wire[944];							inform_R[984][10] = r_cell_wire[945];							inform_R[473][10] = r_cell_wire[946];							inform_R[985][10] = r_cell_wire[947];							inform_R[474][10] = r_cell_wire[948];							inform_R[986][10] = r_cell_wire[949];							inform_R[475][10] = r_cell_wire[950];							inform_R[987][10] = r_cell_wire[951];							inform_R[476][10] = r_cell_wire[952];							inform_R[988][10] = r_cell_wire[953];							inform_R[477][10] = r_cell_wire[954];							inform_R[989][10] = r_cell_wire[955];							inform_R[478][10] = r_cell_wire[956];							inform_R[990][10] = r_cell_wire[957];							inform_R[479][10] = r_cell_wire[958];							inform_R[991][10] = r_cell_wire[959];							inform_R[480][10] = r_cell_wire[960];							inform_R[992][10] = r_cell_wire[961];							inform_R[481][10] = r_cell_wire[962];							inform_R[993][10] = r_cell_wire[963];							inform_R[482][10] = r_cell_wire[964];							inform_R[994][10] = r_cell_wire[965];							inform_R[483][10] = r_cell_wire[966];							inform_R[995][10] = r_cell_wire[967];							inform_R[484][10] = r_cell_wire[968];							inform_R[996][10] = r_cell_wire[969];							inform_R[485][10] = r_cell_wire[970];							inform_R[997][10] = r_cell_wire[971];							inform_R[486][10] = r_cell_wire[972];							inform_R[998][10] = r_cell_wire[973];							inform_R[487][10] = r_cell_wire[974];							inform_R[999][10] = r_cell_wire[975];							inform_R[488][10] = r_cell_wire[976];							inform_R[1000][10] = r_cell_wire[977];							inform_R[489][10] = r_cell_wire[978];							inform_R[1001][10] = r_cell_wire[979];							inform_R[490][10] = r_cell_wire[980];							inform_R[1002][10] = r_cell_wire[981];							inform_R[491][10] = r_cell_wire[982];							inform_R[1003][10] = r_cell_wire[983];							inform_R[492][10] = r_cell_wire[984];							inform_R[1004][10] = r_cell_wire[985];							inform_R[493][10] = r_cell_wire[986];							inform_R[1005][10] = r_cell_wire[987];							inform_R[494][10] = r_cell_wire[988];							inform_R[1006][10] = r_cell_wire[989];							inform_R[495][10] = r_cell_wire[990];							inform_R[1007][10] = r_cell_wire[991];							inform_R[496][10] = r_cell_wire[992];							inform_R[1008][10] = r_cell_wire[993];							inform_R[497][10] = r_cell_wire[994];							inform_R[1009][10] = r_cell_wire[995];							inform_R[498][10] = r_cell_wire[996];							inform_R[1010][10] = r_cell_wire[997];							inform_R[499][10] = r_cell_wire[998];							inform_R[1011][10] = r_cell_wire[999];							inform_R[500][10] = r_cell_wire[1000];							inform_R[1012][10] = r_cell_wire[1001];							inform_R[501][10] = r_cell_wire[1002];							inform_R[1013][10] = r_cell_wire[1003];							inform_R[502][10] = r_cell_wire[1004];							inform_R[1014][10] = r_cell_wire[1005];							inform_R[503][10] = r_cell_wire[1006];							inform_R[1015][10] = r_cell_wire[1007];							inform_R[504][10] = r_cell_wire[1008];							inform_R[1016][10] = r_cell_wire[1009];							inform_R[505][10] = r_cell_wire[1010];							inform_R[1017][10] = r_cell_wire[1011];							inform_R[506][10] = r_cell_wire[1012];							inform_R[1018][10] = r_cell_wire[1013];							inform_R[507][10] = r_cell_wire[1014];							inform_R[1019][10] = r_cell_wire[1015];							inform_R[508][10] = r_cell_wire[1016];							inform_R[1020][10] = r_cell_wire[1017];							inform_R[509][10] = r_cell_wire[1018];							inform_R[1021][10] = r_cell_wire[1019];							inform_R[510][10] = r_cell_wire[1020];							inform_R[1022][10] = r_cell_wire[1021];							inform_R[511][10] = r_cell_wire[1022];							inform_R[1023][10] = r_cell_wire[1023];							inform_L[0][9] = l_cell_wire[0];							inform_L[512][9] = l_cell_wire[1];							inform_L[1][9] = l_cell_wire[2];							inform_L[513][9] = l_cell_wire[3];							inform_L[2][9] = l_cell_wire[4];							inform_L[514][9] = l_cell_wire[5];							inform_L[3][9] = l_cell_wire[6];							inform_L[515][9] = l_cell_wire[7];							inform_L[4][9] = l_cell_wire[8];							inform_L[516][9] = l_cell_wire[9];							inform_L[5][9] = l_cell_wire[10];							inform_L[517][9] = l_cell_wire[11];							inform_L[6][9] = l_cell_wire[12];							inform_L[518][9] = l_cell_wire[13];							inform_L[7][9] = l_cell_wire[14];							inform_L[519][9] = l_cell_wire[15];							inform_L[8][9] = l_cell_wire[16];							inform_L[520][9] = l_cell_wire[17];							inform_L[9][9] = l_cell_wire[18];							inform_L[521][9] = l_cell_wire[19];							inform_L[10][9] = l_cell_wire[20];							inform_L[522][9] = l_cell_wire[21];							inform_L[11][9] = l_cell_wire[22];							inform_L[523][9] = l_cell_wire[23];							inform_L[12][9] = l_cell_wire[24];							inform_L[524][9] = l_cell_wire[25];							inform_L[13][9] = l_cell_wire[26];							inform_L[525][9] = l_cell_wire[27];							inform_L[14][9] = l_cell_wire[28];							inform_L[526][9] = l_cell_wire[29];							inform_L[15][9] = l_cell_wire[30];							inform_L[527][9] = l_cell_wire[31];							inform_L[16][9] = l_cell_wire[32];							inform_L[528][9] = l_cell_wire[33];							inform_L[17][9] = l_cell_wire[34];							inform_L[529][9] = l_cell_wire[35];							inform_L[18][9] = l_cell_wire[36];							inform_L[530][9] = l_cell_wire[37];							inform_L[19][9] = l_cell_wire[38];							inform_L[531][9] = l_cell_wire[39];							inform_L[20][9] = l_cell_wire[40];							inform_L[532][9] = l_cell_wire[41];							inform_L[21][9] = l_cell_wire[42];							inform_L[533][9] = l_cell_wire[43];							inform_L[22][9] = l_cell_wire[44];							inform_L[534][9] = l_cell_wire[45];							inform_L[23][9] = l_cell_wire[46];							inform_L[535][9] = l_cell_wire[47];							inform_L[24][9] = l_cell_wire[48];							inform_L[536][9] = l_cell_wire[49];							inform_L[25][9] = l_cell_wire[50];							inform_L[537][9] = l_cell_wire[51];							inform_L[26][9] = l_cell_wire[52];							inform_L[538][9] = l_cell_wire[53];							inform_L[27][9] = l_cell_wire[54];							inform_L[539][9] = l_cell_wire[55];							inform_L[28][9] = l_cell_wire[56];							inform_L[540][9] = l_cell_wire[57];							inform_L[29][9] = l_cell_wire[58];							inform_L[541][9] = l_cell_wire[59];							inform_L[30][9] = l_cell_wire[60];							inform_L[542][9] = l_cell_wire[61];							inform_L[31][9] = l_cell_wire[62];							inform_L[543][9] = l_cell_wire[63];							inform_L[32][9] = l_cell_wire[64];							inform_L[544][9] = l_cell_wire[65];							inform_L[33][9] = l_cell_wire[66];							inform_L[545][9] = l_cell_wire[67];							inform_L[34][9] = l_cell_wire[68];							inform_L[546][9] = l_cell_wire[69];							inform_L[35][9] = l_cell_wire[70];							inform_L[547][9] = l_cell_wire[71];							inform_L[36][9] = l_cell_wire[72];							inform_L[548][9] = l_cell_wire[73];							inform_L[37][9] = l_cell_wire[74];							inform_L[549][9] = l_cell_wire[75];							inform_L[38][9] = l_cell_wire[76];							inform_L[550][9] = l_cell_wire[77];							inform_L[39][9] = l_cell_wire[78];							inform_L[551][9] = l_cell_wire[79];							inform_L[40][9] = l_cell_wire[80];							inform_L[552][9] = l_cell_wire[81];							inform_L[41][9] = l_cell_wire[82];							inform_L[553][9] = l_cell_wire[83];							inform_L[42][9] = l_cell_wire[84];							inform_L[554][9] = l_cell_wire[85];							inform_L[43][9] = l_cell_wire[86];							inform_L[555][9] = l_cell_wire[87];							inform_L[44][9] = l_cell_wire[88];							inform_L[556][9] = l_cell_wire[89];							inform_L[45][9] = l_cell_wire[90];							inform_L[557][9] = l_cell_wire[91];							inform_L[46][9] = l_cell_wire[92];							inform_L[558][9] = l_cell_wire[93];							inform_L[47][9] = l_cell_wire[94];							inform_L[559][9] = l_cell_wire[95];							inform_L[48][9] = l_cell_wire[96];							inform_L[560][9] = l_cell_wire[97];							inform_L[49][9] = l_cell_wire[98];							inform_L[561][9] = l_cell_wire[99];							inform_L[50][9] = l_cell_wire[100];							inform_L[562][9] = l_cell_wire[101];							inform_L[51][9] = l_cell_wire[102];							inform_L[563][9] = l_cell_wire[103];							inform_L[52][9] = l_cell_wire[104];							inform_L[564][9] = l_cell_wire[105];							inform_L[53][9] = l_cell_wire[106];							inform_L[565][9] = l_cell_wire[107];							inform_L[54][9] = l_cell_wire[108];							inform_L[566][9] = l_cell_wire[109];							inform_L[55][9] = l_cell_wire[110];							inform_L[567][9] = l_cell_wire[111];							inform_L[56][9] = l_cell_wire[112];							inform_L[568][9] = l_cell_wire[113];							inform_L[57][9] = l_cell_wire[114];							inform_L[569][9] = l_cell_wire[115];							inform_L[58][9] = l_cell_wire[116];							inform_L[570][9] = l_cell_wire[117];							inform_L[59][9] = l_cell_wire[118];							inform_L[571][9] = l_cell_wire[119];							inform_L[60][9] = l_cell_wire[120];							inform_L[572][9] = l_cell_wire[121];							inform_L[61][9] = l_cell_wire[122];							inform_L[573][9] = l_cell_wire[123];							inform_L[62][9] = l_cell_wire[124];							inform_L[574][9] = l_cell_wire[125];							inform_L[63][9] = l_cell_wire[126];							inform_L[575][9] = l_cell_wire[127];							inform_L[64][9] = l_cell_wire[128];							inform_L[576][9] = l_cell_wire[129];							inform_L[65][9] = l_cell_wire[130];							inform_L[577][9] = l_cell_wire[131];							inform_L[66][9] = l_cell_wire[132];							inform_L[578][9] = l_cell_wire[133];							inform_L[67][9] = l_cell_wire[134];							inform_L[579][9] = l_cell_wire[135];							inform_L[68][9] = l_cell_wire[136];							inform_L[580][9] = l_cell_wire[137];							inform_L[69][9] = l_cell_wire[138];							inform_L[581][9] = l_cell_wire[139];							inform_L[70][9] = l_cell_wire[140];							inform_L[582][9] = l_cell_wire[141];							inform_L[71][9] = l_cell_wire[142];							inform_L[583][9] = l_cell_wire[143];							inform_L[72][9] = l_cell_wire[144];							inform_L[584][9] = l_cell_wire[145];							inform_L[73][9] = l_cell_wire[146];							inform_L[585][9] = l_cell_wire[147];							inform_L[74][9] = l_cell_wire[148];							inform_L[586][9] = l_cell_wire[149];							inform_L[75][9] = l_cell_wire[150];							inform_L[587][9] = l_cell_wire[151];							inform_L[76][9] = l_cell_wire[152];							inform_L[588][9] = l_cell_wire[153];							inform_L[77][9] = l_cell_wire[154];							inform_L[589][9] = l_cell_wire[155];							inform_L[78][9] = l_cell_wire[156];							inform_L[590][9] = l_cell_wire[157];							inform_L[79][9] = l_cell_wire[158];							inform_L[591][9] = l_cell_wire[159];							inform_L[80][9] = l_cell_wire[160];							inform_L[592][9] = l_cell_wire[161];							inform_L[81][9] = l_cell_wire[162];							inform_L[593][9] = l_cell_wire[163];							inform_L[82][9] = l_cell_wire[164];							inform_L[594][9] = l_cell_wire[165];							inform_L[83][9] = l_cell_wire[166];							inform_L[595][9] = l_cell_wire[167];							inform_L[84][9] = l_cell_wire[168];							inform_L[596][9] = l_cell_wire[169];							inform_L[85][9] = l_cell_wire[170];							inform_L[597][9] = l_cell_wire[171];							inform_L[86][9] = l_cell_wire[172];							inform_L[598][9] = l_cell_wire[173];							inform_L[87][9] = l_cell_wire[174];							inform_L[599][9] = l_cell_wire[175];							inform_L[88][9] = l_cell_wire[176];							inform_L[600][9] = l_cell_wire[177];							inform_L[89][9] = l_cell_wire[178];							inform_L[601][9] = l_cell_wire[179];							inform_L[90][9] = l_cell_wire[180];							inform_L[602][9] = l_cell_wire[181];							inform_L[91][9] = l_cell_wire[182];							inform_L[603][9] = l_cell_wire[183];							inform_L[92][9] = l_cell_wire[184];							inform_L[604][9] = l_cell_wire[185];							inform_L[93][9] = l_cell_wire[186];							inform_L[605][9] = l_cell_wire[187];							inform_L[94][9] = l_cell_wire[188];							inform_L[606][9] = l_cell_wire[189];							inform_L[95][9] = l_cell_wire[190];							inform_L[607][9] = l_cell_wire[191];							inform_L[96][9] = l_cell_wire[192];							inform_L[608][9] = l_cell_wire[193];							inform_L[97][9] = l_cell_wire[194];							inform_L[609][9] = l_cell_wire[195];							inform_L[98][9] = l_cell_wire[196];							inform_L[610][9] = l_cell_wire[197];							inform_L[99][9] = l_cell_wire[198];							inform_L[611][9] = l_cell_wire[199];							inform_L[100][9] = l_cell_wire[200];							inform_L[612][9] = l_cell_wire[201];							inform_L[101][9] = l_cell_wire[202];							inform_L[613][9] = l_cell_wire[203];							inform_L[102][9] = l_cell_wire[204];							inform_L[614][9] = l_cell_wire[205];							inform_L[103][9] = l_cell_wire[206];							inform_L[615][9] = l_cell_wire[207];							inform_L[104][9] = l_cell_wire[208];							inform_L[616][9] = l_cell_wire[209];							inform_L[105][9] = l_cell_wire[210];							inform_L[617][9] = l_cell_wire[211];							inform_L[106][9] = l_cell_wire[212];							inform_L[618][9] = l_cell_wire[213];							inform_L[107][9] = l_cell_wire[214];							inform_L[619][9] = l_cell_wire[215];							inform_L[108][9] = l_cell_wire[216];							inform_L[620][9] = l_cell_wire[217];							inform_L[109][9] = l_cell_wire[218];							inform_L[621][9] = l_cell_wire[219];							inform_L[110][9] = l_cell_wire[220];							inform_L[622][9] = l_cell_wire[221];							inform_L[111][9] = l_cell_wire[222];							inform_L[623][9] = l_cell_wire[223];							inform_L[112][9] = l_cell_wire[224];							inform_L[624][9] = l_cell_wire[225];							inform_L[113][9] = l_cell_wire[226];							inform_L[625][9] = l_cell_wire[227];							inform_L[114][9] = l_cell_wire[228];							inform_L[626][9] = l_cell_wire[229];							inform_L[115][9] = l_cell_wire[230];							inform_L[627][9] = l_cell_wire[231];							inform_L[116][9] = l_cell_wire[232];							inform_L[628][9] = l_cell_wire[233];							inform_L[117][9] = l_cell_wire[234];							inform_L[629][9] = l_cell_wire[235];							inform_L[118][9] = l_cell_wire[236];							inform_L[630][9] = l_cell_wire[237];							inform_L[119][9] = l_cell_wire[238];							inform_L[631][9] = l_cell_wire[239];							inform_L[120][9] = l_cell_wire[240];							inform_L[632][9] = l_cell_wire[241];							inform_L[121][9] = l_cell_wire[242];							inform_L[633][9] = l_cell_wire[243];							inform_L[122][9] = l_cell_wire[244];							inform_L[634][9] = l_cell_wire[245];							inform_L[123][9] = l_cell_wire[246];							inform_L[635][9] = l_cell_wire[247];							inform_L[124][9] = l_cell_wire[248];							inform_L[636][9] = l_cell_wire[249];							inform_L[125][9] = l_cell_wire[250];							inform_L[637][9] = l_cell_wire[251];							inform_L[126][9] = l_cell_wire[252];							inform_L[638][9] = l_cell_wire[253];							inform_L[127][9] = l_cell_wire[254];							inform_L[639][9] = l_cell_wire[255];							inform_L[128][9] = l_cell_wire[256];							inform_L[640][9] = l_cell_wire[257];							inform_L[129][9] = l_cell_wire[258];							inform_L[641][9] = l_cell_wire[259];							inform_L[130][9] = l_cell_wire[260];							inform_L[642][9] = l_cell_wire[261];							inform_L[131][9] = l_cell_wire[262];							inform_L[643][9] = l_cell_wire[263];							inform_L[132][9] = l_cell_wire[264];							inform_L[644][9] = l_cell_wire[265];							inform_L[133][9] = l_cell_wire[266];							inform_L[645][9] = l_cell_wire[267];							inform_L[134][9] = l_cell_wire[268];							inform_L[646][9] = l_cell_wire[269];							inform_L[135][9] = l_cell_wire[270];							inform_L[647][9] = l_cell_wire[271];							inform_L[136][9] = l_cell_wire[272];							inform_L[648][9] = l_cell_wire[273];							inform_L[137][9] = l_cell_wire[274];							inform_L[649][9] = l_cell_wire[275];							inform_L[138][9] = l_cell_wire[276];							inform_L[650][9] = l_cell_wire[277];							inform_L[139][9] = l_cell_wire[278];							inform_L[651][9] = l_cell_wire[279];							inform_L[140][9] = l_cell_wire[280];							inform_L[652][9] = l_cell_wire[281];							inform_L[141][9] = l_cell_wire[282];							inform_L[653][9] = l_cell_wire[283];							inform_L[142][9] = l_cell_wire[284];							inform_L[654][9] = l_cell_wire[285];							inform_L[143][9] = l_cell_wire[286];							inform_L[655][9] = l_cell_wire[287];							inform_L[144][9] = l_cell_wire[288];							inform_L[656][9] = l_cell_wire[289];							inform_L[145][9] = l_cell_wire[290];							inform_L[657][9] = l_cell_wire[291];							inform_L[146][9] = l_cell_wire[292];							inform_L[658][9] = l_cell_wire[293];							inform_L[147][9] = l_cell_wire[294];							inform_L[659][9] = l_cell_wire[295];							inform_L[148][9] = l_cell_wire[296];							inform_L[660][9] = l_cell_wire[297];							inform_L[149][9] = l_cell_wire[298];							inform_L[661][9] = l_cell_wire[299];							inform_L[150][9] = l_cell_wire[300];							inform_L[662][9] = l_cell_wire[301];							inform_L[151][9] = l_cell_wire[302];							inform_L[663][9] = l_cell_wire[303];							inform_L[152][9] = l_cell_wire[304];							inform_L[664][9] = l_cell_wire[305];							inform_L[153][9] = l_cell_wire[306];							inform_L[665][9] = l_cell_wire[307];							inform_L[154][9] = l_cell_wire[308];							inform_L[666][9] = l_cell_wire[309];							inform_L[155][9] = l_cell_wire[310];							inform_L[667][9] = l_cell_wire[311];							inform_L[156][9] = l_cell_wire[312];							inform_L[668][9] = l_cell_wire[313];							inform_L[157][9] = l_cell_wire[314];							inform_L[669][9] = l_cell_wire[315];							inform_L[158][9] = l_cell_wire[316];							inform_L[670][9] = l_cell_wire[317];							inform_L[159][9] = l_cell_wire[318];							inform_L[671][9] = l_cell_wire[319];							inform_L[160][9] = l_cell_wire[320];							inform_L[672][9] = l_cell_wire[321];							inform_L[161][9] = l_cell_wire[322];							inform_L[673][9] = l_cell_wire[323];							inform_L[162][9] = l_cell_wire[324];							inform_L[674][9] = l_cell_wire[325];							inform_L[163][9] = l_cell_wire[326];							inform_L[675][9] = l_cell_wire[327];							inform_L[164][9] = l_cell_wire[328];							inform_L[676][9] = l_cell_wire[329];							inform_L[165][9] = l_cell_wire[330];							inform_L[677][9] = l_cell_wire[331];							inform_L[166][9] = l_cell_wire[332];							inform_L[678][9] = l_cell_wire[333];							inform_L[167][9] = l_cell_wire[334];							inform_L[679][9] = l_cell_wire[335];							inform_L[168][9] = l_cell_wire[336];							inform_L[680][9] = l_cell_wire[337];							inform_L[169][9] = l_cell_wire[338];							inform_L[681][9] = l_cell_wire[339];							inform_L[170][9] = l_cell_wire[340];							inform_L[682][9] = l_cell_wire[341];							inform_L[171][9] = l_cell_wire[342];							inform_L[683][9] = l_cell_wire[343];							inform_L[172][9] = l_cell_wire[344];							inform_L[684][9] = l_cell_wire[345];							inform_L[173][9] = l_cell_wire[346];							inform_L[685][9] = l_cell_wire[347];							inform_L[174][9] = l_cell_wire[348];							inform_L[686][9] = l_cell_wire[349];							inform_L[175][9] = l_cell_wire[350];							inform_L[687][9] = l_cell_wire[351];							inform_L[176][9] = l_cell_wire[352];							inform_L[688][9] = l_cell_wire[353];							inform_L[177][9] = l_cell_wire[354];							inform_L[689][9] = l_cell_wire[355];							inform_L[178][9] = l_cell_wire[356];							inform_L[690][9] = l_cell_wire[357];							inform_L[179][9] = l_cell_wire[358];							inform_L[691][9] = l_cell_wire[359];							inform_L[180][9] = l_cell_wire[360];							inform_L[692][9] = l_cell_wire[361];							inform_L[181][9] = l_cell_wire[362];							inform_L[693][9] = l_cell_wire[363];							inform_L[182][9] = l_cell_wire[364];							inform_L[694][9] = l_cell_wire[365];							inform_L[183][9] = l_cell_wire[366];							inform_L[695][9] = l_cell_wire[367];							inform_L[184][9] = l_cell_wire[368];							inform_L[696][9] = l_cell_wire[369];							inform_L[185][9] = l_cell_wire[370];							inform_L[697][9] = l_cell_wire[371];							inform_L[186][9] = l_cell_wire[372];							inform_L[698][9] = l_cell_wire[373];							inform_L[187][9] = l_cell_wire[374];							inform_L[699][9] = l_cell_wire[375];							inform_L[188][9] = l_cell_wire[376];							inform_L[700][9] = l_cell_wire[377];							inform_L[189][9] = l_cell_wire[378];							inform_L[701][9] = l_cell_wire[379];							inform_L[190][9] = l_cell_wire[380];							inform_L[702][9] = l_cell_wire[381];							inform_L[191][9] = l_cell_wire[382];							inform_L[703][9] = l_cell_wire[383];							inform_L[192][9] = l_cell_wire[384];							inform_L[704][9] = l_cell_wire[385];							inform_L[193][9] = l_cell_wire[386];							inform_L[705][9] = l_cell_wire[387];							inform_L[194][9] = l_cell_wire[388];							inform_L[706][9] = l_cell_wire[389];							inform_L[195][9] = l_cell_wire[390];							inform_L[707][9] = l_cell_wire[391];							inform_L[196][9] = l_cell_wire[392];							inform_L[708][9] = l_cell_wire[393];							inform_L[197][9] = l_cell_wire[394];							inform_L[709][9] = l_cell_wire[395];							inform_L[198][9] = l_cell_wire[396];							inform_L[710][9] = l_cell_wire[397];							inform_L[199][9] = l_cell_wire[398];							inform_L[711][9] = l_cell_wire[399];							inform_L[200][9] = l_cell_wire[400];							inform_L[712][9] = l_cell_wire[401];							inform_L[201][9] = l_cell_wire[402];							inform_L[713][9] = l_cell_wire[403];							inform_L[202][9] = l_cell_wire[404];							inform_L[714][9] = l_cell_wire[405];							inform_L[203][9] = l_cell_wire[406];							inform_L[715][9] = l_cell_wire[407];							inform_L[204][9] = l_cell_wire[408];							inform_L[716][9] = l_cell_wire[409];							inform_L[205][9] = l_cell_wire[410];							inform_L[717][9] = l_cell_wire[411];							inform_L[206][9] = l_cell_wire[412];							inform_L[718][9] = l_cell_wire[413];							inform_L[207][9] = l_cell_wire[414];							inform_L[719][9] = l_cell_wire[415];							inform_L[208][9] = l_cell_wire[416];							inform_L[720][9] = l_cell_wire[417];							inform_L[209][9] = l_cell_wire[418];							inform_L[721][9] = l_cell_wire[419];							inform_L[210][9] = l_cell_wire[420];							inform_L[722][9] = l_cell_wire[421];							inform_L[211][9] = l_cell_wire[422];							inform_L[723][9] = l_cell_wire[423];							inform_L[212][9] = l_cell_wire[424];							inform_L[724][9] = l_cell_wire[425];							inform_L[213][9] = l_cell_wire[426];							inform_L[725][9] = l_cell_wire[427];							inform_L[214][9] = l_cell_wire[428];							inform_L[726][9] = l_cell_wire[429];							inform_L[215][9] = l_cell_wire[430];							inform_L[727][9] = l_cell_wire[431];							inform_L[216][9] = l_cell_wire[432];							inform_L[728][9] = l_cell_wire[433];							inform_L[217][9] = l_cell_wire[434];							inform_L[729][9] = l_cell_wire[435];							inform_L[218][9] = l_cell_wire[436];							inform_L[730][9] = l_cell_wire[437];							inform_L[219][9] = l_cell_wire[438];							inform_L[731][9] = l_cell_wire[439];							inform_L[220][9] = l_cell_wire[440];							inform_L[732][9] = l_cell_wire[441];							inform_L[221][9] = l_cell_wire[442];							inform_L[733][9] = l_cell_wire[443];							inform_L[222][9] = l_cell_wire[444];							inform_L[734][9] = l_cell_wire[445];							inform_L[223][9] = l_cell_wire[446];							inform_L[735][9] = l_cell_wire[447];							inform_L[224][9] = l_cell_wire[448];							inform_L[736][9] = l_cell_wire[449];							inform_L[225][9] = l_cell_wire[450];							inform_L[737][9] = l_cell_wire[451];							inform_L[226][9] = l_cell_wire[452];							inform_L[738][9] = l_cell_wire[453];							inform_L[227][9] = l_cell_wire[454];							inform_L[739][9] = l_cell_wire[455];							inform_L[228][9] = l_cell_wire[456];							inform_L[740][9] = l_cell_wire[457];							inform_L[229][9] = l_cell_wire[458];							inform_L[741][9] = l_cell_wire[459];							inform_L[230][9] = l_cell_wire[460];							inform_L[742][9] = l_cell_wire[461];							inform_L[231][9] = l_cell_wire[462];							inform_L[743][9] = l_cell_wire[463];							inform_L[232][9] = l_cell_wire[464];							inform_L[744][9] = l_cell_wire[465];							inform_L[233][9] = l_cell_wire[466];							inform_L[745][9] = l_cell_wire[467];							inform_L[234][9] = l_cell_wire[468];							inform_L[746][9] = l_cell_wire[469];							inform_L[235][9] = l_cell_wire[470];							inform_L[747][9] = l_cell_wire[471];							inform_L[236][9] = l_cell_wire[472];							inform_L[748][9] = l_cell_wire[473];							inform_L[237][9] = l_cell_wire[474];							inform_L[749][9] = l_cell_wire[475];							inform_L[238][9] = l_cell_wire[476];							inform_L[750][9] = l_cell_wire[477];							inform_L[239][9] = l_cell_wire[478];							inform_L[751][9] = l_cell_wire[479];							inform_L[240][9] = l_cell_wire[480];							inform_L[752][9] = l_cell_wire[481];							inform_L[241][9] = l_cell_wire[482];							inform_L[753][9] = l_cell_wire[483];							inform_L[242][9] = l_cell_wire[484];							inform_L[754][9] = l_cell_wire[485];							inform_L[243][9] = l_cell_wire[486];							inform_L[755][9] = l_cell_wire[487];							inform_L[244][9] = l_cell_wire[488];							inform_L[756][9] = l_cell_wire[489];							inform_L[245][9] = l_cell_wire[490];							inform_L[757][9] = l_cell_wire[491];							inform_L[246][9] = l_cell_wire[492];							inform_L[758][9] = l_cell_wire[493];							inform_L[247][9] = l_cell_wire[494];							inform_L[759][9] = l_cell_wire[495];							inform_L[248][9] = l_cell_wire[496];							inform_L[760][9] = l_cell_wire[497];							inform_L[249][9] = l_cell_wire[498];							inform_L[761][9] = l_cell_wire[499];							inform_L[250][9] = l_cell_wire[500];							inform_L[762][9] = l_cell_wire[501];							inform_L[251][9] = l_cell_wire[502];							inform_L[763][9] = l_cell_wire[503];							inform_L[252][9] = l_cell_wire[504];							inform_L[764][9] = l_cell_wire[505];							inform_L[253][9] = l_cell_wire[506];							inform_L[765][9] = l_cell_wire[507];							inform_L[254][9] = l_cell_wire[508];							inform_L[766][9] = l_cell_wire[509];							inform_L[255][9] = l_cell_wire[510];							inform_L[767][9] = l_cell_wire[511];							inform_L[256][9] = l_cell_wire[512];							inform_L[768][9] = l_cell_wire[513];							inform_L[257][9] = l_cell_wire[514];							inform_L[769][9] = l_cell_wire[515];							inform_L[258][9] = l_cell_wire[516];							inform_L[770][9] = l_cell_wire[517];							inform_L[259][9] = l_cell_wire[518];							inform_L[771][9] = l_cell_wire[519];							inform_L[260][9] = l_cell_wire[520];							inform_L[772][9] = l_cell_wire[521];							inform_L[261][9] = l_cell_wire[522];							inform_L[773][9] = l_cell_wire[523];							inform_L[262][9] = l_cell_wire[524];							inform_L[774][9] = l_cell_wire[525];							inform_L[263][9] = l_cell_wire[526];							inform_L[775][9] = l_cell_wire[527];							inform_L[264][9] = l_cell_wire[528];							inform_L[776][9] = l_cell_wire[529];							inform_L[265][9] = l_cell_wire[530];							inform_L[777][9] = l_cell_wire[531];							inform_L[266][9] = l_cell_wire[532];							inform_L[778][9] = l_cell_wire[533];							inform_L[267][9] = l_cell_wire[534];							inform_L[779][9] = l_cell_wire[535];							inform_L[268][9] = l_cell_wire[536];							inform_L[780][9] = l_cell_wire[537];							inform_L[269][9] = l_cell_wire[538];							inform_L[781][9] = l_cell_wire[539];							inform_L[270][9] = l_cell_wire[540];							inform_L[782][9] = l_cell_wire[541];							inform_L[271][9] = l_cell_wire[542];							inform_L[783][9] = l_cell_wire[543];							inform_L[272][9] = l_cell_wire[544];							inform_L[784][9] = l_cell_wire[545];							inform_L[273][9] = l_cell_wire[546];							inform_L[785][9] = l_cell_wire[547];							inform_L[274][9] = l_cell_wire[548];							inform_L[786][9] = l_cell_wire[549];							inform_L[275][9] = l_cell_wire[550];							inform_L[787][9] = l_cell_wire[551];							inform_L[276][9] = l_cell_wire[552];							inform_L[788][9] = l_cell_wire[553];							inform_L[277][9] = l_cell_wire[554];							inform_L[789][9] = l_cell_wire[555];							inform_L[278][9] = l_cell_wire[556];							inform_L[790][9] = l_cell_wire[557];							inform_L[279][9] = l_cell_wire[558];							inform_L[791][9] = l_cell_wire[559];							inform_L[280][9] = l_cell_wire[560];							inform_L[792][9] = l_cell_wire[561];							inform_L[281][9] = l_cell_wire[562];							inform_L[793][9] = l_cell_wire[563];							inform_L[282][9] = l_cell_wire[564];							inform_L[794][9] = l_cell_wire[565];							inform_L[283][9] = l_cell_wire[566];							inform_L[795][9] = l_cell_wire[567];							inform_L[284][9] = l_cell_wire[568];							inform_L[796][9] = l_cell_wire[569];							inform_L[285][9] = l_cell_wire[570];							inform_L[797][9] = l_cell_wire[571];							inform_L[286][9] = l_cell_wire[572];							inform_L[798][9] = l_cell_wire[573];							inform_L[287][9] = l_cell_wire[574];							inform_L[799][9] = l_cell_wire[575];							inform_L[288][9] = l_cell_wire[576];							inform_L[800][9] = l_cell_wire[577];							inform_L[289][9] = l_cell_wire[578];							inform_L[801][9] = l_cell_wire[579];							inform_L[290][9] = l_cell_wire[580];							inform_L[802][9] = l_cell_wire[581];							inform_L[291][9] = l_cell_wire[582];							inform_L[803][9] = l_cell_wire[583];							inform_L[292][9] = l_cell_wire[584];							inform_L[804][9] = l_cell_wire[585];							inform_L[293][9] = l_cell_wire[586];							inform_L[805][9] = l_cell_wire[587];							inform_L[294][9] = l_cell_wire[588];							inform_L[806][9] = l_cell_wire[589];							inform_L[295][9] = l_cell_wire[590];							inform_L[807][9] = l_cell_wire[591];							inform_L[296][9] = l_cell_wire[592];							inform_L[808][9] = l_cell_wire[593];							inform_L[297][9] = l_cell_wire[594];							inform_L[809][9] = l_cell_wire[595];							inform_L[298][9] = l_cell_wire[596];							inform_L[810][9] = l_cell_wire[597];							inform_L[299][9] = l_cell_wire[598];							inform_L[811][9] = l_cell_wire[599];							inform_L[300][9] = l_cell_wire[600];							inform_L[812][9] = l_cell_wire[601];							inform_L[301][9] = l_cell_wire[602];							inform_L[813][9] = l_cell_wire[603];							inform_L[302][9] = l_cell_wire[604];							inform_L[814][9] = l_cell_wire[605];							inform_L[303][9] = l_cell_wire[606];							inform_L[815][9] = l_cell_wire[607];							inform_L[304][9] = l_cell_wire[608];							inform_L[816][9] = l_cell_wire[609];							inform_L[305][9] = l_cell_wire[610];							inform_L[817][9] = l_cell_wire[611];							inform_L[306][9] = l_cell_wire[612];							inform_L[818][9] = l_cell_wire[613];							inform_L[307][9] = l_cell_wire[614];							inform_L[819][9] = l_cell_wire[615];							inform_L[308][9] = l_cell_wire[616];							inform_L[820][9] = l_cell_wire[617];							inform_L[309][9] = l_cell_wire[618];							inform_L[821][9] = l_cell_wire[619];							inform_L[310][9] = l_cell_wire[620];							inform_L[822][9] = l_cell_wire[621];							inform_L[311][9] = l_cell_wire[622];							inform_L[823][9] = l_cell_wire[623];							inform_L[312][9] = l_cell_wire[624];							inform_L[824][9] = l_cell_wire[625];							inform_L[313][9] = l_cell_wire[626];							inform_L[825][9] = l_cell_wire[627];							inform_L[314][9] = l_cell_wire[628];							inform_L[826][9] = l_cell_wire[629];							inform_L[315][9] = l_cell_wire[630];							inform_L[827][9] = l_cell_wire[631];							inform_L[316][9] = l_cell_wire[632];							inform_L[828][9] = l_cell_wire[633];							inform_L[317][9] = l_cell_wire[634];							inform_L[829][9] = l_cell_wire[635];							inform_L[318][9] = l_cell_wire[636];							inform_L[830][9] = l_cell_wire[637];							inform_L[319][9] = l_cell_wire[638];							inform_L[831][9] = l_cell_wire[639];							inform_L[320][9] = l_cell_wire[640];							inform_L[832][9] = l_cell_wire[641];							inform_L[321][9] = l_cell_wire[642];							inform_L[833][9] = l_cell_wire[643];							inform_L[322][9] = l_cell_wire[644];							inform_L[834][9] = l_cell_wire[645];							inform_L[323][9] = l_cell_wire[646];							inform_L[835][9] = l_cell_wire[647];							inform_L[324][9] = l_cell_wire[648];							inform_L[836][9] = l_cell_wire[649];							inform_L[325][9] = l_cell_wire[650];							inform_L[837][9] = l_cell_wire[651];							inform_L[326][9] = l_cell_wire[652];							inform_L[838][9] = l_cell_wire[653];							inform_L[327][9] = l_cell_wire[654];							inform_L[839][9] = l_cell_wire[655];							inform_L[328][9] = l_cell_wire[656];							inform_L[840][9] = l_cell_wire[657];							inform_L[329][9] = l_cell_wire[658];							inform_L[841][9] = l_cell_wire[659];							inform_L[330][9] = l_cell_wire[660];							inform_L[842][9] = l_cell_wire[661];							inform_L[331][9] = l_cell_wire[662];							inform_L[843][9] = l_cell_wire[663];							inform_L[332][9] = l_cell_wire[664];							inform_L[844][9] = l_cell_wire[665];							inform_L[333][9] = l_cell_wire[666];							inform_L[845][9] = l_cell_wire[667];							inform_L[334][9] = l_cell_wire[668];							inform_L[846][9] = l_cell_wire[669];							inform_L[335][9] = l_cell_wire[670];							inform_L[847][9] = l_cell_wire[671];							inform_L[336][9] = l_cell_wire[672];							inform_L[848][9] = l_cell_wire[673];							inform_L[337][9] = l_cell_wire[674];							inform_L[849][9] = l_cell_wire[675];							inform_L[338][9] = l_cell_wire[676];							inform_L[850][9] = l_cell_wire[677];							inform_L[339][9] = l_cell_wire[678];							inform_L[851][9] = l_cell_wire[679];							inform_L[340][9] = l_cell_wire[680];							inform_L[852][9] = l_cell_wire[681];							inform_L[341][9] = l_cell_wire[682];							inform_L[853][9] = l_cell_wire[683];							inform_L[342][9] = l_cell_wire[684];							inform_L[854][9] = l_cell_wire[685];							inform_L[343][9] = l_cell_wire[686];							inform_L[855][9] = l_cell_wire[687];							inform_L[344][9] = l_cell_wire[688];							inform_L[856][9] = l_cell_wire[689];							inform_L[345][9] = l_cell_wire[690];							inform_L[857][9] = l_cell_wire[691];							inform_L[346][9] = l_cell_wire[692];							inform_L[858][9] = l_cell_wire[693];							inform_L[347][9] = l_cell_wire[694];							inform_L[859][9] = l_cell_wire[695];							inform_L[348][9] = l_cell_wire[696];							inform_L[860][9] = l_cell_wire[697];							inform_L[349][9] = l_cell_wire[698];							inform_L[861][9] = l_cell_wire[699];							inform_L[350][9] = l_cell_wire[700];							inform_L[862][9] = l_cell_wire[701];							inform_L[351][9] = l_cell_wire[702];							inform_L[863][9] = l_cell_wire[703];							inform_L[352][9] = l_cell_wire[704];							inform_L[864][9] = l_cell_wire[705];							inform_L[353][9] = l_cell_wire[706];							inform_L[865][9] = l_cell_wire[707];							inform_L[354][9] = l_cell_wire[708];							inform_L[866][9] = l_cell_wire[709];							inform_L[355][9] = l_cell_wire[710];							inform_L[867][9] = l_cell_wire[711];							inform_L[356][9] = l_cell_wire[712];							inform_L[868][9] = l_cell_wire[713];							inform_L[357][9] = l_cell_wire[714];							inform_L[869][9] = l_cell_wire[715];							inform_L[358][9] = l_cell_wire[716];							inform_L[870][9] = l_cell_wire[717];							inform_L[359][9] = l_cell_wire[718];							inform_L[871][9] = l_cell_wire[719];							inform_L[360][9] = l_cell_wire[720];							inform_L[872][9] = l_cell_wire[721];							inform_L[361][9] = l_cell_wire[722];							inform_L[873][9] = l_cell_wire[723];							inform_L[362][9] = l_cell_wire[724];							inform_L[874][9] = l_cell_wire[725];							inform_L[363][9] = l_cell_wire[726];							inform_L[875][9] = l_cell_wire[727];							inform_L[364][9] = l_cell_wire[728];							inform_L[876][9] = l_cell_wire[729];							inform_L[365][9] = l_cell_wire[730];							inform_L[877][9] = l_cell_wire[731];							inform_L[366][9] = l_cell_wire[732];							inform_L[878][9] = l_cell_wire[733];							inform_L[367][9] = l_cell_wire[734];							inform_L[879][9] = l_cell_wire[735];							inform_L[368][9] = l_cell_wire[736];							inform_L[880][9] = l_cell_wire[737];							inform_L[369][9] = l_cell_wire[738];							inform_L[881][9] = l_cell_wire[739];							inform_L[370][9] = l_cell_wire[740];							inform_L[882][9] = l_cell_wire[741];							inform_L[371][9] = l_cell_wire[742];							inform_L[883][9] = l_cell_wire[743];							inform_L[372][9] = l_cell_wire[744];							inform_L[884][9] = l_cell_wire[745];							inform_L[373][9] = l_cell_wire[746];							inform_L[885][9] = l_cell_wire[747];							inform_L[374][9] = l_cell_wire[748];							inform_L[886][9] = l_cell_wire[749];							inform_L[375][9] = l_cell_wire[750];							inform_L[887][9] = l_cell_wire[751];							inform_L[376][9] = l_cell_wire[752];							inform_L[888][9] = l_cell_wire[753];							inform_L[377][9] = l_cell_wire[754];							inform_L[889][9] = l_cell_wire[755];							inform_L[378][9] = l_cell_wire[756];							inform_L[890][9] = l_cell_wire[757];							inform_L[379][9] = l_cell_wire[758];							inform_L[891][9] = l_cell_wire[759];							inform_L[380][9] = l_cell_wire[760];							inform_L[892][9] = l_cell_wire[761];							inform_L[381][9] = l_cell_wire[762];							inform_L[893][9] = l_cell_wire[763];							inform_L[382][9] = l_cell_wire[764];							inform_L[894][9] = l_cell_wire[765];							inform_L[383][9] = l_cell_wire[766];							inform_L[895][9] = l_cell_wire[767];							inform_L[384][9] = l_cell_wire[768];							inform_L[896][9] = l_cell_wire[769];							inform_L[385][9] = l_cell_wire[770];							inform_L[897][9] = l_cell_wire[771];							inform_L[386][9] = l_cell_wire[772];							inform_L[898][9] = l_cell_wire[773];							inform_L[387][9] = l_cell_wire[774];							inform_L[899][9] = l_cell_wire[775];							inform_L[388][9] = l_cell_wire[776];							inform_L[900][9] = l_cell_wire[777];							inform_L[389][9] = l_cell_wire[778];							inform_L[901][9] = l_cell_wire[779];							inform_L[390][9] = l_cell_wire[780];							inform_L[902][9] = l_cell_wire[781];							inform_L[391][9] = l_cell_wire[782];							inform_L[903][9] = l_cell_wire[783];							inform_L[392][9] = l_cell_wire[784];							inform_L[904][9] = l_cell_wire[785];							inform_L[393][9] = l_cell_wire[786];							inform_L[905][9] = l_cell_wire[787];							inform_L[394][9] = l_cell_wire[788];							inform_L[906][9] = l_cell_wire[789];							inform_L[395][9] = l_cell_wire[790];							inform_L[907][9] = l_cell_wire[791];							inform_L[396][9] = l_cell_wire[792];							inform_L[908][9] = l_cell_wire[793];							inform_L[397][9] = l_cell_wire[794];							inform_L[909][9] = l_cell_wire[795];							inform_L[398][9] = l_cell_wire[796];							inform_L[910][9] = l_cell_wire[797];							inform_L[399][9] = l_cell_wire[798];							inform_L[911][9] = l_cell_wire[799];							inform_L[400][9] = l_cell_wire[800];							inform_L[912][9] = l_cell_wire[801];							inform_L[401][9] = l_cell_wire[802];							inform_L[913][9] = l_cell_wire[803];							inform_L[402][9] = l_cell_wire[804];							inform_L[914][9] = l_cell_wire[805];							inform_L[403][9] = l_cell_wire[806];							inform_L[915][9] = l_cell_wire[807];							inform_L[404][9] = l_cell_wire[808];							inform_L[916][9] = l_cell_wire[809];							inform_L[405][9] = l_cell_wire[810];							inform_L[917][9] = l_cell_wire[811];							inform_L[406][9] = l_cell_wire[812];							inform_L[918][9] = l_cell_wire[813];							inform_L[407][9] = l_cell_wire[814];							inform_L[919][9] = l_cell_wire[815];							inform_L[408][9] = l_cell_wire[816];							inform_L[920][9] = l_cell_wire[817];							inform_L[409][9] = l_cell_wire[818];							inform_L[921][9] = l_cell_wire[819];							inform_L[410][9] = l_cell_wire[820];							inform_L[922][9] = l_cell_wire[821];							inform_L[411][9] = l_cell_wire[822];							inform_L[923][9] = l_cell_wire[823];							inform_L[412][9] = l_cell_wire[824];							inform_L[924][9] = l_cell_wire[825];							inform_L[413][9] = l_cell_wire[826];							inform_L[925][9] = l_cell_wire[827];							inform_L[414][9] = l_cell_wire[828];							inform_L[926][9] = l_cell_wire[829];							inform_L[415][9] = l_cell_wire[830];							inform_L[927][9] = l_cell_wire[831];							inform_L[416][9] = l_cell_wire[832];							inform_L[928][9] = l_cell_wire[833];							inform_L[417][9] = l_cell_wire[834];							inform_L[929][9] = l_cell_wire[835];							inform_L[418][9] = l_cell_wire[836];							inform_L[930][9] = l_cell_wire[837];							inform_L[419][9] = l_cell_wire[838];							inform_L[931][9] = l_cell_wire[839];							inform_L[420][9] = l_cell_wire[840];							inform_L[932][9] = l_cell_wire[841];							inform_L[421][9] = l_cell_wire[842];							inform_L[933][9] = l_cell_wire[843];							inform_L[422][9] = l_cell_wire[844];							inform_L[934][9] = l_cell_wire[845];							inform_L[423][9] = l_cell_wire[846];							inform_L[935][9] = l_cell_wire[847];							inform_L[424][9] = l_cell_wire[848];							inform_L[936][9] = l_cell_wire[849];							inform_L[425][9] = l_cell_wire[850];							inform_L[937][9] = l_cell_wire[851];							inform_L[426][9] = l_cell_wire[852];							inform_L[938][9] = l_cell_wire[853];							inform_L[427][9] = l_cell_wire[854];							inform_L[939][9] = l_cell_wire[855];							inform_L[428][9] = l_cell_wire[856];							inform_L[940][9] = l_cell_wire[857];							inform_L[429][9] = l_cell_wire[858];							inform_L[941][9] = l_cell_wire[859];							inform_L[430][9] = l_cell_wire[860];							inform_L[942][9] = l_cell_wire[861];							inform_L[431][9] = l_cell_wire[862];							inform_L[943][9] = l_cell_wire[863];							inform_L[432][9] = l_cell_wire[864];							inform_L[944][9] = l_cell_wire[865];							inform_L[433][9] = l_cell_wire[866];							inform_L[945][9] = l_cell_wire[867];							inform_L[434][9] = l_cell_wire[868];							inform_L[946][9] = l_cell_wire[869];							inform_L[435][9] = l_cell_wire[870];							inform_L[947][9] = l_cell_wire[871];							inform_L[436][9] = l_cell_wire[872];							inform_L[948][9] = l_cell_wire[873];							inform_L[437][9] = l_cell_wire[874];							inform_L[949][9] = l_cell_wire[875];							inform_L[438][9] = l_cell_wire[876];							inform_L[950][9] = l_cell_wire[877];							inform_L[439][9] = l_cell_wire[878];							inform_L[951][9] = l_cell_wire[879];							inform_L[440][9] = l_cell_wire[880];							inform_L[952][9] = l_cell_wire[881];							inform_L[441][9] = l_cell_wire[882];							inform_L[953][9] = l_cell_wire[883];							inform_L[442][9] = l_cell_wire[884];							inform_L[954][9] = l_cell_wire[885];							inform_L[443][9] = l_cell_wire[886];							inform_L[955][9] = l_cell_wire[887];							inform_L[444][9] = l_cell_wire[888];							inform_L[956][9] = l_cell_wire[889];							inform_L[445][9] = l_cell_wire[890];							inform_L[957][9] = l_cell_wire[891];							inform_L[446][9] = l_cell_wire[892];							inform_L[958][9] = l_cell_wire[893];							inform_L[447][9] = l_cell_wire[894];							inform_L[959][9] = l_cell_wire[895];							inform_L[448][9] = l_cell_wire[896];							inform_L[960][9] = l_cell_wire[897];							inform_L[449][9] = l_cell_wire[898];							inform_L[961][9] = l_cell_wire[899];							inform_L[450][9] = l_cell_wire[900];							inform_L[962][9] = l_cell_wire[901];							inform_L[451][9] = l_cell_wire[902];							inform_L[963][9] = l_cell_wire[903];							inform_L[452][9] = l_cell_wire[904];							inform_L[964][9] = l_cell_wire[905];							inform_L[453][9] = l_cell_wire[906];							inform_L[965][9] = l_cell_wire[907];							inform_L[454][9] = l_cell_wire[908];							inform_L[966][9] = l_cell_wire[909];							inform_L[455][9] = l_cell_wire[910];							inform_L[967][9] = l_cell_wire[911];							inform_L[456][9] = l_cell_wire[912];							inform_L[968][9] = l_cell_wire[913];							inform_L[457][9] = l_cell_wire[914];							inform_L[969][9] = l_cell_wire[915];							inform_L[458][9] = l_cell_wire[916];							inform_L[970][9] = l_cell_wire[917];							inform_L[459][9] = l_cell_wire[918];							inform_L[971][9] = l_cell_wire[919];							inform_L[460][9] = l_cell_wire[920];							inform_L[972][9] = l_cell_wire[921];							inform_L[461][9] = l_cell_wire[922];							inform_L[973][9] = l_cell_wire[923];							inform_L[462][9] = l_cell_wire[924];							inform_L[974][9] = l_cell_wire[925];							inform_L[463][9] = l_cell_wire[926];							inform_L[975][9] = l_cell_wire[927];							inform_L[464][9] = l_cell_wire[928];							inform_L[976][9] = l_cell_wire[929];							inform_L[465][9] = l_cell_wire[930];							inform_L[977][9] = l_cell_wire[931];							inform_L[466][9] = l_cell_wire[932];							inform_L[978][9] = l_cell_wire[933];							inform_L[467][9] = l_cell_wire[934];							inform_L[979][9] = l_cell_wire[935];							inform_L[468][9] = l_cell_wire[936];							inform_L[980][9] = l_cell_wire[937];							inform_L[469][9] = l_cell_wire[938];							inform_L[981][9] = l_cell_wire[939];							inform_L[470][9] = l_cell_wire[940];							inform_L[982][9] = l_cell_wire[941];							inform_L[471][9] = l_cell_wire[942];							inform_L[983][9] = l_cell_wire[943];							inform_L[472][9] = l_cell_wire[944];							inform_L[984][9] = l_cell_wire[945];							inform_L[473][9] = l_cell_wire[946];							inform_L[985][9] = l_cell_wire[947];							inform_L[474][9] = l_cell_wire[948];							inform_L[986][9] = l_cell_wire[949];							inform_L[475][9] = l_cell_wire[950];							inform_L[987][9] = l_cell_wire[951];							inform_L[476][9] = l_cell_wire[952];							inform_L[988][9] = l_cell_wire[953];							inform_L[477][9] = l_cell_wire[954];							inform_L[989][9] = l_cell_wire[955];							inform_L[478][9] = l_cell_wire[956];							inform_L[990][9] = l_cell_wire[957];							inform_L[479][9] = l_cell_wire[958];							inform_L[991][9] = l_cell_wire[959];							inform_L[480][9] = l_cell_wire[960];							inform_L[992][9] = l_cell_wire[961];							inform_L[481][9] = l_cell_wire[962];							inform_L[993][9] = l_cell_wire[963];							inform_L[482][9] = l_cell_wire[964];							inform_L[994][9] = l_cell_wire[965];							inform_L[483][9] = l_cell_wire[966];							inform_L[995][9] = l_cell_wire[967];							inform_L[484][9] = l_cell_wire[968];							inform_L[996][9] = l_cell_wire[969];							inform_L[485][9] = l_cell_wire[970];							inform_L[997][9] = l_cell_wire[971];							inform_L[486][9] = l_cell_wire[972];							inform_L[998][9] = l_cell_wire[973];							inform_L[487][9] = l_cell_wire[974];							inform_L[999][9] = l_cell_wire[975];							inform_L[488][9] = l_cell_wire[976];							inform_L[1000][9] = l_cell_wire[977];							inform_L[489][9] = l_cell_wire[978];							inform_L[1001][9] = l_cell_wire[979];							inform_L[490][9] = l_cell_wire[980];							inform_L[1002][9] = l_cell_wire[981];							inform_L[491][9] = l_cell_wire[982];							inform_L[1003][9] = l_cell_wire[983];							inform_L[492][9] = l_cell_wire[984];							inform_L[1004][9] = l_cell_wire[985];							inform_L[493][9] = l_cell_wire[986];							inform_L[1005][9] = l_cell_wire[987];							inform_L[494][9] = l_cell_wire[988];							inform_L[1006][9] = l_cell_wire[989];							inform_L[495][9] = l_cell_wire[990];							inform_L[1007][9] = l_cell_wire[991];							inform_L[496][9] = l_cell_wire[992];							inform_L[1008][9] = l_cell_wire[993];							inform_L[497][9] = l_cell_wire[994];							inform_L[1009][9] = l_cell_wire[995];							inform_L[498][9] = l_cell_wire[996];							inform_L[1010][9] = l_cell_wire[997];							inform_L[499][9] = l_cell_wire[998];							inform_L[1011][9] = l_cell_wire[999];							inform_L[500][9] = l_cell_wire[1000];							inform_L[1012][9] = l_cell_wire[1001];							inform_L[501][9] = l_cell_wire[1002];							inform_L[1013][9] = l_cell_wire[1003];							inform_L[502][9] = l_cell_wire[1004];							inform_L[1014][9] = l_cell_wire[1005];							inform_L[503][9] = l_cell_wire[1006];							inform_L[1015][9] = l_cell_wire[1007];							inform_L[504][9] = l_cell_wire[1008];							inform_L[1016][9] = l_cell_wire[1009];							inform_L[505][9] = l_cell_wire[1010];							inform_L[1017][9] = l_cell_wire[1011];							inform_L[506][9] = l_cell_wire[1012];							inform_L[1018][9] = l_cell_wire[1013];							inform_L[507][9] = l_cell_wire[1014];							inform_L[1019][9] = l_cell_wire[1015];							inform_L[508][9] = l_cell_wire[1016];							inform_L[1020][9] = l_cell_wire[1017];							inform_L[509][9] = l_cell_wire[1018];							inform_L[1021][9] = l_cell_wire[1019];							inform_L[510][9] = l_cell_wire[1020];							inform_L[1022][9] = l_cell_wire[1021];							inform_L[511][9] = l_cell_wire[1022];							inform_L[1023][9] = l_cell_wire[1023];						end
						default:							for (x = 0; x < 1024; x = x + 1)								for (y = 0; y < 10; y = y + 1)								begin									inform_R[x][y+1] <= 8'd0;									inform_L[x][y] <= 8'd0;								end					endcase				end			end
			BUSY_RIGHT:			begin				if(clk_counter == 2'b11)begin					case (w2r)						1:						begin							inform_R[0][1] = r_cell_wire[0];							inform_R[1][1] = r_cell_wire[1];							inform_R[2][1] = r_cell_wire[2];							inform_R[3][1] = r_cell_wire[3];							inform_R[4][1] = r_cell_wire[4];							inform_R[5][1] = r_cell_wire[5];							inform_R[6][1] = r_cell_wire[6];							inform_R[7][1] = r_cell_wire[7];							inform_R[8][1] = r_cell_wire[8];							inform_R[9][1] = r_cell_wire[9];							inform_R[10][1] = r_cell_wire[10];							inform_R[11][1] = r_cell_wire[11];							inform_R[12][1] = r_cell_wire[12];							inform_R[13][1] = r_cell_wire[13];							inform_R[14][1] = r_cell_wire[14];							inform_R[15][1] = r_cell_wire[15];							inform_R[16][1] = r_cell_wire[16];							inform_R[17][1] = r_cell_wire[17];							inform_R[18][1] = r_cell_wire[18];							inform_R[19][1] = r_cell_wire[19];							inform_R[20][1] = r_cell_wire[20];							inform_R[21][1] = r_cell_wire[21];							inform_R[22][1] = r_cell_wire[22];							inform_R[23][1] = r_cell_wire[23];							inform_R[24][1] = r_cell_wire[24];							inform_R[25][1] = r_cell_wire[25];							inform_R[26][1] = r_cell_wire[26];							inform_R[27][1] = r_cell_wire[27];							inform_R[28][1] = r_cell_wire[28];							inform_R[29][1] = r_cell_wire[29];							inform_R[30][1] = r_cell_wire[30];							inform_R[31][1] = r_cell_wire[31];							inform_R[32][1] = r_cell_wire[32];							inform_R[33][1] = r_cell_wire[33];							inform_R[34][1] = r_cell_wire[34];							inform_R[35][1] = r_cell_wire[35];							inform_R[36][1] = r_cell_wire[36];							inform_R[37][1] = r_cell_wire[37];							inform_R[38][1] = r_cell_wire[38];							inform_R[39][1] = r_cell_wire[39];							inform_R[40][1] = r_cell_wire[40];							inform_R[41][1] = r_cell_wire[41];							inform_R[42][1] = r_cell_wire[42];							inform_R[43][1] = r_cell_wire[43];							inform_R[44][1] = r_cell_wire[44];							inform_R[45][1] = r_cell_wire[45];							inform_R[46][1] = r_cell_wire[46];							inform_R[47][1] = r_cell_wire[47];							inform_R[48][1] = r_cell_wire[48];							inform_R[49][1] = r_cell_wire[49];							inform_R[50][1] = r_cell_wire[50];							inform_R[51][1] = r_cell_wire[51];							inform_R[52][1] = r_cell_wire[52];							inform_R[53][1] = r_cell_wire[53];							inform_R[54][1] = r_cell_wire[54];							inform_R[55][1] = r_cell_wire[55];							inform_R[56][1] = r_cell_wire[56];							inform_R[57][1] = r_cell_wire[57];							inform_R[58][1] = r_cell_wire[58];							inform_R[59][1] = r_cell_wire[59];							inform_R[60][1] = r_cell_wire[60];							inform_R[61][1] = r_cell_wire[61];							inform_R[62][1] = r_cell_wire[62];							inform_R[63][1] = r_cell_wire[63];							inform_R[64][1] = r_cell_wire[64];							inform_R[65][1] = r_cell_wire[65];							inform_R[66][1] = r_cell_wire[66];							inform_R[67][1] = r_cell_wire[67];							inform_R[68][1] = r_cell_wire[68];							inform_R[69][1] = r_cell_wire[69];							inform_R[70][1] = r_cell_wire[70];							inform_R[71][1] = r_cell_wire[71];							inform_R[72][1] = r_cell_wire[72];							inform_R[73][1] = r_cell_wire[73];							inform_R[74][1] = r_cell_wire[74];							inform_R[75][1] = r_cell_wire[75];							inform_R[76][1] = r_cell_wire[76];							inform_R[77][1] = r_cell_wire[77];							inform_R[78][1] = r_cell_wire[78];							inform_R[79][1] = r_cell_wire[79];							inform_R[80][1] = r_cell_wire[80];							inform_R[81][1] = r_cell_wire[81];							inform_R[82][1] = r_cell_wire[82];							inform_R[83][1] = r_cell_wire[83];							inform_R[84][1] = r_cell_wire[84];							inform_R[85][1] = r_cell_wire[85];							inform_R[86][1] = r_cell_wire[86];							inform_R[87][1] = r_cell_wire[87];							inform_R[88][1] = r_cell_wire[88];							inform_R[89][1] = r_cell_wire[89];							inform_R[90][1] = r_cell_wire[90];							inform_R[91][1] = r_cell_wire[91];							inform_R[92][1] = r_cell_wire[92];							inform_R[93][1] = r_cell_wire[93];							inform_R[94][1] = r_cell_wire[94];							inform_R[95][1] = r_cell_wire[95];							inform_R[96][1] = r_cell_wire[96];							inform_R[97][1] = r_cell_wire[97];							inform_R[98][1] = r_cell_wire[98];							inform_R[99][1] = r_cell_wire[99];							inform_R[100][1] = r_cell_wire[100];							inform_R[101][1] = r_cell_wire[101];							inform_R[102][1] = r_cell_wire[102];							inform_R[103][1] = r_cell_wire[103];							inform_R[104][1] = r_cell_wire[104];							inform_R[105][1] = r_cell_wire[105];							inform_R[106][1] = r_cell_wire[106];							inform_R[107][1] = r_cell_wire[107];							inform_R[108][1] = r_cell_wire[108];							inform_R[109][1] = r_cell_wire[109];							inform_R[110][1] = r_cell_wire[110];							inform_R[111][1] = r_cell_wire[111];							inform_R[112][1] = r_cell_wire[112];							inform_R[113][1] = r_cell_wire[113];							inform_R[114][1] = r_cell_wire[114];							inform_R[115][1] = r_cell_wire[115];							inform_R[116][1] = r_cell_wire[116];							inform_R[117][1] = r_cell_wire[117];							inform_R[118][1] = r_cell_wire[118];							inform_R[119][1] = r_cell_wire[119];							inform_R[120][1] = r_cell_wire[120];							inform_R[121][1] = r_cell_wire[121];							inform_R[122][1] = r_cell_wire[122];							inform_R[123][1] = r_cell_wire[123];							inform_R[124][1] = r_cell_wire[124];							inform_R[125][1] = r_cell_wire[125];							inform_R[126][1] = r_cell_wire[126];							inform_R[127][1] = r_cell_wire[127];							inform_R[128][1] = r_cell_wire[128];							inform_R[129][1] = r_cell_wire[129];							inform_R[130][1] = r_cell_wire[130];							inform_R[131][1] = r_cell_wire[131];							inform_R[132][1] = r_cell_wire[132];							inform_R[133][1] = r_cell_wire[133];							inform_R[134][1] = r_cell_wire[134];							inform_R[135][1] = r_cell_wire[135];							inform_R[136][1] = r_cell_wire[136];							inform_R[137][1] = r_cell_wire[137];							inform_R[138][1] = r_cell_wire[138];							inform_R[139][1] = r_cell_wire[139];							inform_R[140][1] = r_cell_wire[140];							inform_R[141][1] = r_cell_wire[141];							inform_R[142][1] = r_cell_wire[142];							inform_R[143][1] = r_cell_wire[143];							inform_R[144][1] = r_cell_wire[144];							inform_R[145][1] = r_cell_wire[145];							inform_R[146][1] = r_cell_wire[146];							inform_R[147][1] = r_cell_wire[147];							inform_R[148][1] = r_cell_wire[148];							inform_R[149][1] = r_cell_wire[149];							inform_R[150][1] = r_cell_wire[150];							inform_R[151][1] = r_cell_wire[151];							inform_R[152][1] = r_cell_wire[152];							inform_R[153][1] = r_cell_wire[153];							inform_R[154][1] = r_cell_wire[154];							inform_R[155][1] = r_cell_wire[155];							inform_R[156][1] = r_cell_wire[156];							inform_R[157][1] = r_cell_wire[157];							inform_R[158][1] = r_cell_wire[158];							inform_R[159][1] = r_cell_wire[159];							inform_R[160][1] = r_cell_wire[160];							inform_R[161][1] = r_cell_wire[161];							inform_R[162][1] = r_cell_wire[162];							inform_R[163][1] = r_cell_wire[163];							inform_R[164][1] = r_cell_wire[164];							inform_R[165][1] = r_cell_wire[165];							inform_R[166][1] = r_cell_wire[166];							inform_R[167][1] = r_cell_wire[167];							inform_R[168][1] = r_cell_wire[168];							inform_R[169][1] = r_cell_wire[169];							inform_R[170][1] = r_cell_wire[170];							inform_R[171][1] = r_cell_wire[171];							inform_R[172][1] = r_cell_wire[172];							inform_R[173][1] = r_cell_wire[173];							inform_R[174][1] = r_cell_wire[174];							inform_R[175][1] = r_cell_wire[175];							inform_R[176][1] = r_cell_wire[176];							inform_R[177][1] = r_cell_wire[177];							inform_R[178][1] = r_cell_wire[178];							inform_R[179][1] = r_cell_wire[179];							inform_R[180][1] = r_cell_wire[180];							inform_R[181][1] = r_cell_wire[181];							inform_R[182][1] = r_cell_wire[182];							inform_R[183][1] = r_cell_wire[183];							inform_R[184][1] = r_cell_wire[184];							inform_R[185][1] = r_cell_wire[185];							inform_R[186][1] = r_cell_wire[186];							inform_R[187][1] = r_cell_wire[187];							inform_R[188][1] = r_cell_wire[188];							inform_R[189][1] = r_cell_wire[189];							inform_R[190][1] = r_cell_wire[190];							inform_R[191][1] = r_cell_wire[191];							inform_R[192][1] = r_cell_wire[192];							inform_R[193][1] = r_cell_wire[193];							inform_R[194][1] = r_cell_wire[194];							inform_R[195][1] = r_cell_wire[195];							inform_R[196][1] = r_cell_wire[196];							inform_R[197][1] = r_cell_wire[197];							inform_R[198][1] = r_cell_wire[198];							inform_R[199][1] = r_cell_wire[199];							inform_R[200][1] = r_cell_wire[200];							inform_R[201][1] = r_cell_wire[201];							inform_R[202][1] = r_cell_wire[202];							inform_R[203][1] = r_cell_wire[203];							inform_R[204][1] = r_cell_wire[204];							inform_R[205][1] = r_cell_wire[205];							inform_R[206][1] = r_cell_wire[206];							inform_R[207][1] = r_cell_wire[207];							inform_R[208][1] = r_cell_wire[208];							inform_R[209][1] = r_cell_wire[209];							inform_R[210][1] = r_cell_wire[210];							inform_R[211][1] = r_cell_wire[211];							inform_R[212][1] = r_cell_wire[212];							inform_R[213][1] = r_cell_wire[213];							inform_R[214][1] = r_cell_wire[214];							inform_R[215][1] = r_cell_wire[215];							inform_R[216][1] = r_cell_wire[216];							inform_R[217][1] = r_cell_wire[217];							inform_R[218][1] = r_cell_wire[218];							inform_R[219][1] = r_cell_wire[219];							inform_R[220][1] = r_cell_wire[220];							inform_R[221][1] = r_cell_wire[221];							inform_R[222][1] = r_cell_wire[222];							inform_R[223][1] = r_cell_wire[223];							inform_R[224][1] = r_cell_wire[224];							inform_R[225][1] = r_cell_wire[225];							inform_R[226][1] = r_cell_wire[226];							inform_R[227][1] = r_cell_wire[227];							inform_R[228][1] = r_cell_wire[228];							inform_R[229][1] = r_cell_wire[229];							inform_R[230][1] = r_cell_wire[230];							inform_R[231][1] = r_cell_wire[231];							inform_R[232][1] = r_cell_wire[232];							inform_R[233][1] = r_cell_wire[233];							inform_R[234][1] = r_cell_wire[234];							inform_R[235][1] = r_cell_wire[235];							inform_R[236][1] = r_cell_wire[236];							inform_R[237][1] = r_cell_wire[237];							inform_R[238][1] = r_cell_wire[238];							inform_R[239][1] = r_cell_wire[239];							inform_R[240][1] = r_cell_wire[240];							inform_R[241][1] = r_cell_wire[241];							inform_R[242][1] = r_cell_wire[242];							inform_R[243][1] = r_cell_wire[243];							inform_R[244][1] = r_cell_wire[244];							inform_R[245][1] = r_cell_wire[245];							inform_R[246][1] = r_cell_wire[246];							inform_R[247][1] = r_cell_wire[247];							inform_R[248][1] = r_cell_wire[248];							inform_R[249][1] = r_cell_wire[249];							inform_R[250][1] = r_cell_wire[250];							inform_R[251][1] = r_cell_wire[251];							inform_R[252][1] = r_cell_wire[252];							inform_R[253][1] = r_cell_wire[253];							inform_R[254][1] = r_cell_wire[254];							inform_R[255][1] = r_cell_wire[255];							inform_R[256][1] = r_cell_wire[256];							inform_R[257][1] = r_cell_wire[257];							inform_R[258][1] = r_cell_wire[258];							inform_R[259][1] = r_cell_wire[259];							inform_R[260][1] = r_cell_wire[260];							inform_R[261][1] = r_cell_wire[261];							inform_R[262][1] = r_cell_wire[262];							inform_R[263][1] = r_cell_wire[263];							inform_R[264][1] = r_cell_wire[264];							inform_R[265][1] = r_cell_wire[265];							inform_R[266][1] = r_cell_wire[266];							inform_R[267][1] = r_cell_wire[267];							inform_R[268][1] = r_cell_wire[268];							inform_R[269][1] = r_cell_wire[269];							inform_R[270][1] = r_cell_wire[270];							inform_R[271][1] = r_cell_wire[271];							inform_R[272][1] = r_cell_wire[272];							inform_R[273][1] = r_cell_wire[273];							inform_R[274][1] = r_cell_wire[274];							inform_R[275][1] = r_cell_wire[275];							inform_R[276][1] = r_cell_wire[276];							inform_R[277][1] = r_cell_wire[277];							inform_R[278][1] = r_cell_wire[278];							inform_R[279][1] = r_cell_wire[279];							inform_R[280][1] = r_cell_wire[280];							inform_R[281][1] = r_cell_wire[281];							inform_R[282][1] = r_cell_wire[282];							inform_R[283][1] = r_cell_wire[283];							inform_R[284][1] = r_cell_wire[284];							inform_R[285][1] = r_cell_wire[285];							inform_R[286][1] = r_cell_wire[286];							inform_R[287][1] = r_cell_wire[287];							inform_R[288][1] = r_cell_wire[288];							inform_R[289][1] = r_cell_wire[289];							inform_R[290][1] = r_cell_wire[290];							inform_R[291][1] = r_cell_wire[291];							inform_R[292][1] = r_cell_wire[292];							inform_R[293][1] = r_cell_wire[293];							inform_R[294][1] = r_cell_wire[294];							inform_R[295][1] = r_cell_wire[295];							inform_R[296][1] = r_cell_wire[296];							inform_R[297][1] = r_cell_wire[297];							inform_R[298][1] = r_cell_wire[298];							inform_R[299][1] = r_cell_wire[299];							inform_R[300][1] = r_cell_wire[300];							inform_R[301][1] = r_cell_wire[301];							inform_R[302][1] = r_cell_wire[302];							inform_R[303][1] = r_cell_wire[303];							inform_R[304][1] = r_cell_wire[304];							inform_R[305][1] = r_cell_wire[305];							inform_R[306][1] = r_cell_wire[306];							inform_R[307][1] = r_cell_wire[307];							inform_R[308][1] = r_cell_wire[308];							inform_R[309][1] = r_cell_wire[309];							inform_R[310][1] = r_cell_wire[310];							inform_R[311][1] = r_cell_wire[311];							inform_R[312][1] = r_cell_wire[312];							inform_R[313][1] = r_cell_wire[313];							inform_R[314][1] = r_cell_wire[314];							inform_R[315][1] = r_cell_wire[315];							inform_R[316][1] = r_cell_wire[316];							inform_R[317][1] = r_cell_wire[317];							inform_R[318][1] = r_cell_wire[318];							inform_R[319][1] = r_cell_wire[319];							inform_R[320][1] = r_cell_wire[320];							inform_R[321][1] = r_cell_wire[321];							inform_R[322][1] = r_cell_wire[322];							inform_R[323][1] = r_cell_wire[323];							inform_R[324][1] = r_cell_wire[324];							inform_R[325][1] = r_cell_wire[325];							inform_R[326][1] = r_cell_wire[326];							inform_R[327][1] = r_cell_wire[327];							inform_R[328][1] = r_cell_wire[328];							inform_R[329][1] = r_cell_wire[329];							inform_R[330][1] = r_cell_wire[330];							inform_R[331][1] = r_cell_wire[331];							inform_R[332][1] = r_cell_wire[332];							inform_R[333][1] = r_cell_wire[333];							inform_R[334][1] = r_cell_wire[334];							inform_R[335][1] = r_cell_wire[335];							inform_R[336][1] = r_cell_wire[336];							inform_R[337][1] = r_cell_wire[337];							inform_R[338][1] = r_cell_wire[338];							inform_R[339][1] = r_cell_wire[339];							inform_R[340][1] = r_cell_wire[340];							inform_R[341][1] = r_cell_wire[341];							inform_R[342][1] = r_cell_wire[342];							inform_R[343][1] = r_cell_wire[343];							inform_R[344][1] = r_cell_wire[344];							inform_R[345][1] = r_cell_wire[345];							inform_R[346][1] = r_cell_wire[346];							inform_R[347][1] = r_cell_wire[347];							inform_R[348][1] = r_cell_wire[348];							inform_R[349][1] = r_cell_wire[349];							inform_R[350][1] = r_cell_wire[350];							inform_R[351][1] = r_cell_wire[351];							inform_R[352][1] = r_cell_wire[352];							inform_R[353][1] = r_cell_wire[353];							inform_R[354][1] = r_cell_wire[354];							inform_R[355][1] = r_cell_wire[355];							inform_R[356][1] = r_cell_wire[356];							inform_R[357][1] = r_cell_wire[357];							inform_R[358][1] = r_cell_wire[358];							inform_R[359][1] = r_cell_wire[359];							inform_R[360][1] = r_cell_wire[360];							inform_R[361][1] = r_cell_wire[361];							inform_R[362][1] = r_cell_wire[362];							inform_R[363][1] = r_cell_wire[363];							inform_R[364][1] = r_cell_wire[364];							inform_R[365][1] = r_cell_wire[365];							inform_R[366][1] = r_cell_wire[366];							inform_R[367][1] = r_cell_wire[367];							inform_R[368][1] = r_cell_wire[368];							inform_R[369][1] = r_cell_wire[369];							inform_R[370][1] = r_cell_wire[370];							inform_R[371][1] = r_cell_wire[371];							inform_R[372][1] = r_cell_wire[372];							inform_R[373][1] = r_cell_wire[373];							inform_R[374][1] = r_cell_wire[374];							inform_R[375][1] = r_cell_wire[375];							inform_R[376][1] = r_cell_wire[376];							inform_R[377][1] = r_cell_wire[377];							inform_R[378][1] = r_cell_wire[378];							inform_R[379][1] = r_cell_wire[379];							inform_R[380][1] = r_cell_wire[380];							inform_R[381][1] = r_cell_wire[381];							inform_R[382][1] = r_cell_wire[382];							inform_R[383][1] = r_cell_wire[383];							inform_R[384][1] = r_cell_wire[384];							inform_R[385][1] = r_cell_wire[385];							inform_R[386][1] = r_cell_wire[386];							inform_R[387][1] = r_cell_wire[387];							inform_R[388][1] = r_cell_wire[388];							inform_R[389][1] = r_cell_wire[389];							inform_R[390][1] = r_cell_wire[390];							inform_R[391][1] = r_cell_wire[391];							inform_R[392][1] = r_cell_wire[392];							inform_R[393][1] = r_cell_wire[393];							inform_R[394][1] = r_cell_wire[394];							inform_R[395][1] = r_cell_wire[395];							inform_R[396][1] = r_cell_wire[396];							inform_R[397][1] = r_cell_wire[397];							inform_R[398][1] = r_cell_wire[398];							inform_R[399][1] = r_cell_wire[399];							inform_R[400][1] = r_cell_wire[400];							inform_R[401][1] = r_cell_wire[401];							inform_R[402][1] = r_cell_wire[402];							inform_R[403][1] = r_cell_wire[403];							inform_R[404][1] = r_cell_wire[404];							inform_R[405][1] = r_cell_wire[405];							inform_R[406][1] = r_cell_wire[406];							inform_R[407][1] = r_cell_wire[407];							inform_R[408][1] = r_cell_wire[408];							inform_R[409][1] = r_cell_wire[409];							inform_R[410][1] = r_cell_wire[410];							inform_R[411][1] = r_cell_wire[411];							inform_R[412][1] = r_cell_wire[412];							inform_R[413][1] = r_cell_wire[413];							inform_R[414][1] = r_cell_wire[414];							inform_R[415][1] = r_cell_wire[415];							inform_R[416][1] = r_cell_wire[416];							inform_R[417][1] = r_cell_wire[417];							inform_R[418][1] = r_cell_wire[418];							inform_R[419][1] = r_cell_wire[419];							inform_R[420][1] = r_cell_wire[420];							inform_R[421][1] = r_cell_wire[421];							inform_R[422][1] = r_cell_wire[422];							inform_R[423][1] = r_cell_wire[423];							inform_R[424][1] = r_cell_wire[424];							inform_R[425][1] = r_cell_wire[425];							inform_R[426][1] = r_cell_wire[426];							inform_R[427][1] = r_cell_wire[427];							inform_R[428][1] = r_cell_wire[428];							inform_R[429][1] = r_cell_wire[429];							inform_R[430][1] = r_cell_wire[430];							inform_R[431][1] = r_cell_wire[431];							inform_R[432][1] = r_cell_wire[432];							inform_R[433][1] = r_cell_wire[433];							inform_R[434][1] = r_cell_wire[434];							inform_R[435][1] = r_cell_wire[435];							inform_R[436][1] = r_cell_wire[436];							inform_R[437][1] = r_cell_wire[437];							inform_R[438][1] = r_cell_wire[438];							inform_R[439][1] = r_cell_wire[439];							inform_R[440][1] = r_cell_wire[440];							inform_R[441][1] = r_cell_wire[441];							inform_R[442][1] = r_cell_wire[442];							inform_R[443][1] = r_cell_wire[443];							inform_R[444][1] = r_cell_wire[444];							inform_R[445][1] = r_cell_wire[445];							inform_R[446][1] = r_cell_wire[446];							inform_R[447][1] = r_cell_wire[447];							inform_R[448][1] = r_cell_wire[448];							inform_R[449][1] = r_cell_wire[449];							inform_R[450][1] = r_cell_wire[450];							inform_R[451][1] = r_cell_wire[451];							inform_R[452][1] = r_cell_wire[452];							inform_R[453][1] = r_cell_wire[453];							inform_R[454][1] = r_cell_wire[454];							inform_R[455][1] = r_cell_wire[455];							inform_R[456][1] = r_cell_wire[456];							inform_R[457][1] = r_cell_wire[457];							inform_R[458][1] = r_cell_wire[458];							inform_R[459][1] = r_cell_wire[459];							inform_R[460][1] = r_cell_wire[460];							inform_R[461][1] = r_cell_wire[461];							inform_R[462][1] = r_cell_wire[462];							inform_R[463][1] = r_cell_wire[463];							inform_R[464][1] = r_cell_wire[464];							inform_R[465][1] = r_cell_wire[465];							inform_R[466][1] = r_cell_wire[466];							inform_R[467][1] = r_cell_wire[467];							inform_R[468][1] = r_cell_wire[468];							inform_R[469][1] = r_cell_wire[469];							inform_R[470][1] = r_cell_wire[470];							inform_R[471][1] = r_cell_wire[471];							inform_R[472][1] = r_cell_wire[472];							inform_R[473][1] = r_cell_wire[473];							inform_R[474][1] = r_cell_wire[474];							inform_R[475][1] = r_cell_wire[475];							inform_R[476][1] = r_cell_wire[476];							inform_R[477][1] = r_cell_wire[477];							inform_R[478][1] = r_cell_wire[478];							inform_R[479][1] = r_cell_wire[479];							inform_R[480][1] = r_cell_wire[480];							inform_R[481][1] = r_cell_wire[481];							inform_R[482][1] = r_cell_wire[482];							inform_R[483][1] = r_cell_wire[483];							inform_R[484][1] = r_cell_wire[484];							inform_R[485][1] = r_cell_wire[485];							inform_R[486][1] = r_cell_wire[486];							inform_R[487][1] = r_cell_wire[487];							inform_R[488][1] = r_cell_wire[488];							inform_R[489][1] = r_cell_wire[489];							inform_R[490][1] = r_cell_wire[490];							inform_R[491][1] = r_cell_wire[491];							inform_R[492][1] = r_cell_wire[492];							inform_R[493][1] = r_cell_wire[493];							inform_R[494][1] = r_cell_wire[494];							inform_R[495][1] = r_cell_wire[495];							inform_R[496][1] = r_cell_wire[496];							inform_R[497][1] = r_cell_wire[497];							inform_R[498][1] = r_cell_wire[498];							inform_R[499][1] = r_cell_wire[499];							inform_R[500][1] = r_cell_wire[500];							inform_R[501][1] = r_cell_wire[501];							inform_R[502][1] = r_cell_wire[502];							inform_R[503][1] = r_cell_wire[503];							inform_R[504][1] = r_cell_wire[504];							inform_R[505][1] = r_cell_wire[505];							inform_R[506][1] = r_cell_wire[506];							inform_R[507][1] = r_cell_wire[507];							inform_R[508][1] = r_cell_wire[508];							inform_R[509][1] = r_cell_wire[509];							inform_R[510][1] = r_cell_wire[510];							inform_R[511][1] = r_cell_wire[511];							inform_R[512][1] = r_cell_wire[512];							inform_R[513][1] = r_cell_wire[513];							inform_R[514][1] = r_cell_wire[514];							inform_R[515][1] = r_cell_wire[515];							inform_R[516][1] = r_cell_wire[516];							inform_R[517][1] = r_cell_wire[517];							inform_R[518][1] = r_cell_wire[518];							inform_R[519][1] = r_cell_wire[519];							inform_R[520][1] = r_cell_wire[520];							inform_R[521][1] = r_cell_wire[521];							inform_R[522][1] = r_cell_wire[522];							inform_R[523][1] = r_cell_wire[523];							inform_R[524][1] = r_cell_wire[524];							inform_R[525][1] = r_cell_wire[525];							inform_R[526][1] = r_cell_wire[526];							inform_R[527][1] = r_cell_wire[527];							inform_R[528][1] = r_cell_wire[528];							inform_R[529][1] = r_cell_wire[529];							inform_R[530][1] = r_cell_wire[530];							inform_R[531][1] = r_cell_wire[531];							inform_R[532][1] = r_cell_wire[532];							inform_R[533][1] = r_cell_wire[533];							inform_R[534][1] = r_cell_wire[534];							inform_R[535][1] = r_cell_wire[535];							inform_R[536][1] = r_cell_wire[536];							inform_R[537][1] = r_cell_wire[537];							inform_R[538][1] = r_cell_wire[538];							inform_R[539][1] = r_cell_wire[539];							inform_R[540][1] = r_cell_wire[540];							inform_R[541][1] = r_cell_wire[541];							inform_R[542][1] = r_cell_wire[542];							inform_R[543][1] = r_cell_wire[543];							inform_R[544][1] = r_cell_wire[544];							inform_R[545][1] = r_cell_wire[545];							inform_R[546][1] = r_cell_wire[546];							inform_R[547][1] = r_cell_wire[547];							inform_R[548][1] = r_cell_wire[548];							inform_R[549][1] = r_cell_wire[549];							inform_R[550][1] = r_cell_wire[550];							inform_R[551][1] = r_cell_wire[551];							inform_R[552][1] = r_cell_wire[552];							inform_R[553][1] = r_cell_wire[553];							inform_R[554][1] = r_cell_wire[554];							inform_R[555][1] = r_cell_wire[555];							inform_R[556][1] = r_cell_wire[556];							inform_R[557][1] = r_cell_wire[557];							inform_R[558][1] = r_cell_wire[558];							inform_R[559][1] = r_cell_wire[559];							inform_R[560][1] = r_cell_wire[560];							inform_R[561][1] = r_cell_wire[561];							inform_R[562][1] = r_cell_wire[562];							inform_R[563][1] = r_cell_wire[563];							inform_R[564][1] = r_cell_wire[564];							inform_R[565][1] = r_cell_wire[565];							inform_R[566][1] = r_cell_wire[566];							inform_R[567][1] = r_cell_wire[567];							inform_R[568][1] = r_cell_wire[568];							inform_R[569][1] = r_cell_wire[569];							inform_R[570][1] = r_cell_wire[570];							inform_R[571][1] = r_cell_wire[571];							inform_R[572][1] = r_cell_wire[572];							inform_R[573][1] = r_cell_wire[573];							inform_R[574][1] = r_cell_wire[574];							inform_R[575][1] = r_cell_wire[575];							inform_R[576][1] = r_cell_wire[576];							inform_R[577][1] = r_cell_wire[577];							inform_R[578][1] = r_cell_wire[578];							inform_R[579][1] = r_cell_wire[579];							inform_R[580][1] = r_cell_wire[580];							inform_R[581][1] = r_cell_wire[581];							inform_R[582][1] = r_cell_wire[582];							inform_R[583][1] = r_cell_wire[583];							inform_R[584][1] = r_cell_wire[584];							inform_R[585][1] = r_cell_wire[585];							inform_R[586][1] = r_cell_wire[586];							inform_R[587][1] = r_cell_wire[587];							inform_R[588][1] = r_cell_wire[588];							inform_R[589][1] = r_cell_wire[589];							inform_R[590][1] = r_cell_wire[590];							inform_R[591][1] = r_cell_wire[591];							inform_R[592][1] = r_cell_wire[592];							inform_R[593][1] = r_cell_wire[593];							inform_R[594][1] = r_cell_wire[594];							inform_R[595][1] = r_cell_wire[595];							inform_R[596][1] = r_cell_wire[596];							inform_R[597][1] = r_cell_wire[597];							inform_R[598][1] = r_cell_wire[598];							inform_R[599][1] = r_cell_wire[599];							inform_R[600][1] = r_cell_wire[600];							inform_R[601][1] = r_cell_wire[601];							inform_R[602][1] = r_cell_wire[602];							inform_R[603][1] = r_cell_wire[603];							inform_R[604][1] = r_cell_wire[604];							inform_R[605][1] = r_cell_wire[605];							inform_R[606][1] = r_cell_wire[606];							inform_R[607][1] = r_cell_wire[607];							inform_R[608][1] = r_cell_wire[608];							inform_R[609][1] = r_cell_wire[609];							inform_R[610][1] = r_cell_wire[610];							inform_R[611][1] = r_cell_wire[611];							inform_R[612][1] = r_cell_wire[612];							inform_R[613][1] = r_cell_wire[613];							inform_R[614][1] = r_cell_wire[614];							inform_R[615][1] = r_cell_wire[615];							inform_R[616][1] = r_cell_wire[616];							inform_R[617][1] = r_cell_wire[617];							inform_R[618][1] = r_cell_wire[618];							inform_R[619][1] = r_cell_wire[619];							inform_R[620][1] = r_cell_wire[620];							inform_R[621][1] = r_cell_wire[621];							inform_R[622][1] = r_cell_wire[622];							inform_R[623][1] = r_cell_wire[623];							inform_R[624][1] = r_cell_wire[624];							inform_R[625][1] = r_cell_wire[625];							inform_R[626][1] = r_cell_wire[626];							inform_R[627][1] = r_cell_wire[627];							inform_R[628][1] = r_cell_wire[628];							inform_R[629][1] = r_cell_wire[629];							inform_R[630][1] = r_cell_wire[630];							inform_R[631][1] = r_cell_wire[631];							inform_R[632][1] = r_cell_wire[632];							inform_R[633][1] = r_cell_wire[633];							inform_R[634][1] = r_cell_wire[634];							inform_R[635][1] = r_cell_wire[635];							inform_R[636][1] = r_cell_wire[636];							inform_R[637][1] = r_cell_wire[637];							inform_R[638][1] = r_cell_wire[638];							inform_R[639][1] = r_cell_wire[639];							inform_R[640][1] = r_cell_wire[640];							inform_R[641][1] = r_cell_wire[641];							inform_R[642][1] = r_cell_wire[642];							inform_R[643][1] = r_cell_wire[643];							inform_R[644][1] = r_cell_wire[644];							inform_R[645][1] = r_cell_wire[645];							inform_R[646][1] = r_cell_wire[646];							inform_R[647][1] = r_cell_wire[647];							inform_R[648][1] = r_cell_wire[648];							inform_R[649][1] = r_cell_wire[649];							inform_R[650][1] = r_cell_wire[650];							inform_R[651][1] = r_cell_wire[651];							inform_R[652][1] = r_cell_wire[652];							inform_R[653][1] = r_cell_wire[653];							inform_R[654][1] = r_cell_wire[654];							inform_R[655][1] = r_cell_wire[655];							inform_R[656][1] = r_cell_wire[656];							inform_R[657][1] = r_cell_wire[657];							inform_R[658][1] = r_cell_wire[658];							inform_R[659][1] = r_cell_wire[659];							inform_R[660][1] = r_cell_wire[660];							inform_R[661][1] = r_cell_wire[661];							inform_R[662][1] = r_cell_wire[662];							inform_R[663][1] = r_cell_wire[663];							inform_R[664][1] = r_cell_wire[664];							inform_R[665][1] = r_cell_wire[665];							inform_R[666][1] = r_cell_wire[666];							inform_R[667][1] = r_cell_wire[667];							inform_R[668][1] = r_cell_wire[668];							inform_R[669][1] = r_cell_wire[669];							inform_R[670][1] = r_cell_wire[670];							inform_R[671][1] = r_cell_wire[671];							inform_R[672][1] = r_cell_wire[672];							inform_R[673][1] = r_cell_wire[673];							inform_R[674][1] = r_cell_wire[674];							inform_R[675][1] = r_cell_wire[675];							inform_R[676][1] = r_cell_wire[676];							inform_R[677][1] = r_cell_wire[677];							inform_R[678][1] = r_cell_wire[678];							inform_R[679][1] = r_cell_wire[679];							inform_R[680][1] = r_cell_wire[680];							inform_R[681][1] = r_cell_wire[681];							inform_R[682][1] = r_cell_wire[682];							inform_R[683][1] = r_cell_wire[683];							inform_R[684][1] = r_cell_wire[684];							inform_R[685][1] = r_cell_wire[685];							inform_R[686][1] = r_cell_wire[686];							inform_R[687][1] = r_cell_wire[687];							inform_R[688][1] = r_cell_wire[688];							inform_R[689][1] = r_cell_wire[689];							inform_R[690][1] = r_cell_wire[690];							inform_R[691][1] = r_cell_wire[691];							inform_R[692][1] = r_cell_wire[692];							inform_R[693][1] = r_cell_wire[693];							inform_R[694][1] = r_cell_wire[694];							inform_R[695][1] = r_cell_wire[695];							inform_R[696][1] = r_cell_wire[696];							inform_R[697][1] = r_cell_wire[697];							inform_R[698][1] = r_cell_wire[698];							inform_R[699][1] = r_cell_wire[699];							inform_R[700][1] = r_cell_wire[700];							inform_R[701][1] = r_cell_wire[701];							inform_R[702][1] = r_cell_wire[702];							inform_R[703][1] = r_cell_wire[703];							inform_R[704][1] = r_cell_wire[704];							inform_R[705][1] = r_cell_wire[705];							inform_R[706][1] = r_cell_wire[706];							inform_R[707][1] = r_cell_wire[707];							inform_R[708][1] = r_cell_wire[708];							inform_R[709][1] = r_cell_wire[709];							inform_R[710][1] = r_cell_wire[710];							inform_R[711][1] = r_cell_wire[711];							inform_R[712][1] = r_cell_wire[712];							inform_R[713][1] = r_cell_wire[713];							inform_R[714][1] = r_cell_wire[714];							inform_R[715][1] = r_cell_wire[715];							inform_R[716][1] = r_cell_wire[716];							inform_R[717][1] = r_cell_wire[717];							inform_R[718][1] = r_cell_wire[718];							inform_R[719][1] = r_cell_wire[719];							inform_R[720][1] = r_cell_wire[720];							inform_R[721][1] = r_cell_wire[721];							inform_R[722][1] = r_cell_wire[722];							inform_R[723][1] = r_cell_wire[723];							inform_R[724][1] = r_cell_wire[724];							inform_R[725][1] = r_cell_wire[725];							inform_R[726][1] = r_cell_wire[726];							inform_R[727][1] = r_cell_wire[727];							inform_R[728][1] = r_cell_wire[728];							inform_R[729][1] = r_cell_wire[729];							inform_R[730][1] = r_cell_wire[730];							inform_R[731][1] = r_cell_wire[731];							inform_R[732][1] = r_cell_wire[732];							inform_R[733][1] = r_cell_wire[733];							inform_R[734][1] = r_cell_wire[734];							inform_R[735][1] = r_cell_wire[735];							inform_R[736][1] = r_cell_wire[736];							inform_R[737][1] = r_cell_wire[737];							inform_R[738][1] = r_cell_wire[738];							inform_R[739][1] = r_cell_wire[739];							inform_R[740][1] = r_cell_wire[740];							inform_R[741][1] = r_cell_wire[741];							inform_R[742][1] = r_cell_wire[742];							inform_R[743][1] = r_cell_wire[743];							inform_R[744][1] = r_cell_wire[744];							inform_R[745][1] = r_cell_wire[745];							inform_R[746][1] = r_cell_wire[746];							inform_R[747][1] = r_cell_wire[747];							inform_R[748][1] = r_cell_wire[748];							inform_R[749][1] = r_cell_wire[749];							inform_R[750][1] = r_cell_wire[750];							inform_R[751][1] = r_cell_wire[751];							inform_R[752][1] = r_cell_wire[752];							inform_R[753][1] = r_cell_wire[753];							inform_R[754][1] = r_cell_wire[754];							inform_R[755][1] = r_cell_wire[755];							inform_R[756][1] = r_cell_wire[756];							inform_R[757][1] = r_cell_wire[757];							inform_R[758][1] = r_cell_wire[758];							inform_R[759][1] = r_cell_wire[759];							inform_R[760][1] = r_cell_wire[760];							inform_R[761][1] = r_cell_wire[761];							inform_R[762][1] = r_cell_wire[762];							inform_R[763][1] = r_cell_wire[763];							inform_R[764][1] = r_cell_wire[764];							inform_R[765][1] = r_cell_wire[765];							inform_R[766][1] = r_cell_wire[766];							inform_R[767][1] = r_cell_wire[767];							inform_R[768][1] = r_cell_wire[768];							inform_R[769][1] = r_cell_wire[769];							inform_R[770][1] = r_cell_wire[770];							inform_R[771][1] = r_cell_wire[771];							inform_R[772][1] = r_cell_wire[772];							inform_R[773][1] = r_cell_wire[773];							inform_R[774][1] = r_cell_wire[774];							inform_R[775][1] = r_cell_wire[775];							inform_R[776][1] = r_cell_wire[776];							inform_R[777][1] = r_cell_wire[777];							inform_R[778][1] = r_cell_wire[778];							inform_R[779][1] = r_cell_wire[779];							inform_R[780][1] = r_cell_wire[780];							inform_R[781][1] = r_cell_wire[781];							inform_R[782][1] = r_cell_wire[782];							inform_R[783][1] = r_cell_wire[783];							inform_R[784][1] = r_cell_wire[784];							inform_R[785][1] = r_cell_wire[785];							inform_R[786][1] = r_cell_wire[786];							inform_R[787][1] = r_cell_wire[787];							inform_R[788][1] = r_cell_wire[788];							inform_R[789][1] = r_cell_wire[789];							inform_R[790][1] = r_cell_wire[790];							inform_R[791][1] = r_cell_wire[791];							inform_R[792][1] = r_cell_wire[792];							inform_R[793][1] = r_cell_wire[793];							inform_R[794][1] = r_cell_wire[794];							inform_R[795][1] = r_cell_wire[795];							inform_R[796][1] = r_cell_wire[796];							inform_R[797][1] = r_cell_wire[797];							inform_R[798][1] = r_cell_wire[798];							inform_R[799][1] = r_cell_wire[799];							inform_R[800][1] = r_cell_wire[800];							inform_R[801][1] = r_cell_wire[801];							inform_R[802][1] = r_cell_wire[802];							inform_R[803][1] = r_cell_wire[803];							inform_R[804][1] = r_cell_wire[804];							inform_R[805][1] = r_cell_wire[805];							inform_R[806][1] = r_cell_wire[806];							inform_R[807][1] = r_cell_wire[807];							inform_R[808][1] = r_cell_wire[808];							inform_R[809][1] = r_cell_wire[809];							inform_R[810][1] = r_cell_wire[810];							inform_R[811][1] = r_cell_wire[811];							inform_R[812][1] = r_cell_wire[812];							inform_R[813][1] = r_cell_wire[813];							inform_R[814][1] = r_cell_wire[814];							inform_R[815][1] = r_cell_wire[815];							inform_R[816][1] = r_cell_wire[816];							inform_R[817][1] = r_cell_wire[817];							inform_R[818][1] = r_cell_wire[818];							inform_R[819][1] = r_cell_wire[819];							inform_R[820][1] = r_cell_wire[820];							inform_R[821][1] = r_cell_wire[821];							inform_R[822][1] = r_cell_wire[822];							inform_R[823][1] = r_cell_wire[823];							inform_R[824][1] = r_cell_wire[824];							inform_R[825][1] = r_cell_wire[825];							inform_R[826][1] = r_cell_wire[826];							inform_R[827][1] = r_cell_wire[827];							inform_R[828][1] = r_cell_wire[828];							inform_R[829][1] = r_cell_wire[829];							inform_R[830][1] = r_cell_wire[830];							inform_R[831][1] = r_cell_wire[831];							inform_R[832][1] = r_cell_wire[832];							inform_R[833][1] = r_cell_wire[833];							inform_R[834][1] = r_cell_wire[834];							inform_R[835][1] = r_cell_wire[835];							inform_R[836][1] = r_cell_wire[836];							inform_R[837][1] = r_cell_wire[837];							inform_R[838][1] = r_cell_wire[838];							inform_R[839][1] = r_cell_wire[839];							inform_R[840][1] = r_cell_wire[840];							inform_R[841][1] = r_cell_wire[841];							inform_R[842][1] = r_cell_wire[842];							inform_R[843][1] = r_cell_wire[843];							inform_R[844][1] = r_cell_wire[844];							inform_R[845][1] = r_cell_wire[845];							inform_R[846][1] = r_cell_wire[846];							inform_R[847][1] = r_cell_wire[847];							inform_R[848][1] = r_cell_wire[848];							inform_R[849][1] = r_cell_wire[849];							inform_R[850][1] = r_cell_wire[850];							inform_R[851][1] = r_cell_wire[851];							inform_R[852][1] = r_cell_wire[852];							inform_R[853][1] = r_cell_wire[853];							inform_R[854][1] = r_cell_wire[854];							inform_R[855][1] = r_cell_wire[855];							inform_R[856][1] = r_cell_wire[856];							inform_R[857][1] = r_cell_wire[857];							inform_R[858][1] = r_cell_wire[858];							inform_R[859][1] = r_cell_wire[859];							inform_R[860][1] = r_cell_wire[860];							inform_R[861][1] = r_cell_wire[861];							inform_R[862][1] = r_cell_wire[862];							inform_R[863][1] = r_cell_wire[863];							inform_R[864][1] = r_cell_wire[864];							inform_R[865][1] = r_cell_wire[865];							inform_R[866][1] = r_cell_wire[866];							inform_R[867][1] = r_cell_wire[867];							inform_R[868][1] = r_cell_wire[868];							inform_R[869][1] = r_cell_wire[869];							inform_R[870][1] = r_cell_wire[870];							inform_R[871][1] = r_cell_wire[871];							inform_R[872][1] = r_cell_wire[872];							inform_R[873][1] = r_cell_wire[873];							inform_R[874][1] = r_cell_wire[874];							inform_R[875][1] = r_cell_wire[875];							inform_R[876][1] = r_cell_wire[876];							inform_R[877][1] = r_cell_wire[877];							inform_R[878][1] = r_cell_wire[878];							inform_R[879][1] = r_cell_wire[879];							inform_R[880][1] = r_cell_wire[880];							inform_R[881][1] = r_cell_wire[881];							inform_R[882][1] = r_cell_wire[882];							inform_R[883][1] = r_cell_wire[883];							inform_R[884][1] = r_cell_wire[884];							inform_R[885][1] = r_cell_wire[885];							inform_R[886][1] = r_cell_wire[886];							inform_R[887][1] = r_cell_wire[887];							inform_R[888][1] = r_cell_wire[888];							inform_R[889][1] = r_cell_wire[889];							inform_R[890][1] = r_cell_wire[890];							inform_R[891][1] = r_cell_wire[891];							inform_R[892][1] = r_cell_wire[892];							inform_R[893][1] = r_cell_wire[893];							inform_R[894][1] = r_cell_wire[894];							inform_R[895][1] = r_cell_wire[895];							inform_R[896][1] = r_cell_wire[896];							inform_R[897][1] = r_cell_wire[897];							inform_R[898][1] = r_cell_wire[898];							inform_R[899][1] = r_cell_wire[899];							inform_R[900][1] = r_cell_wire[900];							inform_R[901][1] = r_cell_wire[901];							inform_R[902][1] = r_cell_wire[902];							inform_R[903][1] = r_cell_wire[903];							inform_R[904][1] = r_cell_wire[904];							inform_R[905][1] = r_cell_wire[905];							inform_R[906][1] = r_cell_wire[906];							inform_R[907][1] = r_cell_wire[907];							inform_R[908][1] = r_cell_wire[908];							inform_R[909][1] = r_cell_wire[909];							inform_R[910][1] = r_cell_wire[910];							inform_R[911][1] = r_cell_wire[911];							inform_R[912][1] = r_cell_wire[912];							inform_R[913][1] = r_cell_wire[913];							inform_R[914][1] = r_cell_wire[914];							inform_R[915][1] = r_cell_wire[915];							inform_R[916][1] = r_cell_wire[916];							inform_R[917][1] = r_cell_wire[917];							inform_R[918][1] = r_cell_wire[918];							inform_R[919][1] = r_cell_wire[919];							inform_R[920][1] = r_cell_wire[920];							inform_R[921][1] = r_cell_wire[921];							inform_R[922][1] = r_cell_wire[922];							inform_R[923][1] = r_cell_wire[923];							inform_R[924][1] = r_cell_wire[924];							inform_R[925][1] = r_cell_wire[925];							inform_R[926][1] = r_cell_wire[926];							inform_R[927][1] = r_cell_wire[927];							inform_R[928][1] = r_cell_wire[928];							inform_R[929][1] = r_cell_wire[929];							inform_R[930][1] = r_cell_wire[930];							inform_R[931][1] = r_cell_wire[931];							inform_R[932][1] = r_cell_wire[932];							inform_R[933][1] = r_cell_wire[933];							inform_R[934][1] = r_cell_wire[934];							inform_R[935][1] = r_cell_wire[935];							inform_R[936][1] = r_cell_wire[936];							inform_R[937][1] = r_cell_wire[937];							inform_R[938][1] = r_cell_wire[938];							inform_R[939][1] = r_cell_wire[939];							inform_R[940][1] = r_cell_wire[940];							inform_R[941][1] = r_cell_wire[941];							inform_R[942][1] = r_cell_wire[942];							inform_R[943][1] = r_cell_wire[943];							inform_R[944][1] = r_cell_wire[944];							inform_R[945][1] = r_cell_wire[945];							inform_R[946][1] = r_cell_wire[946];							inform_R[947][1] = r_cell_wire[947];							inform_R[948][1] = r_cell_wire[948];							inform_R[949][1] = r_cell_wire[949];							inform_R[950][1] = r_cell_wire[950];							inform_R[951][1] = r_cell_wire[951];							inform_R[952][1] = r_cell_wire[952];							inform_R[953][1] = r_cell_wire[953];							inform_R[954][1] = r_cell_wire[954];							inform_R[955][1] = r_cell_wire[955];							inform_R[956][1] = r_cell_wire[956];							inform_R[957][1] = r_cell_wire[957];							inform_R[958][1] = r_cell_wire[958];							inform_R[959][1] = r_cell_wire[959];							inform_R[960][1] = r_cell_wire[960];							inform_R[961][1] = r_cell_wire[961];							inform_R[962][1] = r_cell_wire[962];							inform_R[963][1] = r_cell_wire[963];							inform_R[964][1] = r_cell_wire[964];							inform_R[965][1] = r_cell_wire[965];							inform_R[966][1] = r_cell_wire[966];							inform_R[967][1] = r_cell_wire[967];							inform_R[968][1] = r_cell_wire[968];							inform_R[969][1] = r_cell_wire[969];							inform_R[970][1] = r_cell_wire[970];							inform_R[971][1] = r_cell_wire[971];							inform_R[972][1] = r_cell_wire[972];							inform_R[973][1] = r_cell_wire[973];							inform_R[974][1] = r_cell_wire[974];							inform_R[975][1] = r_cell_wire[975];							inform_R[976][1] = r_cell_wire[976];							inform_R[977][1] = r_cell_wire[977];							inform_R[978][1] = r_cell_wire[978];							inform_R[979][1] = r_cell_wire[979];							inform_R[980][1] = r_cell_wire[980];							inform_R[981][1] = r_cell_wire[981];							inform_R[982][1] = r_cell_wire[982];							inform_R[983][1] = r_cell_wire[983];							inform_R[984][1] = r_cell_wire[984];							inform_R[985][1] = r_cell_wire[985];							inform_R[986][1] = r_cell_wire[986];							inform_R[987][1] = r_cell_wire[987];							inform_R[988][1] = r_cell_wire[988];							inform_R[989][1] = r_cell_wire[989];							inform_R[990][1] = r_cell_wire[990];							inform_R[991][1] = r_cell_wire[991];							inform_R[992][1] = r_cell_wire[992];							inform_R[993][1] = r_cell_wire[993];							inform_R[994][1] = r_cell_wire[994];							inform_R[995][1] = r_cell_wire[995];							inform_R[996][1] = r_cell_wire[996];							inform_R[997][1] = r_cell_wire[997];							inform_R[998][1] = r_cell_wire[998];							inform_R[999][1] = r_cell_wire[999];							inform_R[1000][1] = r_cell_wire[1000];							inform_R[1001][1] = r_cell_wire[1001];							inform_R[1002][1] = r_cell_wire[1002];							inform_R[1003][1] = r_cell_wire[1003];							inform_R[1004][1] = r_cell_wire[1004];							inform_R[1005][1] = r_cell_wire[1005];							inform_R[1006][1] = r_cell_wire[1006];							inform_R[1007][1] = r_cell_wire[1007];							inform_R[1008][1] = r_cell_wire[1008];							inform_R[1009][1] = r_cell_wire[1009];							inform_R[1010][1] = r_cell_wire[1010];							inform_R[1011][1] = r_cell_wire[1011];							inform_R[1012][1] = r_cell_wire[1012];							inform_R[1013][1] = r_cell_wire[1013];							inform_R[1014][1] = r_cell_wire[1014];							inform_R[1015][1] = r_cell_wire[1015];							inform_R[1016][1] = r_cell_wire[1016];							inform_R[1017][1] = r_cell_wire[1017];							inform_R[1018][1] = r_cell_wire[1018];							inform_R[1019][1] = r_cell_wire[1019];							inform_R[1020][1] = r_cell_wire[1020];							inform_R[1021][1] = r_cell_wire[1021];							inform_R[1022][1] = r_cell_wire[1022];							inform_R[1023][1] = r_cell_wire[1023];							inform_L[0][0] = l_cell_wire[0];							inform_L[1][0] = l_cell_wire[1];							inform_L[2][0] = l_cell_wire[2];							inform_L[3][0] = l_cell_wire[3];							inform_L[4][0] = l_cell_wire[4];							inform_L[5][0] = l_cell_wire[5];							inform_L[6][0] = l_cell_wire[6];							inform_L[7][0] = l_cell_wire[7];							inform_L[8][0] = l_cell_wire[8];							inform_L[9][0] = l_cell_wire[9];							inform_L[10][0] = l_cell_wire[10];							inform_L[11][0] = l_cell_wire[11];							inform_L[12][0] = l_cell_wire[12];							inform_L[13][0] = l_cell_wire[13];							inform_L[14][0] = l_cell_wire[14];							inform_L[15][0] = l_cell_wire[15];							inform_L[16][0] = l_cell_wire[16];							inform_L[17][0] = l_cell_wire[17];							inform_L[18][0] = l_cell_wire[18];							inform_L[19][0] = l_cell_wire[19];							inform_L[20][0] = l_cell_wire[20];							inform_L[21][0] = l_cell_wire[21];							inform_L[22][0] = l_cell_wire[22];							inform_L[23][0] = l_cell_wire[23];							inform_L[24][0] = l_cell_wire[24];							inform_L[25][0] = l_cell_wire[25];							inform_L[26][0] = l_cell_wire[26];							inform_L[27][0] = l_cell_wire[27];							inform_L[28][0] = l_cell_wire[28];							inform_L[29][0] = l_cell_wire[29];							inform_L[30][0] = l_cell_wire[30];							inform_L[31][0] = l_cell_wire[31];							inform_L[32][0] = l_cell_wire[32];							inform_L[33][0] = l_cell_wire[33];							inform_L[34][0] = l_cell_wire[34];							inform_L[35][0] = l_cell_wire[35];							inform_L[36][0] = l_cell_wire[36];							inform_L[37][0] = l_cell_wire[37];							inform_L[38][0] = l_cell_wire[38];							inform_L[39][0] = l_cell_wire[39];							inform_L[40][0] = l_cell_wire[40];							inform_L[41][0] = l_cell_wire[41];							inform_L[42][0] = l_cell_wire[42];							inform_L[43][0] = l_cell_wire[43];							inform_L[44][0] = l_cell_wire[44];							inform_L[45][0] = l_cell_wire[45];							inform_L[46][0] = l_cell_wire[46];							inform_L[47][0] = l_cell_wire[47];							inform_L[48][0] = l_cell_wire[48];							inform_L[49][0] = l_cell_wire[49];							inform_L[50][0] = l_cell_wire[50];							inform_L[51][0] = l_cell_wire[51];							inform_L[52][0] = l_cell_wire[52];							inform_L[53][0] = l_cell_wire[53];							inform_L[54][0] = l_cell_wire[54];							inform_L[55][0] = l_cell_wire[55];							inform_L[56][0] = l_cell_wire[56];							inform_L[57][0] = l_cell_wire[57];							inform_L[58][0] = l_cell_wire[58];							inform_L[59][0] = l_cell_wire[59];							inform_L[60][0] = l_cell_wire[60];							inform_L[61][0] = l_cell_wire[61];							inform_L[62][0] = l_cell_wire[62];							inform_L[63][0] = l_cell_wire[63];							inform_L[64][0] = l_cell_wire[64];							inform_L[65][0] = l_cell_wire[65];							inform_L[66][0] = l_cell_wire[66];							inform_L[67][0] = l_cell_wire[67];							inform_L[68][0] = l_cell_wire[68];							inform_L[69][0] = l_cell_wire[69];							inform_L[70][0] = l_cell_wire[70];							inform_L[71][0] = l_cell_wire[71];							inform_L[72][0] = l_cell_wire[72];							inform_L[73][0] = l_cell_wire[73];							inform_L[74][0] = l_cell_wire[74];							inform_L[75][0] = l_cell_wire[75];							inform_L[76][0] = l_cell_wire[76];							inform_L[77][0] = l_cell_wire[77];							inform_L[78][0] = l_cell_wire[78];							inform_L[79][0] = l_cell_wire[79];							inform_L[80][0] = l_cell_wire[80];							inform_L[81][0] = l_cell_wire[81];							inform_L[82][0] = l_cell_wire[82];							inform_L[83][0] = l_cell_wire[83];							inform_L[84][0] = l_cell_wire[84];							inform_L[85][0] = l_cell_wire[85];							inform_L[86][0] = l_cell_wire[86];							inform_L[87][0] = l_cell_wire[87];							inform_L[88][0] = l_cell_wire[88];							inform_L[89][0] = l_cell_wire[89];							inform_L[90][0] = l_cell_wire[90];							inform_L[91][0] = l_cell_wire[91];							inform_L[92][0] = l_cell_wire[92];							inform_L[93][0] = l_cell_wire[93];							inform_L[94][0] = l_cell_wire[94];							inform_L[95][0] = l_cell_wire[95];							inform_L[96][0] = l_cell_wire[96];							inform_L[97][0] = l_cell_wire[97];							inform_L[98][0] = l_cell_wire[98];							inform_L[99][0] = l_cell_wire[99];							inform_L[100][0] = l_cell_wire[100];							inform_L[101][0] = l_cell_wire[101];							inform_L[102][0] = l_cell_wire[102];							inform_L[103][0] = l_cell_wire[103];							inform_L[104][0] = l_cell_wire[104];							inform_L[105][0] = l_cell_wire[105];							inform_L[106][0] = l_cell_wire[106];							inform_L[107][0] = l_cell_wire[107];							inform_L[108][0] = l_cell_wire[108];							inform_L[109][0] = l_cell_wire[109];							inform_L[110][0] = l_cell_wire[110];							inform_L[111][0] = l_cell_wire[111];							inform_L[112][0] = l_cell_wire[112];							inform_L[113][0] = l_cell_wire[113];							inform_L[114][0] = l_cell_wire[114];							inform_L[115][0] = l_cell_wire[115];							inform_L[116][0] = l_cell_wire[116];							inform_L[117][0] = l_cell_wire[117];							inform_L[118][0] = l_cell_wire[118];							inform_L[119][0] = l_cell_wire[119];							inform_L[120][0] = l_cell_wire[120];							inform_L[121][0] = l_cell_wire[121];							inform_L[122][0] = l_cell_wire[122];							inform_L[123][0] = l_cell_wire[123];							inform_L[124][0] = l_cell_wire[124];							inform_L[125][0] = l_cell_wire[125];							inform_L[126][0] = l_cell_wire[126];							inform_L[127][0] = l_cell_wire[127];							inform_L[128][0] = l_cell_wire[128];							inform_L[129][0] = l_cell_wire[129];							inform_L[130][0] = l_cell_wire[130];							inform_L[131][0] = l_cell_wire[131];							inform_L[132][0] = l_cell_wire[132];							inform_L[133][0] = l_cell_wire[133];							inform_L[134][0] = l_cell_wire[134];							inform_L[135][0] = l_cell_wire[135];							inform_L[136][0] = l_cell_wire[136];							inform_L[137][0] = l_cell_wire[137];							inform_L[138][0] = l_cell_wire[138];							inform_L[139][0] = l_cell_wire[139];							inform_L[140][0] = l_cell_wire[140];							inform_L[141][0] = l_cell_wire[141];							inform_L[142][0] = l_cell_wire[142];							inform_L[143][0] = l_cell_wire[143];							inform_L[144][0] = l_cell_wire[144];							inform_L[145][0] = l_cell_wire[145];							inform_L[146][0] = l_cell_wire[146];							inform_L[147][0] = l_cell_wire[147];							inform_L[148][0] = l_cell_wire[148];							inform_L[149][0] = l_cell_wire[149];							inform_L[150][0] = l_cell_wire[150];							inform_L[151][0] = l_cell_wire[151];							inform_L[152][0] = l_cell_wire[152];							inform_L[153][0] = l_cell_wire[153];							inform_L[154][0] = l_cell_wire[154];							inform_L[155][0] = l_cell_wire[155];							inform_L[156][0] = l_cell_wire[156];							inform_L[157][0] = l_cell_wire[157];							inform_L[158][0] = l_cell_wire[158];							inform_L[159][0] = l_cell_wire[159];							inform_L[160][0] = l_cell_wire[160];							inform_L[161][0] = l_cell_wire[161];							inform_L[162][0] = l_cell_wire[162];							inform_L[163][0] = l_cell_wire[163];							inform_L[164][0] = l_cell_wire[164];							inform_L[165][0] = l_cell_wire[165];							inform_L[166][0] = l_cell_wire[166];							inform_L[167][0] = l_cell_wire[167];							inform_L[168][0] = l_cell_wire[168];							inform_L[169][0] = l_cell_wire[169];							inform_L[170][0] = l_cell_wire[170];							inform_L[171][0] = l_cell_wire[171];							inform_L[172][0] = l_cell_wire[172];							inform_L[173][0] = l_cell_wire[173];							inform_L[174][0] = l_cell_wire[174];							inform_L[175][0] = l_cell_wire[175];							inform_L[176][0] = l_cell_wire[176];							inform_L[177][0] = l_cell_wire[177];							inform_L[178][0] = l_cell_wire[178];							inform_L[179][0] = l_cell_wire[179];							inform_L[180][0] = l_cell_wire[180];							inform_L[181][0] = l_cell_wire[181];							inform_L[182][0] = l_cell_wire[182];							inform_L[183][0] = l_cell_wire[183];							inform_L[184][0] = l_cell_wire[184];							inform_L[185][0] = l_cell_wire[185];							inform_L[186][0] = l_cell_wire[186];							inform_L[187][0] = l_cell_wire[187];							inform_L[188][0] = l_cell_wire[188];							inform_L[189][0] = l_cell_wire[189];							inform_L[190][0] = l_cell_wire[190];							inform_L[191][0] = l_cell_wire[191];							inform_L[192][0] = l_cell_wire[192];							inform_L[193][0] = l_cell_wire[193];							inform_L[194][0] = l_cell_wire[194];							inform_L[195][0] = l_cell_wire[195];							inform_L[196][0] = l_cell_wire[196];							inform_L[197][0] = l_cell_wire[197];							inform_L[198][0] = l_cell_wire[198];							inform_L[199][0] = l_cell_wire[199];							inform_L[200][0] = l_cell_wire[200];							inform_L[201][0] = l_cell_wire[201];							inform_L[202][0] = l_cell_wire[202];							inform_L[203][0] = l_cell_wire[203];							inform_L[204][0] = l_cell_wire[204];							inform_L[205][0] = l_cell_wire[205];							inform_L[206][0] = l_cell_wire[206];							inform_L[207][0] = l_cell_wire[207];							inform_L[208][0] = l_cell_wire[208];							inform_L[209][0] = l_cell_wire[209];							inform_L[210][0] = l_cell_wire[210];							inform_L[211][0] = l_cell_wire[211];							inform_L[212][0] = l_cell_wire[212];							inform_L[213][0] = l_cell_wire[213];							inform_L[214][0] = l_cell_wire[214];							inform_L[215][0] = l_cell_wire[215];							inform_L[216][0] = l_cell_wire[216];							inform_L[217][0] = l_cell_wire[217];							inform_L[218][0] = l_cell_wire[218];							inform_L[219][0] = l_cell_wire[219];							inform_L[220][0] = l_cell_wire[220];							inform_L[221][0] = l_cell_wire[221];							inform_L[222][0] = l_cell_wire[222];							inform_L[223][0] = l_cell_wire[223];							inform_L[224][0] = l_cell_wire[224];							inform_L[225][0] = l_cell_wire[225];							inform_L[226][0] = l_cell_wire[226];							inform_L[227][0] = l_cell_wire[227];							inform_L[228][0] = l_cell_wire[228];							inform_L[229][0] = l_cell_wire[229];							inform_L[230][0] = l_cell_wire[230];							inform_L[231][0] = l_cell_wire[231];							inform_L[232][0] = l_cell_wire[232];							inform_L[233][0] = l_cell_wire[233];							inform_L[234][0] = l_cell_wire[234];							inform_L[235][0] = l_cell_wire[235];							inform_L[236][0] = l_cell_wire[236];							inform_L[237][0] = l_cell_wire[237];							inform_L[238][0] = l_cell_wire[238];							inform_L[239][0] = l_cell_wire[239];							inform_L[240][0] = l_cell_wire[240];							inform_L[241][0] = l_cell_wire[241];							inform_L[242][0] = l_cell_wire[242];							inform_L[243][0] = l_cell_wire[243];							inform_L[244][0] = l_cell_wire[244];							inform_L[245][0] = l_cell_wire[245];							inform_L[246][0] = l_cell_wire[246];							inform_L[247][0] = l_cell_wire[247];							inform_L[248][0] = l_cell_wire[248];							inform_L[249][0] = l_cell_wire[249];							inform_L[250][0] = l_cell_wire[250];							inform_L[251][0] = l_cell_wire[251];							inform_L[252][0] = l_cell_wire[252];							inform_L[253][0] = l_cell_wire[253];							inform_L[254][0] = l_cell_wire[254];							inform_L[255][0] = l_cell_wire[255];							inform_L[256][0] = l_cell_wire[256];							inform_L[257][0] = l_cell_wire[257];							inform_L[258][0] = l_cell_wire[258];							inform_L[259][0] = l_cell_wire[259];							inform_L[260][0] = l_cell_wire[260];							inform_L[261][0] = l_cell_wire[261];							inform_L[262][0] = l_cell_wire[262];							inform_L[263][0] = l_cell_wire[263];							inform_L[264][0] = l_cell_wire[264];							inform_L[265][0] = l_cell_wire[265];							inform_L[266][0] = l_cell_wire[266];							inform_L[267][0] = l_cell_wire[267];							inform_L[268][0] = l_cell_wire[268];							inform_L[269][0] = l_cell_wire[269];							inform_L[270][0] = l_cell_wire[270];							inform_L[271][0] = l_cell_wire[271];							inform_L[272][0] = l_cell_wire[272];							inform_L[273][0] = l_cell_wire[273];							inform_L[274][0] = l_cell_wire[274];							inform_L[275][0] = l_cell_wire[275];							inform_L[276][0] = l_cell_wire[276];							inform_L[277][0] = l_cell_wire[277];							inform_L[278][0] = l_cell_wire[278];							inform_L[279][0] = l_cell_wire[279];							inform_L[280][0] = l_cell_wire[280];							inform_L[281][0] = l_cell_wire[281];							inform_L[282][0] = l_cell_wire[282];							inform_L[283][0] = l_cell_wire[283];							inform_L[284][0] = l_cell_wire[284];							inform_L[285][0] = l_cell_wire[285];							inform_L[286][0] = l_cell_wire[286];							inform_L[287][0] = l_cell_wire[287];							inform_L[288][0] = l_cell_wire[288];							inform_L[289][0] = l_cell_wire[289];							inform_L[290][0] = l_cell_wire[290];							inform_L[291][0] = l_cell_wire[291];							inform_L[292][0] = l_cell_wire[292];							inform_L[293][0] = l_cell_wire[293];							inform_L[294][0] = l_cell_wire[294];							inform_L[295][0] = l_cell_wire[295];							inform_L[296][0] = l_cell_wire[296];							inform_L[297][0] = l_cell_wire[297];							inform_L[298][0] = l_cell_wire[298];							inform_L[299][0] = l_cell_wire[299];							inform_L[300][0] = l_cell_wire[300];							inform_L[301][0] = l_cell_wire[301];							inform_L[302][0] = l_cell_wire[302];							inform_L[303][0] = l_cell_wire[303];							inform_L[304][0] = l_cell_wire[304];							inform_L[305][0] = l_cell_wire[305];							inform_L[306][0] = l_cell_wire[306];							inform_L[307][0] = l_cell_wire[307];							inform_L[308][0] = l_cell_wire[308];							inform_L[309][0] = l_cell_wire[309];							inform_L[310][0] = l_cell_wire[310];							inform_L[311][0] = l_cell_wire[311];							inform_L[312][0] = l_cell_wire[312];							inform_L[313][0] = l_cell_wire[313];							inform_L[314][0] = l_cell_wire[314];							inform_L[315][0] = l_cell_wire[315];							inform_L[316][0] = l_cell_wire[316];							inform_L[317][0] = l_cell_wire[317];							inform_L[318][0] = l_cell_wire[318];							inform_L[319][0] = l_cell_wire[319];							inform_L[320][0] = l_cell_wire[320];							inform_L[321][0] = l_cell_wire[321];							inform_L[322][0] = l_cell_wire[322];							inform_L[323][0] = l_cell_wire[323];							inform_L[324][0] = l_cell_wire[324];							inform_L[325][0] = l_cell_wire[325];							inform_L[326][0] = l_cell_wire[326];							inform_L[327][0] = l_cell_wire[327];							inform_L[328][0] = l_cell_wire[328];							inform_L[329][0] = l_cell_wire[329];							inform_L[330][0] = l_cell_wire[330];							inform_L[331][0] = l_cell_wire[331];							inform_L[332][0] = l_cell_wire[332];							inform_L[333][0] = l_cell_wire[333];							inform_L[334][0] = l_cell_wire[334];							inform_L[335][0] = l_cell_wire[335];							inform_L[336][0] = l_cell_wire[336];							inform_L[337][0] = l_cell_wire[337];							inform_L[338][0] = l_cell_wire[338];							inform_L[339][0] = l_cell_wire[339];							inform_L[340][0] = l_cell_wire[340];							inform_L[341][0] = l_cell_wire[341];							inform_L[342][0] = l_cell_wire[342];							inform_L[343][0] = l_cell_wire[343];							inform_L[344][0] = l_cell_wire[344];							inform_L[345][0] = l_cell_wire[345];							inform_L[346][0] = l_cell_wire[346];							inform_L[347][0] = l_cell_wire[347];							inform_L[348][0] = l_cell_wire[348];							inform_L[349][0] = l_cell_wire[349];							inform_L[350][0] = l_cell_wire[350];							inform_L[351][0] = l_cell_wire[351];							inform_L[352][0] = l_cell_wire[352];							inform_L[353][0] = l_cell_wire[353];							inform_L[354][0] = l_cell_wire[354];							inform_L[355][0] = l_cell_wire[355];							inform_L[356][0] = l_cell_wire[356];							inform_L[357][0] = l_cell_wire[357];							inform_L[358][0] = l_cell_wire[358];							inform_L[359][0] = l_cell_wire[359];							inform_L[360][0] = l_cell_wire[360];							inform_L[361][0] = l_cell_wire[361];							inform_L[362][0] = l_cell_wire[362];							inform_L[363][0] = l_cell_wire[363];							inform_L[364][0] = l_cell_wire[364];							inform_L[365][0] = l_cell_wire[365];							inform_L[366][0] = l_cell_wire[366];							inform_L[367][0] = l_cell_wire[367];							inform_L[368][0] = l_cell_wire[368];							inform_L[369][0] = l_cell_wire[369];							inform_L[370][0] = l_cell_wire[370];							inform_L[371][0] = l_cell_wire[371];							inform_L[372][0] = l_cell_wire[372];							inform_L[373][0] = l_cell_wire[373];							inform_L[374][0] = l_cell_wire[374];							inform_L[375][0] = l_cell_wire[375];							inform_L[376][0] = l_cell_wire[376];							inform_L[377][0] = l_cell_wire[377];							inform_L[378][0] = l_cell_wire[378];							inform_L[379][0] = l_cell_wire[379];							inform_L[380][0] = l_cell_wire[380];							inform_L[381][0] = l_cell_wire[381];							inform_L[382][0] = l_cell_wire[382];							inform_L[383][0] = l_cell_wire[383];							inform_L[384][0] = l_cell_wire[384];							inform_L[385][0] = l_cell_wire[385];							inform_L[386][0] = l_cell_wire[386];							inform_L[387][0] = l_cell_wire[387];							inform_L[388][0] = l_cell_wire[388];							inform_L[389][0] = l_cell_wire[389];							inform_L[390][0] = l_cell_wire[390];							inform_L[391][0] = l_cell_wire[391];							inform_L[392][0] = l_cell_wire[392];							inform_L[393][0] = l_cell_wire[393];							inform_L[394][0] = l_cell_wire[394];							inform_L[395][0] = l_cell_wire[395];							inform_L[396][0] = l_cell_wire[396];							inform_L[397][0] = l_cell_wire[397];							inform_L[398][0] = l_cell_wire[398];							inform_L[399][0] = l_cell_wire[399];							inform_L[400][0] = l_cell_wire[400];							inform_L[401][0] = l_cell_wire[401];							inform_L[402][0] = l_cell_wire[402];							inform_L[403][0] = l_cell_wire[403];							inform_L[404][0] = l_cell_wire[404];							inform_L[405][0] = l_cell_wire[405];							inform_L[406][0] = l_cell_wire[406];							inform_L[407][0] = l_cell_wire[407];							inform_L[408][0] = l_cell_wire[408];							inform_L[409][0] = l_cell_wire[409];							inform_L[410][0] = l_cell_wire[410];							inform_L[411][0] = l_cell_wire[411];							inform_L[412][0] = l_cell_wire[412];							inform_L[413][0] = l_cell_wire[413];							inform_L[414][0] = l_cell_wire[414];							inform_L[415][0] = l_cell_wire[415];							inform_L[416][0] = l_cell_wire[416];							inform_L[417][0] = l_cell_wire[417];							inform_L[418][0] = l_cell_wire[418];							inform_L[419][0] = l_cell_wire[419];							inform_L[420][0] = l_cell_wire[420];							inform_L[421][0] = l_cell_wire[421];							inform_L[422][0] = l_cell_wire[422];							inform_L[423][0] = l_cell_wire[423];							inform_L[424][0] = l_cell_wire[424];							inform_L[425][0] = l_cell_wire[425];							inform_L[426][0] = l_cell_wire[426];							inform_L[427][0] = l_cell_wire[427];							inform_L[428][0] = l_cell_wire[428];							inform_L[429][0] = l_cell_wire[429];							inform_L[430][0] = l_cell_wire[430];							inform_L[431][0] = l_cell_wire[431];							inform_L[432][0] = l_cell_wire[432];							inform_L[433][0] = l_cell_wire[433];							inform_L[434][0] = l_cell_wire[434];							inform_L[435][0] = l_cell_wire[435];							inform_L[436][0] = l_cell_wire[436];							inform_L[437][0] = l_cell_wire[437];							inform_L[438][0] = l_cell_wire[438];							inform_L[439][0] = l_cell_wire[439];							inform_L[440][0] = l_cell_wire[440];							inform_L[441][0] = l_cell_wire[441];							inform_L[442][0] = l_cell_wire[442];							inform_L[443][0] = l_cell_wire[443];							inform_L[444][0] = l_cell_wire[444];							inform_L[445][0] = l_cell_wire[445];							inform_L[446][0] = l_cell_wire[446];							inform_L[447][0] = l_cell_wire[447];							inform_L[448][0] = l_cell_wire[448];							inform_L[449][0] = l_cell_wire[449];							inform_L[450][0] = l_cell_wire[450];							inform_L[451][0] = l_cell_wire[451];							inform_L[452][0] = l_cell_wire[452];							inform_L[453][0] = l_cell_wire[453];							inform_L[454][0] = l_cell_wire[454];							inform_L[455][0] = l_cell_wire[455];							inform_L[456][0] = l_cell_wire[456];							inform_L[457][0] = l_cell_wire[457];							inform_L[458][0] = l_cell_wire[458];							inform_L[459][0] = l_cell_wire[459];							inform_L[460][0] = l_cell_wire[460];							inform_L[461][0] = l_cell_wire[461];							inform_L[462][0] = l_cell_wire[462];							inform_L[463][0] = l_cell_wire[463];							inform_L[464][0] = l_cell_wire[464];							inform_L[465][0] = l_cell_wire[465];							inform_L[466][0] = l_cell_wire[466];							inform_L[467][0] = l_cell_wire[467];							inform_L[468][0] = l_cell_wire[468];							inform_L[469][0] = l_cell_wire[469];							inform_L[470][0] = l_cell_wire[470];							inform_L[471][0] = l_cell_wire[471];							inform_L[472][0] = l_cell_wire[472];							inform_L[473][0] = l_cell_wire[473];							inform_L[474][0] = l_cell_wire[474];							inform_L[475][0] = l_cell_wire[475];							inform_L[476][0] = l_cell_wire[476];							inform_L[477][0] = l_cell_wire[477];							inform_L[478][0] = l_cell_wire[478];							inform_L[479][0] = l_cell_wire[479];							inform_L[480][0] = l_cell_wire[480];							inform_L[481][0] = l_cell_wire[481];							inform_L[482][0] = l_cell_wire[482];							inform_L[483][0] = l_cell_wire[483];							inform_L[484][0] = l_cell_wire[484];							inform_L[485][0] = l_cell_wire[485];							inform_L[486][0] = l_cell_wire[486];							inform_L[487][0] = l_cell_wire[487];							inform_L[488][0] = l_cell_wire[488];							inform_L[489][0] = l_cell_wire[489];							inform_L[490][0] = l_cell_wire[490];							inform_L[491][0] = l_cell_wire[491];							inform_L[492][0] = l_cell_wire[492];							inform_L[493][0] = l_cell_wire[493];							inform_L[494][0] = l_cell_wire[494];							inform_L[495][0] = l_cell_wire[495];							inform_L[496][0] = l_cell_wire[496];							inform_L[497][0] = l_cell_wire[497];							inform_L[498][0] = l_cell_wire[498];							inform_L[499][0] = l_cell_wire[499];							inform_L[500][0] = l_cell_wire[500];							inform_L[501][0] = l_cell_wire[501];							inform_L[502][0] = l_cell_wire[502];							inform_L[503][0] = l_cell_wire[503];							inform_L[504][0] = l_cell_wire[504];							inform_L[505][0] = l_cell_wire[505];							inform_L[506][0] = l_cell_wire[506];							inform_L[507][0] = l_cell_wire[507];							inform_L[508][0] = l_cell_wire[508];							inform_L[509][0] = l_cell_wire[509];							inform_L[510][0] = l_cell_wire[510];							inform_L[511][0] = l_cell_wire[511];							inform_L[512][0] = l_cell_wire[512];							inform_L[513][0] = l_cell_wire[513];							inform_L[514][0] = l_cell_wire[514];							inform_L[515][0] = l_cell_wire[515];							inform_L[516][0] = l_cell_wire[516];							inform_L[517][0] = l_cell_wire[517];							inform_L[518][0] = l_cell_wire[518];							inform_L[519][0] = l_cell_wire[519];							inform_L[520][0] = l_cell_wire[520];							inform_L[521][0] = l_cell_wire[521];							inform_L[522][0] = l_cell_wire[522];							inform_L[523][0] = l_cell_wire[523];							inform_L[524][0] = l_cell_wire[524];							inform_L[525][0] = l_cell_wire[525];							inform_L[526][0] = l_cell_wire[526];							inform_L[527][0] = l_cell_wire[527];							inform_L[528][0] = l_cell_wire[528];							inform_L[529][0] = l_cell_wire[529];							inform_L[530][0] = l_cell_wire[530];							inform_L[531][0] = l_cell_wire[531];							inform_L[532][0] = l_cell_wire[532];							inform_L[533][0] = l_cell_wire[533];							inform_L[534][0] = l_cell_wire[534];							inform_L[535][0] = l_cell_wire[535];							inform_L[536][0] = l_cell_wire[536];							inform_L[537][0] = l_cell_wire[537];							inform_L[538][0] = l_cell_wire[538];							inform_L[539][0] = l_cell_wire[539];							inform_L[540][0] = l_cell_wire[540];							inform_L[541][0] = l_cell_wire[541];							inform_L[542][0] = l_cell_wire[542];							inform_L[543][0] = l_cell_wire[543];							inform_L[544][0] = l_cell_wire[544];							inform_L[545][0] = l_cell_wire[545];							inform_L[546][0] = l_cell_wire[546];							inform_L[547][0] = l_cell_wire[547];							inform_L[548][0] = l_cell_wire[548];							inform_L[549][0] = l_cell_wire[549];							inform_L[550][0] = l_cell_wire[550];							inform_L[551][0] = l_cell_wire[551];							inform_L[552][0] = l_cell_wire[552];							inform_L[553][0] = l_cell_wire[553];							inform_L[554][0] = l_cell_wire[554];							inform_L[555][0] = l_cell_wire[555];							inform_L[556][0] = l_cell_wire[556];							inform_L[557][0] = l_cell_wire[557];							inform_L[558][0] = l_cell_wire[558];							inform_L[559][0] = l_cell_wire[559];							inform_L[560][0] = l_cell_wire[560];							inform_L[561][0] = l_cell_wire[561];							inform_L[562][0] = l_cell_wire[562];							inform_L[563][0] = l_cell_wire[563];							inform_L[564][0] = l_cell_wire[564];							inform_L[565][0] = l_cell_wire[565];							inform_L[566][0] = l_cell_wire[566];							inform_L[567][0] = l_cell_wire[567];							inform_L[568][0] = l_cell_wire[568];							inform_L[569][0] = l_cell_wire[569];							inform_L[570][0] = l_cell_wire[570];							inform_L[571][0] = l_cell_wire[571];							inform_L[572][0] = l_cell_wire[572];							inform_L[573][0] = l_cell_wire[573];							inform_L[574][0] = l_cell_wire[574];							inform_L[575][0] = l_cell_wire[575];							inform_L[576][0] = l_cell_wire[576];							inform_L[577][0] = l_cell_wire[577];							inform_L[578][0] = l_cell_wire[578];							inform_L[579][0] = l_cell_wire[579];							inform_L[580][0] = l_cell_wire[580];							inform_L[581][0] = l_cell_wire[581];							inform_L[582][0] = l_cell_wire[582];							inform_L[583][0] = l_cell_wire[583];							inform_L[584][0] = l_cell_wire[584];							inform_L[585][0] = l_cell_wire[585];							inform_L[586][0] = l_cell_wire[586];							inform_L[587][0] = l_cell_wire[587];							inform_L[588][0] = l_cell_wire[588];							inform_L[589][0] = l_cell_wire[589];							inform_L[590][0] = l_cell_wire[590];							inform_L[591][0] = l_cell_wire[591];							inform_L[592][0] = l_cell_wire[592];							inform_L[593][0] = l_cell_wire[593];							inform_L[594][0] = l_cell_wire[594];							inform_L[595][0] = l_cell_wire[595];							inform_L[596][0] = l_cell_wire[596];							inform_L[597][0] = l_cell_wire[597];							inform_L[598][0] = l_cell_wire[598];							inform_L[599][0] = l_cell_wire[599];							inform_L[600][0] = l_cell_wire[600];							inform_L[601][0] = l_cell_wire[601];							inform_L[602][0] = l_cell_wire[602];							inform_L[603][0] = l_cell_wire[603];							inform_L[604][0] = l_cell_wire[604];							inform_L[605][0] = l_cell_wire[605];							inform_L[606][0] = l_cell_wire[606];							inform_L[607][0] = l_cell_wire[607];							inform_L[608][0] = l_cell_wire[608];							inform_L[609][0] = l_cell_wire[609];							inform_L[610][0] = l_cell_wire[610];							inform_L[611][0] = l_cell_wire[611];							inform_L[612][0] = l_cell_wire[612];							inform_L[613][0] = l_cell_wire[613];							inform_L[614][0] = l_cell_wire[614];							inform_L[615][0] = l_cell_wire[615];							inform_L[616][0] = l_cell_wire[616];							inform_L[617][0] = l_cell_wire[617];							inform_L[618][0] = l_cell_wire[618];							inform_L[619][0] = l_cell_wire[619];							inform_L[620][0] = l_cell_wire[620];							inform_L[621][0] = l_cell_wire[621];							inform_L[622][0] = l_cell_wire[622];							inform_L[623][0] = l_cell_wire[623];							inform_L[624][0] = l_cell_wire[624];							inform_L[625][0] = l_cell_wire[625];							inform_L[626][0] = l_cell_wire[626];							inform_L[627][0] = l_cell_wire[627];							inform_L[628][0] = l_cell_wire[628];							inform_L[629][0] = l_cell_wire[629];							inform_L[630][0] = l_cell_wire[630];							inform_L[631][0] = l_cell_wire[631];							inform_L[632][0] = l_cell_wire[632];							inform_L[633][0] = l_cell_wire[633];							inform_L[634][0] = l_cell_wire[634];							inform_L[635][0] = l_cell_wire[635];							inform_L[636][0] = l_cell_wire[636];							inform_L[637][0] = l_cell_wire[637];							inform_L[638][0] = l_cell_wire[638];							inform_L[639][0] = l_cell_wire[639];							inform_L[640][0] = l_cell_wire[640];							inform_L[641][0] = l_cell_wire[641];							inform_L[642][0] = l_cell_wire[642];							inform_L[643][0] = l_cell_wire[643];							inform_L[644][0] = l_cell_wire[644];							inform_L[645][0] = l_cell_wire[645];							inform_L[646][0] = l_cell_wire[646];							inform_L[647][0] = l_cell_wire[647];							inform_L[648][0] = l_cell_wire[648];							inform_L[649][0] = l_cell_wire[649];							inform_L[650][0] = l_cell_wire[650];							inform_L[651][0] = l_cell_wire[651];							inform_L[652][0] = l_cell_wire[652];							inform_L[653][0] = l_cell_wire[653];							inform_L[654][0] = l_cell_wire[654];							inform_L[655][0] = l_cell_wire[655];							inform_L[656][0] = l_cell_wire[656];							inform_L[657][0] = l_cell_wire[657];							inform_L[658][0] = l_cell_wire[658];							inform_L[659][0] = l_cell_wire[659];							inform_L[660][0] = l_cell_wire[660];							inform_L[661][0] = l_cell_wire[661];							inform_L[662][0] = l_cell_wire[662];							inform_L[663][0] = l_cell_wire[663];							inform_L[664][0] = l_cell_wire[664];							inform_L[665][0] = l_cell_wire[665];							inform_L[666][0] = l_cell_wire[666];							inform_L[667][0] = l_cell_wire[667];							inform_L[668][0] = l_cell_wire[668];							inform_L[669][0] = l_cell_wire[669];							inform_L[670][0] = l_cell_wire[670];							inform_L[671][0] = l_cell_wire[671];							inform_L[672][0] = l_cell_wire[672];							inform_L[673][0] = l_cell_wire[673];							inform_L[674][0] = l_cell_wire[674];							inform_L[675][0] = l_cell_wire[675];							inform_L[676][0] = l_cell_wire[676];							inform_L[677][0] = l_cell_wire[677];							inform_L[678][0] = l_cell_wire[678];							inform_L[679][0] = l_cell_wire[679];							inform_L[680][0] = l_cell_wire[680];							inform_L[681][0] = l_cell_wire[681];							inform_L[682][0] = l_cell_wire[682];							inform_L[683][0] = l_cell_wire[683];							inform_L[684][0] = l_cell_wire[684];							inform_L[685][0] = l_cell_wire[685];							inform_L[686][0] = l_cell_wire[686];							inform_L[687][0] = l_cell_wire[687];							inform_L[688][0] = l_cell_wire[688];							inform_L[689][0] = l_cell_wire[689];							inform_L[690][0] = l_cell_wire[690];							inform_L[691][0] = l_cell_wire[691];							inform_L[692][0] = l_cell_wire[692];							inform_L[693][0] = l_cell_wire[693];							inform_L[694][0] = l_cell_wire[694];							inform_L[695][0] = l_cell_wire[695];							inform_L[696][0] = l_cell_wire[696];							inform_L[697][0] = l_cell_wire[697];							inform_L[698][0] = l_cell_wire[698];							inform_L[699][0] = l_cell_wire[699];							inform_L[700][0] = l_cell_wire[700];							inform_L[701][0] = l_cell_wire[701];							inform_L[702][0] = l_cell_wire[702];							inform_L[703][0] = l_cell_wire[703];							inform_L[704][0] = l_cell_wire[704];							inform_L[705][0] = l_cell_wire[705];							inform_L[706][0] = l_cell_wire[706];							inform_L[707][0] = l_cell_wire[707];							inform_L[708][0] = l_cell_wire[708];							inform_L[709][0] = l_cell_wire[709];							inform_L[710][0] = l_cell_wire[710];							inform_L[711][0] = l_cell_wire[711];							inform_L[712][0] = l_cell_wire[712];							inform_L[713][0] = l_cell_wire[713];							inform_L[714][0] = l_cell_wire[714];							inform_L[715][0] = l_cell_wire[715];							inform_L[716][0] = l_cell_wire[716];							inform_L[717][0] = l_cell_wire[717];							inform_L[718][0] = l_cell_wire[718];							inform_L[719][0] = l_cell_wire[719];							inform_L[720][0] = l_cell_wire[720];							inform_L[721][0] = l_cell_wire[721];							inform_L[722][0] = l_cell_wire[722];							inform_L[723][0] = l_cell_wire[723];							inform_L[724][0] = l_cell_wire[724];							inform_L[725][0] = l_cell_wire[725];							inform_L[726][0] = l_cell_wire[726];							inform_L[727][0] = l_cell_wire[727];							inform_L[728][0] = l_cell_wire[728];							inform_L[729][0] = l_cell_wire[729];							inform_L[730][0] = l_cell_wire[730];							inform_L[731][0] = l_cell_wire[731];							inform_L[732][0] = l_cell_wire[732];							inform_L[733][0] = l_cell_wire[733];							inform_L[734][0] = l_cell_wire[734];							inform_L[735][0] = l_cell_wire[735];							inform_L[736][0] = l_cell_wire[736];							inform_L[737][0] = l_cell_wire[737];							inform_L[738][0] = l_cell_wire[738];							inform_L[739][0] = l_cell_wire[739];							inform_L[740][0] = l_cell_wire[740];							inform_L[741][0] = l_cell_wire[741];							inform_L[742][0] = l_cell_wire[742];							inform_L[743][0] = l_cell_wire[743];							inform_L[744][0] = l_cell_wire[744];							inform_L[745][0] = l_cell_wire[745];							inform_L[746][0] = l_cell_wire[746];							inform_L[747][0] = l_cell_wire[747];							inform_L[748][0] = l_cell_wire[748];							inform_L[749][0] = l_cell_wire[749];							inform_L[750][0] = l_cell_wire[750];							inform_L[751][0] = l_cell_wire[751];							inform_L[752][0] = l_cell_wire[752];							inform_L[753][0] = l_cell_wire[753];							inform_L[754][0] = l_cell_wire[754];							inform_L[755][0] = l_cell_wire[755];							inform_L[756][0] = l_cell_wire[756];							inform_L[757][0] = l_cell_wire[757];							inform_L[758][0] = l_cell_wire[758];							inform_L[759][0] = l_cell_wire[759];							inform_L[760][0] = l_cell_wire[760];							inform_L[761][0] = l_cell_wire[761];							inform_L[762][0] = l_cell_wire[762];							inform_L[763][0] = l_cell_wire[763];							inform_L[764][0] = l_cell_wire[764];							inform_L[765][0] = l_cell_wire[765];							inform_L[766][0] = l_cell_wire[766];							inform_L[767][0] = l_cell_wire[767];							inform_L[768][0] = l_cell_wire[768];							inform_L[769][0] = l_cell_wire[769];							inform_L[770][0] = l_cell_wire[770];							inform_L[771][0] = l_cell_wire[771];							inform_L[772][0] = l_cell_wire[772];							inform_L[773][0] = l_cell_wire[773];							inform_L[774][0] = l_cell_wire[774];							inform_L[775][0] = l_cell_wire[775];							inform_L[776][0] = l_cell_wire[776];							inform_L[777][0] = l_cell_wire[777];							inform_L[778][0] = l_cell_wire[778];							inform_L[779][0] = l_cell_wire[779];							inform_L[780][0] = l_cell_wire[780];							inform_L[781][0] = l_cell_wire[781];							inform_L[782][0] = l_cell_wire[782];							inform_L[783][0] = l_cell_wire[783];							inform_L[784][0] = l_cell_wire[784];							inform_L[785][0] = l_cell_wire[785];							inform_L[786][0] = l_cell_wire[786];							inform_L[787][0] = l_cell_wire[787];							inform_L[788][0] = l_cell_wire[788];							inform_L[789][0] = l_cell_wire[789];							inform_L[790][0] = l_cell_wire[790];							inform_L[791][0] = l_cell_wire[791];							inform_L[792][0] = l_cell_wire[792];							inform_L[793][0] = l_cell_wire[793];							inform_L[794][0] = l_cell_wire[794];							inform_L[795][0] = l_cell_wire[795];							inform_L[796][0] = l_cell_wire[796];							inform_L[797][0] = l_cell_wire[797];							inform_L[798][0] = l_cell_wire[798];							inform_L[799][0] = l_cell_wire[799];							inform_L[800][0] = l_cell_wire[800];							inform_L[801][0] = l_cell_wire[801];							inform_L[802][0] = l_cell_wire[802];							inform_L[803][0] = l_cell_wire[803];							inform_L[804][0] = l_cell_wire[804];							inform_L[805][0] = l_cell_wire[805];							inform_L[806][0] = l_cell_wire[806];							inform_L[807][0] = l_cell_wire[807];							inform_L[808][0] = l_cell_wire[808];							inform_L[809][0] = l_cell_wire[809];							inform_L[810][0] = l_cell_wire[810];							inform_L[811][0] = l_cell_wire[811];							inform_L[812][0] = l_cell_wire[812];							inform_L[813][0] = l_cell_wire[813];							inform_L[814][0] = l_cell_wire[814];							inform_L[815][0] = l_cell_wire[815];							inform_L[816][0] = l_cell_wire[816];							inform_L[817][0] = l_cell_wire[817];							inform_L[818][0] = l_cell_wire[818];							inform_L[819][0] = l_cell_wire[819];							inform_L[820][0] = l_cell_wire[820];							inform_L[821][0] = l_cell_wire[821];							inform_L[822][0] = l_cell_wire[822];							inform_L[823][0] = l_cell_wire[823];							inform_L[824][0] = l_cell_wire[824];							inform_L[825][0] = l_cell_wire[825];							inform_L[826][0] = l_cell_wire[826];							inform_L[827][0] = l_cell_wire[827];							inform_L[828][0] = l_cell_wire[828];							inform_L[829][0] = l_cell_wire[829];							inform_L[830][0] = l_cell_wire[830];							inform_L[831][0] = l_cell_wire[831];							inform_L[832][0] = l_cell_wire[832];							inform_L[833][0] = l_cell_wire[833];							inform_L[834][0] = l_cell_wire[834];							inform_L[835][0] = l_cell_wire[835];							inform_L[836][0] = l_cell_wire[836];							inform_L[837][0] = l_cell_wire[837];							inform_L[838][0] = l_cell_wire[838];							inform_L[839][0] = l_cell_wire[839];							inform_L[840][0] = l_cell_wire[840];							inform_L[841][0] = l_cell_wire[841];							inform_L[842][0] = l_cell_wire[842];							inform_L[843][0] = l_cell_wire[843];							inform_L[844][0] = l_cell_wire[844];							inform_L[845][0] = l_cell_wire[845];							inform_L[846][0] = l_cell_wire[846];							inform_L[847][0] = l_cell_wire[847];							inform_L[848][0] = l_cell_wire[848];							inform_L[849][0] = l_cell_wire[849];							inform_L[850][0] = l_cell_wire[850];							inform_L[851][0] = l_cell_wire[851];							inform_L[852][0] = l_cell_wire[852];							inform_L[853][0] = l_cell_wire[853];							inform_L[854][0] = l_cell_wire[854];							inform_L[855][0] = l_cell_wire[855];							inform_L[856][0] = l_cell_wire[856];							inform_L[857][0] = l_cell_wire[857];							inform_L[858][0] = l_cell_wire[858];							inform_L[859][0] = l_cell_wire[859];							inform_L[860][0] = l_cell_wire[860];							inform_L[861][0] = l_cell_wire[861];							inform_L[862][0] = l_cell_wire[862];							inform_L[863][0] = l_cell_wire[863];							inform_L[864][0] = l_cell_wire[864];							inform_L[865][0] = l_cell_wire[865];							inform_L[866][0] = l_cell_wire[866];							inform_L[867][0] = l_cell_wire[867];							inform_L[868][0] = l_cell_wire[868];							inform_L[869][0] = l_cell_wire[869];							inform_L[870][0] = l_cell_wire[870];							inform_L[871][0] = l_cell_wire[871];							inform_L[872][0] = l_cell_wire[872];							inform_L[873][0] = l_cell_wire[873];							inform_L[874][0] = l_cell_wire[874];							inform_L[875][0] = l_cell_wire[875];							inform_L[876][0] = l_cell_wire[876];							inform_L[877][0] = l_cell_wire[877];							inform_L[878][0] = l_cell_wire[878];							inform_L[879][0] = l_cell_wire[879];							inform_L[880][0] = l_cell_wire[880];							inform_L[881][0] = l_cell_wire[881];							inform_L[882][0] = l_cell_wire[882];							inform_L[883][0] = l_cell_wire[883];							inform_L[884][0] = l_cell_wire[884];							inform_L[885][0] = l_cell_wire[885];							inform_L[886][0] = l_cell_wire[886];							inform_L[887][0] = l_cell_wire[887];							inform_L[888][0] = l_cell_wire[888];							inform_L[889][0] = l_cell_wire[889];							inform_L[890][0] = l_cell_wire[890];							inform_L[891][0] = l_cell_wire[891];							inform_L[892][0] = l_cell_wire[892];							inform_L[893][0] = l_cell_wire[893];							inform_L[894][0] = l_cell_wire[894];							inform_L[895][0] = l_cell_wire[895];							inform_L[896][0] = l_cell_wire[896];							inform_L[897][0] = l_cell_wire[897];							inform_L[898][0] = l_cell_wire[898];							inform_L[899][0] = l_cell_wire[899];							inform_L[900][0] = l_cell_wire[900];							inform_L[901][0] = l_cell_wire[901];							inform_L[902][0] = l_cell_wire[902];							inform_L[903][0] = l_cell_wire[903];							inform_L[904][0] = l_cell_wire[904];							inform_L[905][0] = l_cell_wire[905];							inform_L[906][0] = l_cell_wire[906];							inform_L[907][0] = l_cell_wire[907];							inform_L[908][0] = l_cell_wire[908];							inform_L[909][0] = l_cell_wire[909];							inform_L[910][0] = l_cell_wire[910];							inform_L[911][0] = l_cell_wire[911];							inform_L[912][0] = l_cell_wire[912];							inform_L[913][0] = l_cell_wire[913];							inform_L[914][0] = l_cell_wire[914];							inform_L[915][0] = l_cell_wire[915];							inform_L[916][0] = l_cell_wire[916];							inform_L[917][0] = l_cell_wire[917];							inform_L[918][0] = l_cell_wire[918];							inform_L[919][0] = l_cell_wire[919];							inform_L[920][0] = l_cell_wire[920];							inform_L[921][0] = l_cell_wire[921];							inform_L[922][0] = l_cell_wire[922];							inform_L[923][0] = l_cell_wire[923];							inform_L[924][0] = l_cell_wire[924];							inform_L[925][0] = l_cell_wire[925];							inform_L[926][0] = l_cell_wire[926];							inform_L[927][0] = l_cell_wire[927];							inform_L[928][0] = l_cell_wire[928];							inform_L[929][0] = l_cell_wire[929];							inform_L[930][0] = l_cell_wire[930];							inform_L[931][0] = l_cell_wire[931];							inform_L[932][0] = l_cell_wire[932];							inform_L[933][0] = l_cell_wire[933];							inform_L[934][0] = l_cell_wire[934];							inform_L[935][0] = l_cell_wire[935];							inform_L[936][0] = l_cell_wire[936];							inform_L[937][0] = l_cell_wire[937];							inform_L[938][0] = l_cell_wire[938];							inform_L[939][0] = l_cell_wire[939];							inform_L[940][0] = l_cell_wire[940];							inform_L[941][0] = l_cell_wire[941];							inform_L[942][0] = l_cell_wire[942];							inform_L[943][0] = l_cell_wire[943];							inform_L[944][0] = l_cell_wire[944];							inform_L[945][0] = l_cell_wire[945];							inform_L[946][0] = l_cell_wire[946];							inform_L[947][0] = l_cell_wire[947];							inform_L[948][0] = l_cell_wire[948];							inform_L[949][0] = l_cell_wire[949];							inform_L[950][0] = l_cell_wire[950];							inform_L[951][0] = l_cell_wire[951];							inform_L[952][0] = l_cell_wire[952];							inform_L[953][0] = l_cell_wire[953];							inform_L[954][0] = l_cell_wire[954];							inform_L[955][0] = l_cell_wire[955];							inform_L[956][0] = l_cell_wire[956];							inform_L[957][0] = l_cell_wire[957];							inform_L[958][0] = l_cell_wire[958];							inform_L[959][0] = l_cell_wire[959];							inform_L[960][0] = l_cell_wire[960];							inform_L[961][0] = l_cell_wire[961];							inform_L[962][0] = l_cell_wire[962];							inform_L[963][0] = l_cell_wire[963];							inform_L[964][0] = l_cell_wire[964];							inform_L[965][0] = l_cell_wire[965];							inform_L[966][0] = l_cell_wire[966];							inform_L[967][0] = l_cell_wire[967];							inform_L[968][0] = l_cell_wire[968];							inform_L[969][0] = l_cell_wire[969];							inform_L[970][0] = l_cell_wire[970];							inform_L[971][0] = l_cell_wire[971];							inform_L[972][0] = l_cell_wire[972];							inform_L[973][0] = l_cell_wire[973];							inform_L[974][0] = l_cell_wire[974];							inform_L[975][0] = l_cell_wire[975];							inform_L[976][0] = l_cell_wire[976];							inform_L[977][0] = l_cell_wire[977];							inform_L[978][0] = l_cell_wire[978];							inform_L[979][0] = l_cell_wire[979];							inform_L[980][0] = l_cell_wire[980];							inform_L[981][0] = l_cell_wire[981];							inform_L[982][0] = l_cell_wire[982];							inform_L[983][0] = l_cell_wire[983];							inform_L[984][0] = l_cell_wire[984];							inform_L[985][0] = l_cell_wire[985];							inform_L[986][0] = l_cell_wire[986];							inform_L[987][0] = l_cell_wire[987];							inform_L[988][0] = l_cell_wire[988];							inform_L[989][0] = l_cell_wire[989];							inform_L[990][0] = l_cell_wire[990];							inform_L[991][0] = l_cell_wire[991];							inform_L[992][0] = l_cell_wire[992];							inform_L[993][0] = l_cell_wire[993];							inform_L[994][0] = l_cell_wire[994];							inform_L[995][0] = l_cell_wire[995];							inform_L[996][0] = l_cell_wire[996];							inform_L[997][0] = l_cell_wire[997];							inform_L[998][0] = l_cell_wire[998];							inform_L[999][0] = l_cell_wire[999];							inform_L[1000][0] = l_cell_wire[1000];							inform_L[1001][0] = l_cell_wire[1001];							inform_L[1002][0] = l_cell_wire[1002];							inform_L[1003][0] = l_cell_wire[1003];							inform_L[1004][0] = l_cell_wire[1004];							inform_L[1005][0] = l_cell_wire[1005];							inform_L[1006][0] = l_cell_wire[1006];							inform_L[1007][0] = l_cell_wire[1007];							inform_L[1008][0] = l_cell_wire[1008];							inform_L[1009][0] = l_cell_wire[1009];							inform_L[1010][0] = l_cell_wire[1010];							inform_L[1011][0] = l_cell_wire[1011];							inform_L[1012][0] = l_cell_wire[1012];							inform_L[1013][0] = l_cell_wire[1013];							inform_L[1014][0] = l_cell_wire[1014];							inform_L[1015][0] = l_cell_wire[1015];							inform_L[1016][0] = l_cell_wire[1016];							inform_L[1017][0] = l_cell_wire[1017];							inform_L[1018][0] = l_cell_wire[1018];							inform_L[1019][0] = l_cell_wire[1019];							inform_L[1020][0] = l_cell_wire[1020];							inform_L[1021][0] = l_cell_wire[1021];							inform_L[1022][0] = l_cell_wire[1022];							inform_L[1023][0] = l_cell_wire[1023];						end
						2:						begin							inform_R[0][2] = r_cell_wire[0];							inform_R[2][2] = r_cell_wire[1];							inform_R[1][2] = r_cell_wire[2];							inform_R[3][2] = r_cell_wire[3];							inform_R[4][2] = r_cell_wire[4];							inform_R[6][2] = r_cell_wire[5];							inform_R[5][2] = r_cell_wire[6];							inform_R[7][2] = r_cell_wire[7];							inform_R[8][2] = r_cell_wire[8];							inform_R[10][2] = r_cell_wire[9];							inform_R[9][2] = r_cell_wire[10];							inform_R[11][2] = r_cell_wire[11];							inform_R[12][2] = r_cell_wire[12];							inform_R[14][2] = r_cell_wire[13];							inform_R[13][2] = r_cell_wire[14];							inform_R[15][2] = r_cell_wire[15];							inform_R[16][2] = r_cell_wire[16];							inform_R[18][2] = r_cell_wire[17];							inform_R[17][2] = r_cell_wire[18];							inform_R[19][2] = r_cell_wire[19];							inform_R[20][2] = r_cell_wire[20];							inform_R[22][2] = r_cell_wire[21];							inform_R[21][2] = r_cell_wire[22];							inform_R[23][2] = r_cell_wire[23];							inform_R[24][2] = r_cell_wire[24];							inform_R[26][2] = r_cell_wire[25];							inform_R[25][2] = r_cell_wire[26];							inform_R[27][2] = r_cell_wire[27];							inform_R[28][2] = r_cell_wire[28];							inform_R[30][2] = r_cell_wire[29];							inform_R[29][2] = r_cell_wire[30];							inform_R[31][2] = r_cell_wire[31];							inform_R[32][2] = r_cell_wire[32];							inform_R[34][2] = r_cell_wire[33];							inform_R[33][2] = r_cell_wire[34];							inform_R[35][2] = r_cell_wire[35];							inform_R[36][2] = r_cell_wire[36];							inform_R[38][2] = r_cell_wire[37];							inform_R[37][2] = r_cell_wire[38];							inform_R[39][2] = r_cell_wire[39];							inform_R[40][2] = r_cell_wire[40];							inform_R[42][2] = r_cell_wire[41];							inform_R[41][2] = r_cell_wire[42];							inform_R[43][2] = r_cell_wire[43];							inform_R[44][2] = r_cell_wire[44];							inform_R[46][2] = r_cell_wire[45];							inform_R[45][2] = r_cell_wire[46];							inform_R[47][2] = r_cell_wire[47];							inform_R[48][2] = r_cell_wire[48];							inform_R[50][2] = r_cell_wire[49];							inform_R[49][2] = r_cell_wire[50];							inform_R[51][2] = r_cell_wire[51];							inform_R[52][2] = r_cell_wire[52];							inform_R[54][2] = r_cell_wire[53];							inform_R[53][2] = r_cell_wire[54];							inform_R[55][2] = r_cell_wire[55];							inform_R[56][2] = r_cell_wire[56];							inform_R[58][2] = r_cell_wire[57];							inform_R[57][2] = r_cell_wire[58];							inform_R[59][2] = r_cell_wire[59];							inform_R[60][2] = r_cell_wire[60];							inform_R[62][2] = r_cell_wire[61];							inform_R[61][2] = r_cell_wire[62];							inform_R[63][2] = r_cell_wire[63];							inform_R[64][2] = r_cell_wire[64];							inform_R[66][2] = r_cell_wire[65];							inform_R[65][2] = r_cell_wire[66];							inform_R[67][2] = r_cell_wire[67];							inform_R[68][2] = r_cell_wire[68];							inform_R[70][2] = r_cell_wire[69];							inform_R[69][2] = r_cell_wire[70];							inform_R[71][2] = r_cell_wire[71];							inform_R[72][2] = r_cell_wire[72];							inform_R[74][2] = r_cell_wire[73];							inform_R[73][2] = r_cell_wire[74];							inform_R[75][2] = r_cell_wire[75];							inform_R[76][2] = r_cell_wire[76];							inform_R[78][2] = r_cell_wire[77];							inform_R[77][2] = r_cell_wire[78];							inform_R[79][2] = r_cell_wire[79];							inform_R[80][2] = r_cell_wire[80];							inform_R[82][2] = r_cell_wire[81];							inform_R[81][2] = r_cell_wire[82];							inform_R[83][2] = r_cell_wire[83];							inform_R[84][2] = r_cell_wire[84];							inform_R[86][2] = r_cell_wire[85];							inform_R[85][2] = r_cell_wire[86];							inform_R[87][2] = r_cell_wire[87];							inform_R[88][2] = r_cell_wire[88];							inform_R[90][2] = r_cell_wire[89];							inform_R[89][2] = r_cell_wire[90];							inform_R[91][2] = r_cell_wire[91];							inform_R[92][2] = r_cell_wire[92];							inform_R[94][2] = r_cell_wire[93];							inform_R[93][2] = r_cell_wire[94];							inform_R[95][2] = r_cell_wire[95];							inform_R[96][2] = r_cell_wire[96];							inform_R[98][2] = r_cell_wire[97];							inform_R[97][2] = r_cell_wire[98];							inform_R[99][2] = r_cell_wire[99];							inform_R[100][2] = r_cell_wire[100];							inform_R[102][2] = r_cell_wire[101];							inform_R[101][2] = r_cell_wire[102];							inform_R[103][2] = r_cell_wire[103];							inform_R[104][2] = r_cell_wire[104];							inform_R[106][2] = r_cell_wire[105];							inform_R[105][2] = r_cell_wire[106];							inform_R[107][2] = r_cell_wire[107];							inform_R[108][2] = r_cell_wire[108];							inform_R[110][2] = r_cell_wire[109];							inform_R[109][2] = r_cell_wire[110];							inform_R[111][2] = r_cell_wire[111];							inform_R[112][2] = r_cell_wire[112];							inform_R[114][2] = r_cell_wire[113];							inform_R[113][2] = r_cell_wire[114];							inform_R[115][2] = r_cell_wire[115];							inform_R[116][2] = r_cell_wire[116];							inform_R[118][2] = r_cell_wire[117];							inform_R[117][2] = r_cell_wire[118];							inform_R[119][2] = r_cell_wire[119];							inform_R[120][2] = r_cell_wire[120];							inform_R[122][2] = r_cell_wire[121];							inform_R[121][2] = r_cell_wire[122];							inform_R[123][2] = r_cell_wire[123];							inform_R[124][2] = r_cell_wire[124];							inform_R[126][2] = r_cell_wire[125];							inform_R[125][2] = r_cell_wire[126];							inform_R[127][2] = r_cell_wire[127];							inform_R[128][2] = r_cell_wire[128];							inform_R[130][2] = r_cell_wire[129];							inform_R[129][2] = r_cell_wire[130];							inform_R[131][2] = r_cell_wire[131];							inform_R[132][2] = r_cell_wire[132];							inform_R[134][2] = r_cell_wire[133];							inform_R[133][2] = r_cell_wire[134];							inform_R[135][2] = r_cell_wire[135];							inform_R[136][2] = r_cell_wire[136];							inform_R[138][2] = r_cell_wire[137];							inform_R[137][2] = r_cell_wire[138];							inform_R[139][2] = r_cell_wire[139];							inform_R[140][2] = r_cell_wire[140];							inform_R[142][2] = r_cell_wire[141];							inform_R[141][2] = r_cell_wire[142];							inform_R[143][2] = r_cell_wire[143];							inform_R[144][2] = r_cell_wire[144];							inform_R[146][2] = r_cell_wire[145];							inform_R[145][2] = r_cell_wire[146];							inform_R[147][2] = r_cell_wire[147];							inform_R[148][2] = r_cell_wire[148];							inform_R[150][2] = r_cell_wire[149];							inform_R[149][2] = r_cell_wire[150];							inform_R[151][2] = r_cell_wire[151];							inform_R[152][2] = r_cell_wire[152];							inform_R[154][2] = r_cell_wire[153];							inform_R[153][2] = r_cell_wire[154];							inform_R[155][2] = r_cell_wire[155];							inform_R[156][2] = r_cell_wire[156];							inform_R[158][2] = r_cell_wire[157];							inform_R[157][2] = r_cell_wire[158];							inform_R[159][2] = r_cell_wire[159];							inform_R[160][2] = r_cell_wire[160];							inform_R[162][2] = r_cell_wire[161];							inform_R[161][2] = r_cell_wire[162];							inform_R[163][2] = r_cell_wire[163];							inform_R[164][2] = r_cell_wire[164];							inform_R[166][2] = r_cell_wire[165];							inform_R[165][2] = r_cell_wire[166];							inform_R[167][2] = r_cell_wire[167];							inform_R[168][2] = r_cell_wire[168];							inform_R[170][2] = r_cell_wire[169];							inform_R[169][2] = r_cell_wire[170];							inform_R[171][2] = r_cell_wire[171];							inform_R[172][2] = r_cell_wire[172];							inform_R[174][2] = r_cell_wire[173];							inform_R[173][2] = r_cell_wire[174];							inform_R[175][2] = r_cell_wire[175];							inform_R[176][2] = r_cell_wire[176];							inform_R[178][2] = r_cell_wire[177];							inform_R[177][2] = r_cell_wire[178];							inform_R[179][2] = r_cell_wire[179];							inform_R[180][2] = r_cell_wire[180];							inform_R[182][2] = r_cell_wire[181];							inform_R[181][2] = r_cell_wire[182];							inform_R[183][2] = r_cell_wire[183];							inform_R[184][2] = r_cell_wire[184];							inform_R[186][2] = r_cell_wire[185];							inform_R[185][2] = r_cell_wire[186];							inform_R[187][2] = r_cell_wire[187];							inform_R[188][2] = r_cell_wire[188];							inform_R[190][2] = r_cell_wire[189];							inform_R[189][2] = r_cell_wire[190];							inform_R[191][2] = r_cell_wire[191];							inform_R[192][2] = r_cell_wire[192];							inform_R[194][2] = r_cell_wire[193];							inform_R[193][2] = r_cell_wire[194];							inform_R[195][2] = r_cell_wire[195];							inform_R[196][2] = r_cell_wire[196];							inform_R[198][2] = r_cell_wire[197];							inform_R[197][2] = r_cell_wire[198];							inform_R[199][2] = r_cell_wire[199];							inform_R[200][2] = r_cell_wire[200];							inform_R[202][2] = r_cell_wire[201];							inform_R[201][2] = r_cell_wire[202];							inform_R[203][2] = r_cell_wire[203];							inform_R[204][2] = r_cell_wire[204];							inform_R[206][2] = r_cell_wire[205];							inform_R[205][2] = r_cell_wire[206];							inform_R[207][2] = r_cell_wire[207];							inform_R[208][2] = r_cell_wire[208];							inform_R[210][2] = r_cell_wire[209];							inform_R[209][2] = r_cell_wire[210];							inform_R[211][2] = r_cell_wire[211];							inform_R[212][2] = r_cell_wire[212];							inform_R[214][2] = r_cell_wire[213];							inform_R[213][2] = r_cell_wire[214];							inform_R[215][2] = r_cell_wire[215];							inform_R[216][2] = r_cell_wire[216];							inform_R[218][2] = r_cell_wire[217];							inform_R[217][2] = r_cell_wire[218];							inform_R[219][2] = r_cell_wire[219];							inform_R[220][2] = r_cell_wire[220];							inform_R[222][2] = r_cell_wire[221];							inform_R[221][2] = r_cell_wire[222];							inform_R[223][2] = r_cell_wire[223];							inform_R[224][2] = r_cell_wire[224];							inform_R[226][2] = r_cell_wire[225];							inform_R[225][2] = r_cell_wire[226];							inform_R[227][2] = r_cell_wire[227];							inform_R[228][2] = r_cell_wire[228];							inform_R[230][2] = r_cell_wire[229];							inform_R[229][2] = r_cell_wire[230];							inform_R[231][2] = r_cell_wire[231];							inform_R[232][2] = r_cell_wire[232];							inform_R[234][2] = r_cell_wire[233];							inform_R[233][2] = r_cell_wire[234];							inform_R[235][2] = r_cell_wire[235];							inform_R[236][2] = r_cell_wire[236];							inform_R[238][2] = r_cell_wire[237];							inform_R[237][2] = r_cell_wire[238];							inform_R[239][2] = r_cell_wire[239];							inform_R[240][2] = r_cell_wire[240];							inform_R[242][2] = r_cell_wire[241];							inform_R[241][2] = r_cell_wire[242];							inform_R[243][2] = r_cell_wire[243];							inform_R[244][2] = r_cell_wire[244];							inform_R[246][2] = r_cell_wire[245];							inform_R[245][2] = r_cell_wire[246];							inform_R[247][2] = r_cell_wire[247];							inform_R[248][2] = r_cell_wire[248];							inform_R[250][2] = r_cell_wire[249];							inform_R[249][2] = r_cell_wire[250];							inform_R[251][2] = r_cell_wire[251];							inform_R[252][2] = r_cell_wire[252];							inform_R[254][2] = r_cell_wire[253];							inform_R[253][2] = r_cell_wire[254];							inform_R[255][2] = r_cell_wire[255];							inform_R[256][2] = r_cell_wire[256];							inform_R[258][2] = r_cell_wire[257];							inform_R[257][2] = r_cell_wire[258];							inform_R[259][2] = r_cell_wire[259];							inform_R[260][2] = r_cell_wire[260];							inform_R[262][2] = r_cell_wire[261];							inform_R[261][2] = r_cell_wire[262];							inform_R[263][2] = r_cell_wire[263];							inform_R[264][2] = r_cell_wire[264];							inform_R[266][2] = r_cell_wire[265];							inform_R[265][2] = r_cell_wire[266];							inform_R[267][2] = r_cell_wire[267];							inform_R[268][2] = r_cell_wire[268];							inform_R[270][2] = r_cell_wire[269];							inform_R[269][2] = r_cell_wire[270];							inform_R[271][2] = r_cell_wire[271];							inform_R[272][2] = r_cell_wire[272];							inform_R[274][2] = r_cell_wire[273];							inform_R[273][2] = r_cell_wire[274];							inform_R[275][2] = r_cell_wire[275];							inform_R[276][2] = r_cell_wire[276];							inform_R[278][2] = r_cell_wire[277];							inform_R[277][2] = r_cell_wire[278];							inform_R[279][2] = r_cell_wire[279];							inform_R[280][2] = r_cell_wire[280];							inform_R[282][2] = r_cell_wire[281];							inform_R[281][2] = r_cell_wire[282];							inform_R[283][2] = r_cell_wire[283];							inform_R[284][2] = r_cell_wire[284];							inform_R[286][2] = r_cell_wire[285];							inform_R[285][2] = r_cell_wire[286];							inform_R[287][2] = r_cell_wire[287];							inform_R[288][2] = r_cell_wire[288];							inform_R[290][2] = r_cell_wire[289];							inform_R[289][2] = r_cell_wire[290];							inform_R[291][2] = r_cell_wire[291];							inform_R[292][2] = r_cell_wire[292];							inform_R[294][2] = r_cell_wire[293];							inform_R[293][2] = r_cell_wire[294];							inform_R[295][2] = r_cell_wire[295];							inform_R[296][2] = r_cell_wire[296];							inform_R[298][2] = r_cell_wire[297];							inform_R[297][2] = r_cell_wire[298];							inform_R[299][2] = r_cell_wire[299];							inform_R[300][2] = r_cell_wire[300];							inform_R[302][2] = r_cell_wire[301];							inform_R[301][2] = r_cell_wire[302];							inform_R[303][2] = r_cell_wire[303];							inform_R[304][2] = r_cell_wire[304];							inform_R[306][2] = r_cell_wire[305];							inform_R[305][2] = r_cell_wire[306];							inform_R[307][2] = r_cell_wire[307];							inform_R[308][2] = r_cell_wire[308];							inform_R[310][2] = r_cell_wire[309];							inform_R[309][2] = r_cell_wire[310];							inform_R[311][2] = r_cell_wire[311];							inform_R[312][2] = r_cell_wire[312];							inform_R[314][2] = r_cell_wire[313];							inform_R[313][2] = r_cell_wire[314];							inform_R[315][2] = r_cell_wire[315];							inform_R[316][2] = r_cell_wire[316];							inform_R[318][2] = r_cell_wire[317];							inform_R[317][2] = r_cell_wire[318];							inform_R[319][2] = r_cell_wire[319];							inform_R[320][2] = r_cell_wire[320];							inform_R[322][2] = r_cell_wire[321];							inform_R[321][2] = r_cell_wire[322];							inform_R[323][2] = r_cell_wire[323];							inform_R[324][2] = r_cell_wire[324];							inform_R[326][2] = r_cell_wire[325];							inform_R[325][2] = r_cell_wire[326];							inform_R[327][2] = r_cell_wire[327];							inform_R[328][2] = r_cell_wire[328];							inform_R[330][2] = r_cell_wire[329];							inform_R[329][2] = r_cell_wire[330];							inform_R[331][2] = r_cell_wire[331];							inform_R[332][2] = r_cell_wire[332];							inform_R[334][2] = r_cell_wire[333];							inform_R[333][2] = r_cell_wire[334];							inform_R[335][2] = r_cell_wire[335];							inform_R[336][2] = r_cell_wire[336];							inform_R[338][2] = r_cell_wire[337];							inform_R[337][2] = r_cell_wire[338];							inform_R[339][2] = r_cell_wire[339];							inform_R[340][2] = r_cell_wire[340];							inform_R[342][2] = r_cell_wire[341];							inform_R[341][2] = r_cell_wire[342];							inform_R[343][2] = r_cell_wire[343];							inform_R[344][2] = r_cell_wire[344];							inform_R[346][2] = r_cell_wire[345];							inform_R[345][2] = r_cell_wire[346];							inform_R[347][2] = r_cell_wire[347];							inform_R[348][2] = r_cell_wire[348];							inform_R[350][2] = r_cell_wire[349];							inform_R[349][2] = r_cell_wire[350];							inform_R[351][2] = r_cell_wire[351];							inform_R[352][2] = r_cell_wire[352];							inform_R[354][2] = r_cell_wire[353];							inform_R[353][2] = r_cell_wire[354];							inform_R[355][2] = r_cell_wire[355];							inform_R[356][2] = r_cell_wire[356];							inform_R[358][2] = r_cell_wire[357];							inform_R[357][2] = r_cell_wire[358];							inform_R[359][2] = r_cell_wire[359];							inform_R[360][2] = r_cell_wire[360];							inform_R[362][2] = r_cell_wire[361];							inform_R[361][2] = r_cell_wire[362];							inform_R[363][2] = r_cell_wire[363];							inform_R[364][2] = r_cell_wire[364];							inform_R[366][2] = r_cell_wire[365];							inform_R[365][2] = r_cell_wire[366];							inform_R[367][2] = r_cell_wire[367];							inform_R[368][2] = r_cell_wire[368];							inform_R[370][2] = r_cell_wire[369];							inform_R[369][2] = r_cell_wire[370];							inform_R[371][2] = r_cell_wire[371];							inform_R[372][2] = r_cell_wire[372];							inform_R[374][2] = r_cell_wire[373];							inform_R[373][2] = r_cell_wire[374];							inform_R[375][2] = r_cell_wire[375];							inform_R[376][2] = r_cell_wire[376];							inform_R[378][2] = r_cell_wire[377];							inform_R[377][2] = r_cell_wire[378];							inform_R[379][2] = r_cell_wire[379];							inform_R[380][2] = r_cell_wire[380];							inform_R[382][2] = r_cell_wire[381];							inform_R[381][2] = r_cell_wire[382];							inform_R[383][2] = r_cell_wire[383];							inform_R[384][2] = r_cell_wire[384];							inform_R[386][2] = r_cell_wire[385];							inform_R[385][2] = r_cell_wire[386];							inform_R[387][2] = r_cell_wire[387];							inform_R[388][2] = r_cell_wire[388];							inform_R[390][2] = r_cell_wire[389];							inform_R[389][2] = r_cell_wire[390];							inform_R[391][2] = r_cell_wire[391];							inform_R[392][2] = r_cell_wire[392];							inform_R[394][2] = r_cell_wire[393];							inform_R[393][2] = r_cell_wire[394];							inform_R[395][2] = r_cell_wire[395];							inform_R[396][2] = r_cell_wire[396];							inform_R[398][2] = r_cell_wire[397];							inform_R[397][2] = r_cell_wire[398];							inform_R[399][2] = r_cell_wire[399];							inform_R[400][2] = r_cell_wire[400];							inform_R[402][2] = r_cell_wire[401];							inform_R[401][2] = r_cell_wire[402];							inform_R[403][2] = r_cell_wire[403];							inform_R[404][2] = r_cell_wire[404];							inform_R[406][2] = r_cell_wire[405];							inform_R[405][2] = r_cell_wire[406];							inform_R[407][2] = r_cell_wire[407];							inform_R[408][2] = r_cell_wire[408];							inform_R[410][2] = r_cell_wire[409];							inform_R[409][2] = r_cell_wire[410];							inform_R[411][2] = r_cell_wire[411];							inform_R[412][2] = r_cell_wire[412];							inform_R[414][2] = r_cell_wire[413];							inform_R[413][2] = r_cell_wire[414];							inform_R[415][2] = r_cell_wire[415];							inform_R[416][2] = r_cell_wire[416];							inform_R[418][2] = r_cell_wire[417];							inform_R[417][2] = r_cell_wire[418];							inform_R[419][2] = r_cell_wire[419];							inform_R[420][2] = r_cell_wire[420];							inform_R[422][2] = r_cell_wire[421];							inform_R[421][2] = r_cell_wire[422];							inform_R[423][2] = r_cell_wire[423];							inform_R[424][2] = r_cell_wire[424];							inform_R[426][2] = r_cell_wire[425];							inform_R[425][2] = r_cell_wire[426];							inform_R[427][2] = r_cell_wire[427];							inform_R[428][2] = r_cell_wire[428];							inform_R[430][2] = r_cell_wire[429];							inform_R[429][2] = r_cell_wire[430];							inform_R[431][2] = r_cell_wire[431];							inform_R[432][2] = r_cell_wire[432];							inform_R[434][2] = r_cell_wire[433];							inform_R[433][2] = r_cell_wire[434];							inform_R[435][2] = r_cell_wire[435];							inform_R[436][2] = r_cell_wire[436];							inform_R[438][2] = r_cell_wire[437];							inform_R[437][2] = r_cell_wire[438];							inform_R[439][2] = r_cell_wire[439];							inform_R[440][2] = r_cell_wire[440];							inform_R[442][2] = r_cell_wire[441];							inform_R[441][2] = r_cell_wire[442];							inform_R[443][2] = r_cell_wire[443];							inform_R[444][2] = r_cell_wire[444];							inform_R[446][2] = r_cell_wire[445];							inform_R[445][2] = r_cell_wire[446];							inform_R[447][2] = r_cell_wire[447];							inform_R[448][2] = r_cell_wire[448];							inform_R[450][2] = r_cell_wire[449];							inform_R[449][2] = r_cell_wire[450];							inform_R[451][2] = r_cell_wire[451];							inform_R[452][2] = r_cell_wire[452];							inform_R[454][2] = r_cell_wire[453];							inform_R[453][2] = r_cell_wire[454];							inform_R[455][2] = r_cell_wire[455];							inform_R[456][2] = r_cell_wire[456];							inform_R[458][2] = r_cell_wire[457];							inform_R[457][2] = r_cell_wire[458];							inform_R[459][2] = r_cell_wire[459];							inform_R[460][2] = r_cell_wire[460];							inform_R[462][2] = r_cell_wire[461];							inform_R[461][2] = r_cell_wire[462];							inform_R[463][2] = r_cell_wire[463];							inform_R[464][2] = r_cell_wire[464];							inform_R[466][2] = r_cell_wire[465];							inform_R[465][2] = r_cell_wire[466];							inform_R[467][2] = r_cell_wire[467];							inform_R[468][2] = r_cell_wire[468];							inform_R[470][2] = r_cell_wire[469];							inform_R[469][2] = r_cell_wire[470];							inform_R[471][2] = r_cell_wire[471];							inform_R[472][2] = r_cell_wire[472];							inform_R[474][2] = r_cell_wire[473];							inform_R[473][2] = r_cell_wire[474];							inform_R[475][2] = r_cell_wire[475];							inform_R[476][2] = r_cell_wire[476];							inform_R[478][2] = r_cell_wire[477];							inform_R[477][2] = r_cell_wire[478];							inform_R[479][2] = r_cell_wire[479];							inform_R[480][2] = r_cell_wire[480];							inform_R[482][2] = r_cell_wire[481];							inform_R[481][2] = r_cell_wire[482];							inform_R[483][2] = r_cell_wire[483];							inform_R[484][2] = r_cell_wire[484];							inform_R[486][2] = r_cell_wire[485];							inform_R[485][2] = r_cell_wire[486];							inform_R[487][2] = r_cell_wire[487];							inform_R[488][2] = r_cell_wire[488];							inform_R[490][2] = r_cell_wire[489];							inform_R[489][2] = r_cell_wire[490];							inform_R[491][2] = r_cell_wire[491];							inform_R[492][2] = r_cell_wire[492];							inform_R[494][2] = r_cell_wire[493];							inform_R[493][2] = r_cell_wire[494];							inform_R[495][2] = r_cell_wire[495];							inform_R[496][2] = r_cell_wire[496];							inform_R[498][2] = r_cell_wire[497];							inform_R[497][2] = r_cell_wire[498];							inform_R[499][2] = r_cell_wire[499];							inform_R[500][2] = r_cell_wire[500];							inform_R[502][2] = r_cell_wire[501];							inform_R[501][2] = r_cell_wire[502];							inform_R[503][2] = r_cell_wire[503];							inform_R[504][2] = r_cell_wire[504];							inform_R[506][2] = r_cell_wire[505];							inform_R[505][2] = r_cell_wire[506];							inform_R[507][2] = r_cell_wire[507];							inform_R[508][2] = r_cell_wire[508];							inform_R[510][2] = r_cell_wire[509];							inform_R[509][2] = r_cell_wire[510];							inform_R[511][2] = r_cell_wire[511];							inform_R[512][2] = r_cell_wire[512];							inform_R[514][2] = r_cell_wire[513];							inform_R[513][2] = r_cell_wire[514];							inform_R[515][2] = r_cell_wire[515];							inform_R[516][2] = r_cell_wire[516];							inform_R[518][2] = r_cell_wire[517];							inform_R[517][2] = r_cell_wire[518];							inform_R[519][2] = r_cell_wire[519];							inform_R[520][2] = r_cell_wire[520];							inform_R[522][2] = r_cell_wire[521];							inform_R[521][2] = r_cell_wire[522];							inform_R[523][2] = r_cell_wire[523];							inform_R[524][2] = r_cell_wire[524];							inform_R[526][2] = r_cell_wire[525];							inform_R[525][2] = r_cell_wire[526];							inform_R[527][2] = r_cell_wire[527];							inform_R[528][2] = r_cell_wire[528];							inform_R[530][2] = r_cell_wire[529];							inform_R[529][2] = r_cell_wire[530];							inform_R[531][2] = r_cell_wire[531];							inform_R[532][2] = r_cell_wire[532];							inform_R[534][2] = r_cell_wire[533];							inform_R[533][2] = r_cell_wire[534];							inform_R[535][2] = r_cell_wire[535];							inform_R[536][2] = r_cell_wire[536];							inform_R[538][2] = r_cell_wire[537];							inform_R[537][2] = r_cell_wire[538];							inform_R[539][2] = r_cell_wire[539];							inform_R[540][2] = r_cell_wire[540];							inform_R[542][2] = r_cell_wire[541];							inform_R[541][2] = r_cell_wire[542];							inform_R[543][2] = r_cell_wire[543];							inform_R[544][2] = r_cell_wire[544];							inform_R[546][2] = r_cell_wire[545];							inform_R[545][2] = r_cell_wire[546];							inform_R[547][2] = r_cell_wire[547];							inform_R[548][2] = r_cell_wire[548];							inform_R[550][2] = r_cell_wire[549];							inform_R[549][2] = r_cell_wire[550];							inform_R[551][2] = r_cell_wire[551];							inform_R[552][2] = r_cell_wire[552];							inform_R[554][2] = r_cell_wire[553];							inform_R[553][2] = r_cell_wire[554];							inform_R[555][2] = r_cell_wire[555];							inform_R[556][2] = r_cell_wire[556];							inform_R[558][2] = r_cell_wire[557];							inform_R[557][2] = r_cell_wire[558];							inform_R[559][2] = r_cell_wire[559];							inform_R[560][2] = r_cell_wire[560];							inform_R[562][2] = r_cell_wire[561];							inform_R[561][2] = r_cell_wire[562];							inform_R[563][2] = r_cell_wire[563];							inform_R[564][2] = r_cell_wire[564];							inform_R[566][2] = r_cell_wire[565];							inform_R[565][2] = r_cell_wire[566];							inform_R[567][2] = r_cell_wire[567];							inform_R[568][2] = r_cell_wire[568];							inform_R[570][2] = r_cell_wire[569];							inform_R[569][2] = r_cell_wire[570];							inform_R[571][2] = r_cell_wire[571];							inform_R[572][2] = r_cell_wire[572];							inform_R[574][2] = r_cell_wire[573];							inform_R[573][2] = r_cell_wire[574];							inform_R[575][2] = r_cell_wire[575];							inform_R[576][2] = r_cell_wire[576];							inform_R[578][2] = r_cell_wire[577];							inform_R[577][2] = r_cell_wire[578];							inform_R[579][2] = r_cell_wire[579];							inform_R[580][2] = r_cell_wire[580];							inform_R[582][2] = r_cell_wire[581];							inform_R[581][2] = r_cell_wire[582];							inform_R[583][2] = r_cell_wire[583];							inform_R[584][2] = r_cell_wire[584];							inform_R[586][2] = r_cell_wire[585];							inform_R[585][2] = r_cell_wire[586];							inform_R[587][2] = r_cell_wire[587];							inform_R[588][2] = r_cell_wire[588];							inform_R[590][2] = r_cell_wire[589];							inform_R[589][2] = r_cell_wire[590];							inform_R[591][2] = r_cell_wire[591];							inform_R[592][2] = r_cell_wire[592];							inform_R[594][2] = r_cell_wire[593];							inform_R[593][2] = r_cell_wire[594];							inform_R[595][2] = r_cell_wire[595];							inform_R[596][2] = r_cell_wire[596];							inform_R[598][2] = r_cell_wire[597];							inform_R[597][2] = r_cell_wire[598];							inform_R[599][2] = r_cell_wire[599];							inform_R[600][2] = r_cell_wire[600];							inform_R[602][2] = r_cell_wire[601];							inform_R[601][2] = r_cell_wire[602];							inform_R[603][2] = r_cell_wire[603];							inform_R[604][2] = r_cell_wire[604];							inform_R[606][2] = r_cell_wire[605];							inform_R[605][2] = r_cell_wire[606];							inform_R[607][2] = r_cell_wire[607];							inform_R[608][2] = r_cell_wire[608];							inform_R[610][2] = r_cell_wire[609];							inform_R[609][2] = r_cell_wire[610];							inform_R[611][2] = r_cell_wire[611];							inform_R[612][2] = r_cell_wire[612];							inform_R[614][2] = r_cell_wire[613];							inform_R[613][2] = r_cell_wire[614];							inform_R[615][2] = r_cell_wire[615];							inform_R[616][2] = r_cell_wire[616];							inform_R[618][2] = r_cell_wire[617];							inform_R[617][2] = r_cell_wire[618];							inform_R[619][2] = r_cell_wire[619];							inform_R[620][2] = r_cell_wire[620];							inform_R[622][2] = r_cell_wire[621];							inform_R[621][2] = r_cell_wire[622];							inform_R[623][2] = r_cell_wire[623];							inform_R[624][2] = r_cell_wire[624];							inform_R[626][2] = r_cell_wire[625];							inform_R[625][2] = r_cell_wire[626];							inform_R[627][2] = r_cell_wire[627];							inform_R[628][2] = r_cell_wire[628];							inform_R[630][2] = r_cell_wire[629];							inform_R[629][2] = r_cell_wire[630];							inform_R[631][2] = r_cell_wire[631];							inform_R[632][2] = r_cell_wire[632];							inform_R[634][2] = r_cell_wire[633];							inform_R[633][2] = r_cell_wire[634];							inform_R[635][2] = r_cell_wire[635];							inform_R[636][2] = r_cell_wire[636];							inform_R[638][2] = r_cell_wire[637];							inform_R[637][2] = r_cell_wire[638];							inform_R[639][2] = r_cell_wire[639];							inform_R[640][2] = r_cell_wire[640];							inform_R[642][2] = r_cell_wire[641];							inform_R[641][2] = r_cell_wire[642];							inform_R[643][2] = r_cell_wire[643];							inform_R[644][2] = r_cell_wire[644];							inform_R[646][2] = r_cell_wire[645];							inform_R[645][2] = r_cell_wire[646];							inform_R[647][2] = r_cell_wire[647];							inform_R[648][2] = r_cell_wire[648];							inform_R[650][2] = r_cell_wire[649];							inform_R[649][2] = r_cell_wire[650];							inform_R[651][2] = r_cell_wire[651];							inform_R[652][2] = r_cell_wire[652];							inform_R[654][2] = r_cell_wire[653];							inform_R[653][2] = r_cell_wire[654];							inform_R[655][2] = r_cell_wire[655];							inform_R[656][2] = r_cell_wire[656];							inform_R[658][2] = r_cell_wire[657];							inform_R[657][2] = r_cell_wire[658];							inform_R[659][2] = r_cell_wire[659];							inform_R[660][2] = r_cell_wire[660];							inform_R[662][2] = r_cell_wire[661];							inform_R[661][2] = r_cell_wire[662];							inform_R[663][2] = r_cell_wire[663];							inform_R[664][2] = r_cell_wire[664];							inform_R[666][2] = r_cell_wire[665];							inform_R[665][2] = r_cell_wire[666];							inform_R[667][2] = r_cell_wire[667];							inform_R[668][2] = r_cell_wire[668];							inform_R[670][2] = r_cell_wire[669];							inform_R[669][2] = r_cell_wire[670];							inform_R[671][2] = r_cell_wire[671];							inform_R[672][2] = r_cell_wire[672];							inform_R[674][2] = r_cell_wire[673];							inform_R[673][2] = r_cell_wire[674];							inform_R[675][2] = r_cell_wire[675];							inform_R[676][2] = r_cell_wire[676];							inform_R[678][2] = r_cell_wire[677];							inform_R[677][2] = r_cell_wire[678];							inform_R[679][2] = r_cell_wire[679];							inform_R[680][2] = r_cell_wire[680];							inform_R[682][2] = r_cell_wire[681];							inform_R[681][2] = r_cell_wire[682];							inform_R[683][2] = r_cell_wire[683];							inform_R[684][2] = r_cell_wire[684];							inform_R[686][2] = r_cell_wire[685];							inform_R[685][2] = r_cell_wire[686];							inform_R[687][2] = r_cell_wire[687];							inform_R[688][2] = r_cell_wire[688];							inform_R[690][2] = r_cell_wire[689];							inform_R[689][2] = r_cell_wire[690];							inform_R[691][2] = r_cell_wire[691];							inform_R[692][2] = r_cell_wire[692];							inform_R[694][2] = r_cell_wire[693];							inform_R[693][2] = r_cell_wire[694];							inform_R[695][2] = r_cell_wire[695];							inform_R[696][2] = r_cell_wire[696];							inform_R[698][2] = r_cell_wire[697];							inform_R[697][2] = r_cell_wire[698];							inform_R[699][2] = r_cell_wire[699];							inform_R[700][2] = r_cell_wire[700];							inform_R[702][2] = r_cell_wire[701];							inform_R[701][2] = r_cell_wire[702];							inform_R[703][2] = r_cell_wire[703];							inform_R[704][2] = r_cell_wire[704];							inform_R[706][2] = r_cell_wire[705];							inform_R[705][2] = r_cell_wire[706];							inform_R[707][2] = r_cell_wire[707];							inform_R[708][2] = r_cell_wire[708];							inform_R[710][2] = r_cell_wire[709];							inform_R[709][2] = r_cell_wire[710];							inform_R[711][2] = r_cell_wire[711];							inform_R[712][2] = r_cell_wire[712];							inform_R[714][2] = r_cell_wire[713];							inform_R[713][2] = r_cell_wire[714];							inform_R[715][2] = r_cell_wire[715];							inform_R[716][2] = r_cell_wire[716];							inform_R[718][2] = r_cell_wire[717];							inform_R[717][2] = r_cell_wire[718];							inform_R[719][2] = r_cell_wire[719];							inform_R[720][2] = r_cell_wire[720];							inform_R[722][2] = r_cell_wire[721];							inform_R[721][2] = r_cell_wire[722];							inform_R[723][2] = r_cell_wire[723];							inform_R[724][2] = r_cell_wire[724];							inform_R[726][2] = r_cell_wire[725];							inform_R[725][2] = r_cell_wire[726];							inform_R[727][2] = r_cell_wire[727];							inform_R[728][2] = r_cell_wire[728];							inform_R[730][2] = r_cell_wire[729];							inform_R[729][2] = r_cell_wire[730];							inform_R[731][2] = r_cell_wire[731];							inform_R[732][2] = r_cell_wire[732];							inform_R[734][2] = r_cell_wire[733];							inform_R[733][2] = r_cell_wire[734];							inform_R[735][2] = r_cell_wire[735];							inform_R[736][2] = r_cell_wire[736];							inform_R[738][2] = r_cell_wire[737];							inform_R[737][2] = r_cell_wire[738];							inform_R[739][2] = r_cell_wire[739];							inform_R[740][2] = r_cell_wire[740];							inform_R[742][2] = r_cell_wire[741];							inform_R[741][2] = r_cell_wire[742];							inform_R[743][2] = r_cell_wire[743];							inform_R[744][2] = r_cell_wire[744];							inform_R[746][2] = r_cell_wire[745];							inform_R[745][2] = r_cell_wire[746];							inform_R[747][2] = r_cell_wire[747];							inform_R[748][2] = r_cell_wire[748];							inform_R[750][2] = r_cell_wire[749];							inform_R[749][2] = r_cell_wire[750];							inform_R[751][2] = r_cell_wire[751];							inform_R[752][2] = r_cell_wire[752];							inform_R[754][2] = r_cell_wire[753];							inform_R[753][2] = r_cell_wire[754];							inform_R[755][2] = r_cell_wire[755];							inform_R[756][2] = r_cell_wire[756];							inform_R[758][2] = r_cell_wire[757];							inform_R[757][2] = r_cell_wire[758];							inform_R[759][2] = r_cell_wire[759];							inform_R[760][2] = r_cell_wire[760];							inform_R[762][2] = r_cell_wire[761];							inform_R[761][2] = r_cell_wire[762];							inform_R[763][2] = r_cell_wire[763];							inform_R[764][2] = r_cell_wire[764];							inform_R[766][2] = r_cell_wire[765];							inform_R[765][2] = r_cell_wire[766];							inform_R[767][2] = r_cell_wire[767];							inform_R[768][2] = r_cell_wire[768];							inform_R[770][2] = r_cell_wire[769];							inform_R[769][2] = r_cell_wire[770];							inform_R[771][2] = r_cell_wire[771];							inform_R[772][2] = r_cell_wire[772];							inform_R[774][2] = r_cell_wire[773];							inform_R[773][2] = r_cell_wire[774];							inform_R[775][2] = r_cell_wire[775];							inform_R[776][2] = r_cell_wire[776];							inform_R[778][2] = r_cell_wire[777];							inform_R[777][2] = r_cell_wire[778];							inform_R[779][2] = r_cell_wire[779];							inform_R[780][2] = r_cell_wire[780];							inform_R[782][2] = r_cell_wire[781];							inform_R[781][2] = r_cell_wire[782];							inform_R[783][2] = r_cell_wire[783];							inform_R[784][2] = r_cell_wire[784];							inform_R[786][2] = r_cell_wire[785];							inform_R[785][2] = r_cell_wire[786];							inform_R[787][2] = r_cell_wire[787];							inform_R[788][2] = r_cell_wire[788];							inform_R[790][2] = r_cell_wire[789];							inform_R[789][2] = r_cell_wire[790];							inform_R[791][2] = r_cell_wire[791];							inform_R[792][2] = r_cell_wire[792];							inform_R[794][2] = r_cell_wire[793];							inform_R[793][2] = r_cell_wire[794];							inform_R[795][2] = r_cell_wire[795];							inform_R[796][2] = r_cell_wire[796];							inform_R[798][2] = r_cell_wire[797];							inform_R[797][2] = r_cell_wire[798];							inform_R[799][2] = r_cell_wire[799];							inform_R[800][2] = r_cell_wire[800];							inform_R[802][2] = r_cell_wire[801];							inform_R[801][2] = r_cell_wire[802];							inform_R[803][2] = r_cell_wire[803];							inform_R[804][2] = r_cell_wire[804];							inform_R[806][2] = r_cell_wire[805];							inform_R[805][2] = r_cell_wire[806];							inform_R[807][2] = r_cell_wire[807];							inform_R[808][2] = r_cell_wire[808];							inform_R[810][2] = r_cell_wire[809];							inform_R[809][2] = r_cell_wire[810];							inform_R[811][2] = r_cell_wire[811];							inform_R[812][2] = r_cell_wire[812];							inform_R[814][2] = r_cell_wire[813];							inform_R[813][2] = r_cell_wire[814];							inform_R[815][2] = r_cell_wire[815];							inform_R[816][2] = r_cell_wire[816];							inform_R[818][2] = r_cell_wire[817];							inform_R[817][2] = r_cell_wire[818];							inform_R[819][2] = r_cell_wire[819];							inform_R[820][2] = r_cell_wire[820];							inform_R[822][2] = r_cell_wire[821];							inform_R[821][2] = r_cell_wire[822];							inform_R[823][2] = r_cell_wire[823];							inform_R[824][2] = r_cell_wire[824];							inform_R[826][2] = r_cell_wire[825];							inform_R[825][2] = r_cell_wire[826];							inform_R[827][2] = r_cell_wire[827];							inform_R[828][2] = r_cell_wire[828];							inform_R[830][2] = r_cell_wire[829];							inform_R[829][2] = r_cell_wire[830];							inform_R[831][2] = r_cell_wire[831];							inform_R[832][2] = r_cell_wire[832];							inform_R[834][2] = r_cell_wire[833];							inform_R[833][2] = r_cell_wire[834];							inform_R[835][2] = r_cell_wire[835];							inform_R[836][2] = r_cell_wire[836];							inform_R[838][2] = r_cell_wire[837];							inform_R[837][2] = r_cell_wire[838];							inform_R[839][2] = r_cell_wire[839];							inform_R[840][2] = r_cell_wire[840];							inform_R[842][2] = r_cell_wire[841];							inform_R[841][2] = r_cell_wire[842];							inform_R[843][2] = r_cell_wire[843];							inform_R[844][2] = r_cell_wire[844];							inform_R[846][2] = r_cell_wire[845];							inform_R[845][2] = r_cell_wire[846];							inform_R[847][2] = r_cell_wire[847];							inform_R[848][2] = r_cell_wire[848];							inform_R[850][2] = r_cell_wire[849];							inform_R[849][2] = r_cell_wire[850];							inform_R[851][2] = r_cell_wire[851];							inform_R[852][2] = r_cell_wire[852];							inform_R[854][2] = r_cell_wire[853];							inform_R[853][2] = r_cell_wire[854];							inform_R[855][2] = r_cell_wire[855];							inform_R[856][2] = r_cell_wire[856];							inform_R[858][2] = r_cell_wire[857];							inform_R[857][2] = r_cell_wire[858];							inform_R[859][2] = r_cell_wire[859];							inform_R[860][2] = r_cell_wire[860];							inform_R[862][2] = r_cell_wire[861];							inform_R[861][2] = r_cell_wire[862];							inform_R[863][2] = r_cell_wire[863];							inform_R[864][2] = r_cell_wire[864];							inform_R[866][2] = r_cell_wire[865];							inform_R[865][2] = r_cell_wire[866];							inform_R[867][2] = r_cell_wire[867];							inform_R[868][2] = r_cell_wire[868];							inform_R[870][2] = r_cell_wire[869];							inform_R[869][2] = r_cell_wire[870];							inform_R[871][2] = r_cell_wire[871];							inform_R[872][2] = r_cell_wire[872];							inform_R[874][2] = r_cell_wire[873];							inform_R[873][2] = r_cell_wire[874];							inform_R[875][2] = r_cell_wire[875];							inform_R[876][2] = r_cell_wire[876];							inform_R[878][2] = r_cell_wire[877];							inform_R[877][2] = r_cell_wire[878];							inform_R[879][2] = r_cell_wire[879];							inform_R[880][2] = r_cell_wire[880];							inform_R[882][2] = r_cell_wire[881];							inform_R[881][2] = r_cell_wire[882];							inform_R[883][2] = r_cell_wire[883];							inform_R[884][2] = r_cell_wire[884];							inform_R[886][2] = r_cell_wire[885];							inform_R[885][2] = r_cell_wire[886];							inform_R[887][2] = r_cell_wire[887];							inform_R[888][2] = r_cell_wire[888];							inform_R[890][2] = r_cell_wire[889];							inform_R[889][2] = r_cell_wire[890];							inform_R[891][2] = r_cell_wire[891];							inform_R[892][2] = r_cell_wire[892];							inform_R[894][2] = r_cell_wire[893];							inform_R[893][2] = r_cell_wire[894];							inform_R[895][2] = r_cell_wire[895];							inform_R[896][2] = r_cell_wire[896];							inform_R[898][2] = r_cell_wire[897];							inform_R[897][2] = r_cell_wire[898];							inform_R[899][2] = r_cell_wire[899];							inform_R[900][2] = r_cell_wire[900];							inform_R[902][2] = r_cell_wire[901];							inform_R[901][2] = r_cell_wire[902];							inform_R[903][2] = r_cell_wire[903];							inform_R[904][2] = r_cell_wire[904];							inform_R[906][2] = r_cell_wire[905];							inform_R[905][2] = r_cell_wire[906];							inform_R[907][2] = r_cell_wire[907];							inform_R[908][2] = r_cell_wire[908];							inform_R[910][2] = r_cell_wire[909];							inform_R[909][2] = r_cell_wire[910];							inform_R[911][2] = r_cell_wire[911];							inform_R[912][2] = r_cell_wire[912];							inform_R[914][2] = r_cell_wire[913];							inform_R[913][2] = r_cell_wire[914];							inform_R[915][2] = r_cell_wire[915];							inform_R[916][2] = r_cell_wire[916];							inform_R[918][2] = r_cell_wire[917];							inform_R[917][2] = r_cell_wire[918];							inform_R[919][2] = r_cell_wire[919];							inform_R[920][2] = r_cell_wire[920];							inform_R[922][2] = r_cell_wire[921];							inform_R[921][2] = r_cell_wire[922];							inform_R[923][2] = r_cell_wire[923];							inform_R[924][2] = r_cell_wire[924];							inform_R[926][2] = r_cell_wire[925];							inform_R[925][2] = r_cell_wire[926];							inform_R[927][2] = r_cell_wire[927];							inform_R[928][2] = r_cell_wire[928];							inform_R[930][2] = r_cell_wire[929];							inform_R[929][2] = r_cell_wire[930];							inform_R[931][2] = r_cell_wire[931];							inform_R[932][2] = r_cell_wire[932];							inform_R[934][2] = r_cell_wire[933];							inform_R[933][2] = r_cell_wire[934];							inform_R[935][2] = r_cell_wire[935];							inform_R[936][2] = r_cell_wire[936];							inform_R[938][2] = r_cell_wire[937];							inform_R[937][2] = r_cell_wire[938];							inform_R[939][2] = r_cell_wire[939];							inform_R[940][2] = r_cell_wire[940];							inform_R[942][2] = r_cell_wire[941];							inform_R[941][2] = r_cell_wire[942];							inform_R[943][2] = r_cell_wire[943];							inform_R[944][2] = r_cell_wire[944];							inform_R[946][2] = r_cell_wire[945];							inform_R[945][2] = r_cell_wire[946];							inform_R[947][2] = r_cell_wire[947];							inform_R[948][2] = r_cell_wire[948];							inform_R[950][2] = r_cell_wire[949];							inform_R[949][2] = r_cell_wire[950];							inform_R[951][2] = r_cell_wire[951];							inform_R[952][2] = r_cell_wire[952];							inform_R[954][2] = r_cell_wire[953];							inform_R[953][2] = r_cell_wire[954];							inform_R[955][2] = r_cell_wire[955];							inform_R[956][2] = r_cell_wire[956];							inform_R[958][2] = r_cell_wire[957];							inform_R[957][2] = r_cell_wire[958];							inform_R[959][2] = r_cell_wire[959];							inform_R[960][2] = r_cell_wire[960];							inform_R[962][2] = r_cell_wire[961];							inform_R[961][2] = r_cell_wire[962];							inform_R[963][2] = r_cell_wire[963];							inform_R[964][2] = r_cell_wire[964];							inform_R[966][2] = r_cell_wire[965];							inform_R[965][2] = r_cell_wire[966];							inform_R[967][2] = r_cell_wire[967];							inform_R[968][2] = r_cell_wire[968];							inform_R[970][2] = r_cell_wire[969];							inform_R[969][2] = r_cell_wire[970];							inform_R[971][2] = r_cell_wire[971];							inform_R[972][2] = r_cell_wire[972];							inform_R[974][2] = r_cell_wire[973];							inform_R[973][2] = r_cell_wire[974];							inform_R[975][2] = r_cell_wire[975];							inform_R[976][2] = r_cell_wire[976];							inform_R[978][2] = r_cell_wire[977];							inform_R[977][2] = r_cell_wire[978];							inform_R[979][2] = r_cell_wire[979];							inform_R[980][2] = r_cell_wire[980];							inform_R[982][2] = r_cell_wire[981];							inform_R[981][2] = r_cell_wire[982];							inform_R[983][2] = r_cell_wire[983];							inform_R[984][2] = r_cell_wire[984];							inform_R[986][2] = r_cell_wire[985];							inform_R[985][2] = r_cell_wire[986];							inform_R[987][2] = r_cell_wire[987];							inform_R[988][2] = r_cell_wire[988];							inform_R[990][2] = r_cell_wire[989];							inform_R[989][2] = r_cell_wire[990];							inform_R[991][2] = r_cell_wire[991];							inform_R[992][2] = r_cell_wire[992];							inform_R[994][2] = r_cell_wire[993];							inform_R[993][2] = r_cell_wire[994];							inform_R[995][2] = r_cell_wire[995];							inform_R[996][2] = r_cell_wire[996];							inform_R[998][2] = r_cell_wire[997];							inform_R[997][2] = r_cell_wire[998];							inform_R[999][2] = r_cell_wire[999];							inform_R[1000][2] = r_cell_wire[1000];							inform_R[1002][2] = r_cell_wire[1001];							inform_R[1001][2] = r_cell_wire[1002];							inform_R[1003][2] = r_cell_wire[1003];							inform_R[1004][2] = r_cell_wire[1004];							inform_R[1006][2] = r_cell_wire[1005];							inform_R[1005][2] = r_cell_wire[1006];							inform_R[1007][2] = r_cell_wire[1007];							inform_R[1008][2] = r_cell_wire[1008];							inform_R[1010][2] = r_cell_wire[1009];							inform_R[1009][2] = r_cell_wire[1010];							inform_R[1011][2] = r_cell_wire[1011];							inform_R[1012][2] = r_cell_wire[1012];							inform_R[1014][2] = r_cell_wire[1013];							inform_R[1013][2] = r_cell_wire[1014];							inform_R[1015][2] = r_cell_wire[1015];							inform_R[1016][2] = r_cell_wire[1016];							inform_R[1018][2] = r_cell_wire[1017];							inform_R[1017][2] = r_cell_wire[1018];							inform_R[1019][2] = r_cell_wire[1019];							inform_R[1020][2] = r_cell_wire[1020];							inform_R[1022][2] = r_cell_wire[1021];							inform_R[1021][2] = r_cell_wire[1022];							inform_R[1023][2] = r_cell_wire[1023];							inform_L[0][1] = l_cell_wire[0];							inform_L[2][1] = l_cell_wire[1];							inform_L[1][1] = l_cell_wire[2];							inform_L[3][1] = l_cell_wire[3];							inform_L[4][1] = l_cell_wire[4];							inform_L[6][1] = l_cell_wire[5];							inform_L[5][1] = l_cell_wire[6];							inform_L[7][1] = l_cell_wire[7];							inform_L[8][1] = l_cell_wire[8];							inform_L[10][1] = l_cell_wire[9];							inform_L[9][1] = l_cell_wire[10];							inform_L[11][1] = l_cell_wire[11];							inform_L[12][1] = l_cell_wire[12];							inform_L[14][1] = l_cell_wire[13];							inform_L[13][1] = l_cell_wire[14];							inform_L[15][1] = l_cell_wire[15];							inform_L[16][1] = l_cell_wire[16];							inform_L[18][1] = l_cell_wire[17];							inform_L[17][1] = l_cell_wire[18];							inform_L[19][1] = l_cell_wire[19];							inform_L[20][1] = l_cell_wire[20];							inform_L[22][1] = l_cell_wire[21];							inform_L[21][1] = l_cell_wire[22];							inform_L[23][1] = l_cell_wire[23];							inform_L[24][1] = l_cell_wire[24];							inform_L[26][1] = l_cell_wire[25];							inform_L[25][1] = l_cell_wire[26];							inform_L[27][1] = l_cell_wire[27];							inform_L[28][1] = l_cell_wire[28];							inform_L[30][1] = l_cell_wire[29];							inform_L[29][1] = l_cell_wire[30];							inform_L[31][1] = l_cell_wire[31];							inform_L[32][1] = l_cell_wire[32];							inform_L[34][1] = l_cell_wire[33];							inform_L[33][1] = l_cell_wire[34];							inform_L[35][1] = l_cell_wire[35];							inform_L[36][1] = l_cell_wire[36];							inform_L[38][1] = l_cell_wire[37];							inform_L[37][1] = l_cell_wire[38];							inform_L[39][1] = l_cell_wire[39];							inform_L[40][1] = l_cell_wire[40];							inform_L[42][1] = l_cell_wire[41];							inform_L[41][1] = l_cell_wire[42];							inform_L[43][1] = l_cell_wire[43];							inform_L[44][1] = l_cell_wire[44];							inform_L[46][1] = l_cell_wire[45];							inform_L[45][1] = l_cell_wire[46];							inform_L[47][1] = l_cell_wire[47];							inform_L[48][1] = l_cell_wire[48];							inform_L[50][1] = l_cell_wire[49];							inform_L[49][1] = l_cell_wire[50];							inform_L[51][1] = l_cell_wire[51];							inform_L[52][1] = l_cell_wire[52];							inform_L[54][1] = l_cell_wire[53];							inform_L[53][1] = l_cell_wire[54];							inform_L[55][1] = l_cell_wire[55];							inform_L[56][1] = l_cell_wire[56];							inform_L[58][1] = l_cell_wire[57];							inform_L[57][1] = l_cell_wire[58];							inform_L[59][1] = l_cell_wire[59];							inform_L[60][1] = l_cell_wire[60];							inform_L[62][1] = l_cell_wire[61];							inform_L[61][1] = l_cell_wire[62];							inform_L[63][1] = l_cell_wire[63];							inform_L[64][1] = l_cell_wire[64];							inform_L[66][1] = l_cell_wire[65];							inform_L[65][1] = l_cell_wire[66];							inform_L[67][1] = l_cell_wire[67];							inform_L[68][1] = l_cell_wire[68];							inform_L[70][1] = l_cell_wire[69];							inform_L[69][1] = l_cell_wire[70];							inform_L[71][1] = l_cell_wire[71];							inform_L[72][1] = l_cell_wire[72];							inform_L[74][1] = l_cell_wire[73];							inform_L[73][1] = l_cell_wire[74];							inform_L[75][1] = l_cell_wire[75];							inform_L[76][1] = l_cell_wire[76];							inform_L[78][1] = l_cell_wire[77];							inform_L[77][1] = l_cell_wire[78];							inform_L[79][1] = l_cell_wire[79];							inform_L[80][1] = l_cell_wire[80];							inform_L[82][1] = l_cell_wire[81];							inform_L[81][1] = l_cell_wire[82];							inform_L[83][1] = l_cell_wire[83];							inform_L[84][1] = l_cell_wire[84];							inform_L[86][1] = l_cell_wire[85];							inform_L[85][1] = l_cell_wire[86];							inform_L[87][1] = l_cell_wire[87];							inform_L[88][1] = l_cell_wire[88];							inform_L[90][1] = l_cell_wire[89];							inform_L[89][1] = l_cell_wire[90];							inform_L[91][1] = l_cell_wire[91];							inform_L[92][1] = l_cell_wire[92];							inform_L[94][1] = l_cell_wire[93];							inform_L[93][1] = l_cell_wire[94];							inform_L[95][1] = l_cell_wire[95];							inform_L[96][1] = l_cell_wire[96];							inform_L[98][1] = l_cell_wire[97];							inform_L[97][1] = l_cell_wire[98];							inform_L[99][1] = l_cell_wire[99];							inform_L[100][1] = l_cell_wire[100];							inform_L[102][1] = l_cell_wire[101];							inform_L[101][1] = l_cell_wire[102];							inform_L[103][1] = l_cell_wire[103];							inform_L[104][1] = l_cell_wire[104];							inform_L[106][1] = l_cell_wire[105];							inform_L[105][1] = l_cell_wire[106];							inform_L[107][1] = l_cell_wire[107];							inform_L[108][1] = l_cell_wire[108];							inform_L[110][1] = l_cell_wire[109];							inform_L[109][1] = l_cell_wire[110];							inform_L[111][1] = l_cell_wire[111];							inform_L[112][1] = l_cell_wire[112];							inform_L[114][1] = l_cell_wire[113];							inform_L[113][1] = l_cell_wire[114];							inform_L[115][1] = l_cell_wire[115];							inform_L[116][1] = l_cell_wire[116];							inform_L[118][1] = l_cell_wire[117];							inform_L[117][1] = l_cell_wire[118];							inform_L[119][1] = l_cell_wire[119];							inform_L[120][1] = l_cell_wire[120];							inform_L[122][1] = l_cell_wire[121];							inform_L[121][1] = l_cell_wire[122];							inform_L[123][1] = l_cell_wire[123];							inform_L[124][1] = l_cell_wire[124];							inform_L[126][1] = l_cell_wire[125];							inform_L[125][1] = l_cell_wire[126];							inform_L[127][1] = l_cell_wire[127];							inform_L[128][1] = l_cell_wire[128];							inform_L[130][1] = l_cell_wire[129];							inform_L[129][1] = l_cell_wire[130];							inform_L[131][1] = l_cell_wire[131];							inform_L[132][1] = l_cell_wire[132];							inform_L[134][1] = l_cell_wire[133];							inform_L[133][1] = l_cell_wire[134];							inform_L[135][1] = l_cell_wire[135];							inform_L[136][1] = l_cell_wire[136];							inform_L[138][1] = l_cell_wire[137];							inform_L[137][1] = l_cell_wire[138];							inform_L[139][1] = l_cell_wire[139];							inform_L[140][1] = l_cell_wire[140];							inform_L[142][1] = l_cell_wire[141];							inform_L[141][1] = l_cell_wire[142];							inform_L[143][1] = l_cell_wire[143];							inform_L[144][1] = l_cell_wire[144];							inform_L[146][1] = l_cell_wire[145];							inform_L[145][1] = l_cell_wire[146];							inform_L[147][1] = l_cell_wire[147];							inform_L[148][1] = l_cell_wire[148];							inform_L[150][1] = l_cell_wire[149];							inform_L[149][1] = l_cell_wire[150];							inform_L[151][1] = l_cell_wire[151];							inform_L[152][1] = l_cell_wire[152];							inform_L[154][1] = l_cell_wire[153];							inform_L[153][1] = l_cell_wire[154];							inform_L[155][1] = l_cell_wire[155];							inform_L[156][1] = l_cell_wire[156];							inform_L[158][1] = l_cell_wire[157];							inform_L[157][1] = l_cell_wire[158];							inform_L[159][1] = l_cell_wire[159];							inform_L[160][1] = l_cell_wire[160];							inform_L[162][1] = l_cell_wire[161];							inform_L[161][1] = l_cell_wire[162];							inform_L[163][1] = l_cell_wire[163];							inform_L[164][1] = l_cell_wire[164];							inform_L[166][1] = l_cell_wire[165];							inform_L[165][1] = l_cell_wire[166];							inform_L[167][1] = l_cell_wire[167];							inform_L[168][1] = l_cell_wire[168];							inform_L[170][1] = l_cell_wire[169];							inform_L[169][1] = l_cell_wire[170];							inform_L[171][1] = l_cell_wire[171];							inform_L[172][1] = l_cell_wire[172];							inform_L[174][1] = l_cell_wire[173];							inform_L[173][1] = l_cell_wire[174];							inform_L[175][1] = l_cell_wire[175];							inform_L[176][1] = l_cell_wire[176];							inform_L[178][1] = l_cell_wire[177];							inform_L[177][1] = l_cell_wire[178];							inform_L[179][1] = l_cell_wire[179];							inform_L[180][1] = l_cell_wire[180];							inform_L[182][1] = l_cell_wire[181];							inform_L[181][1] = l_cell_wire[182];							inform_L[183][1] = l_cell_wire[183];							inform_L[184][1] = l_cell_wire[184];							inform_L[186][1] = l_cell_wire[185];							inform_L[185][1] = l_cell_wire[186];							inform_L[187][1] = l_cell_wire[187];							inform_L[188][1] = l_cell_wire[188];							inform_L[190][1] = l_cell_wire[189];							inform_L[189][1] = l_cell_wire[190];							inform_L[191][1] = l_cell_wire[191];							inform_L[192][1] = l_cell_wire[192];							inform_L[194][1] = l_cell_wire[193];							inform_L[193][1] = l_cell_wire[194];							inform_L[195][1] = l_cell_wire[195];							inform_L[196][1] = l_cell_wire[196];							inform_L[198][1] = l_cell_wire[197];							inform_L[197][1] = l_cell_wire[198];							inform_L[199][1] = l_cell_wire[199];							inform_L[200][1] = l_cell_wire[200];							inform_L[202][1] = l_cell_wire[201];							inform_L[201][1] = l_cell_wire[202];							inform_L[203][1] = l_cell_wire[203];							inform_L[204][1] = l_cell_wire[204];							inform_L[206][1] = l_cell_wire[205];							inform_L[205][1] = l_cell_wire[206];							inform_L[207][1] = l_cell_wire[207];							inform_L[208][1] = l_cell_wire[208];							inform_L[210][1] = l_cell_wire[209];							inform_L[209][1] = l_cell_wire[210];							inform_L[211][1] = l_cell_wire[211];							inform_L[212][1] = l_cell_wire[212];							inform_L[214][1] = l_cell_wire[213];							inform_L[213][1] = l_cell_wire[214];							inform_L[215][1] = l_cell_wire[215];							inform_L[216][1] = l_cell_wire[216];							inform_L[218][1] = l_cell_wire[217];							inform_L[217][1] = l_cell_wire[218];							inform_L[219][1] = l_cell_wire[219];							inform_L[220][1] = l_cell_wire[220];							inform_L[222][1] = l_cell_wire[221];							inform_L[221][1] = l_cell_wire[222];							inform_L[223][1] = l_cell_wire[223];							inform_L[224][1] = l_cell_wire[224];							inform_L[226][1] = l_cell_wire[225];							inform_L[225][1] = l_cell_wire[226];							inform_L[227][1] = l_cell_wire[227];							inform_L[228][1] = l_cell_wire[228];							inform_L[230][1] = l_cell_wire[229];							inform_L[229][1] = l_cell_wire[230];							inform_L[231][1] = l_cell_wire[231];							inform_L[232][1] = l_cell_wire[232];							inform_L[234][1] = l_cell_wire[233];							inform_L[233][1] = l_cell_wire[234];							inform_L[235][1] = l_cell_wire[235];							inform_L[236][1] = l_cell_wire[236];							inform_L[238][1] = l_cell_wire[237];							inform_L[237][1] = l_cell_wire[238];							inform_L[239][1] = l_cell_wire[239];							inform_L[240][1] = l_cell_wire[240];							inform_L[242][1] = l_cell_wire[241];							inform_L[241][1] = l_cell_wire[242];							inform_L[243][1] = l_cell_wire[243];							inform_L[244][1] = l_cell_wire[244];							inform_L[246][1] = l_cell_wire[245];							inform_L[245][1] = l_cell_wire[246];							inform_L[247][1] = l_cell_wire[247];							inform_L[248][1] = l_cell_wire[248];							inform_L[250][1] = l_cell_wire[249];							inform_L[249][1] = l_cell_wire[250];							inform_L[251][1] = l_cell_wire[251];							inform_L[252][1] = l_cell_wire[252];							inform_L[254][1] = l_cell_wire[253];							inform_L[253][1] = l_cell_wire[254];							inform_L[255][1] = l_cell_wire[255];							inform_L[256][1] = l_cell_wire[256];							inform_L[258][1] = l_cell_wire[257];							inform_L[257][1] = l_cell_wire[258];							inform_L[259][1] = l_cell_wire[259];							inform_L[260][1] = l_cell_wire[260];							inform_L[262][1] = l_cell_wire[261];							inform_L[261][1] = l_cell_wire[262];							inform_L[263][1] = l_cell_wire[263];							inform_L[264][1] = l_cell_wire[264];							inform_L[266][1] = l_cell_wire[265];							inform_L[265][1] = l_cell_wire[266];							inform_L[267][1] = l_cell_wire[267];							inform_L[268][1] = l_cell_wire[268];							inform_L[270][1] = l_cell_wire[269];							inform_L[269][1] = l_cell_wire[270];							inform_L[271][1] = l_cell_wire[271];							inform_L[272][1] = l_cell_wire[272];							inform_L[274][1] = l_cell_wire[273];							inform_L[273][1] = l_cell_wire[274];							inform_L[275][1] = l_cell_wire[275];							inform_L[276][1] = l_cell_wire[276];							inform_L[278][1] = l_cell_wire[277];							inform_L[277][1] = l_cell_wire[278];							inform_L[279][1] = l_cell_wire[279];							inform_L[280][1] = l_cell_wire[280];							inform_L[282][1] = l_cell_wire[281];							inform_L[281][1] = l_cell_wire[282];							inform_L[283][1] = l_cell_wire[283];							inform_L[284][1] = l_cell_wire[284];							inform_L[286][1] = l_cell_wire[285];							inform_L[285][1] = l_cell_wire[286];							inform_L[287][1] = l_cell_wire[287];							inform_L[288][1] = l_cell_wire[288];							inform_L[290][1] = l_cell_wire[289];							inform_L[289][1] = l_cell_wire[290];							inform_L[291][1] = l_cell_wire[291];							inform_L[292][1] = l_cell_wire[292];							inform_L[294][1] = l_cell_wire[293];							inform_L[293][1] = l_cell_wire[294];							inform_L[295][1] = l_cell_wire[295];							inform_L[296][1] = l_cell_wire[296];							inform_L[298][1] = l_cell_wire[297];							inform_L[297][1] = l_cell_wire[298];							inform_L[299][1] = l_cell_wire[299];							inform_L[300][1] = l_cell_wire[300];							inform_L[302][1] = l_cell_wire[301];							inform_L[301][1] = l_cell_wire[302];							inform_L[303][1] = l_cell_wire[303];							inform_L[304][1] = l_cell_wire[304];							inform_L[306][1] = l_cell_wire[305];							inform_L[305][1] = l_cell_wire[306];							inform_L[307][1] = l_cell_wire[307];							inform_L[308][1] = l_cell_wire[308];							inform_L[310][1] = l_cell_wire[309];							inform_L[309][1] = l_cell_wire[310];							inform_L[311][1] = l_cell_wire[311];							inform_L[312][1] = l_cell_wire[312];							inform_L[314][1] = l_cell_wire[313];							inform_L[313][1] = l_cell_wire[314];							inform_L[315][1] = l_cell_wire[315];							inform_L[316][1] = l_cell_wire[316];							inform_L[318][1] = l_cell_wire[317];							inform_L[317][1] = l_cell_wire[318];							inform_L[319][1] = l_cell_wire[319];							inform_L[320][1] = l_cell_wire[320];							inform_L[322][1] = l_cell_wire[321];							inform_L[321][1] = l_cell_wire[322];							inform_L[323][1] = l_cell_wire[323];							inform_L[324][1] = l_cell_wire[324];							inform_L[326][1] = l_cell_wire[325];							inform_L[325][1] = l_cell_wire[326];							inform_L[327][1] = l_cell_wire[327];							inform_L[328][1] = l_cell_wire[328];							inform_L[330][1] = l_cell_wire[329];							inform_L[329][1] = l_cell_wire[330];							inform_L[331][1] = l_cell_wire[331];							inform_L[332][1] = l_cell_wire[332];							inform_L[334][1] = l_cell_wire[333];							inform_L[333][1] = l_cell_wire[334];							inform_L[335][1] = l_cell_wire[335];							inform_L[336][1] = l_cell_wire[336];							inform_L[338][1] = l_cell_wire[337];							inform_L[337][1] = l_cell_wire[338];							inform_L[339][1] = l_cell_wire[339];							inform_L[340][1] = l_cell_wire[340];							inform_L[342][1] = l_cell_wire[341];							inform_L[341][1] = l_cell_wire[342];							inform_L[343][1] = l_cell_wire[343];							inform_L[344][1] = l_cell_wire[344];							inform_L[346][1] = l_cell_wire[345];							inform_L[345][1] = l_cell_wire[346];							inform_L[347][1] = l_cell_wire[347];							inform_L[348][1] = l_cell_wire[348];							inform_L[350][1] = l_cell_wire[349];							inform_L[349][1] = l_cell_wire[350];							inform_L[351][1] = l_cell_wire[351];							inform_L[352][1] = l_cell_wire[352];							inform_L[354][1] = l_cell_wire[353];							inform_L[353][1] = l_cell_wire[354];							inform_L[355][1] = l_cell_wire[355];							inform_L[356][1] = l_cell_wire[356];							inform_L[358][1] = l_cell_wire[357];							inform_L[357][1] = l_cell_wire[358];							inform_L[359][1] = l_cell_wire[359];							inform_L[360][1] = l_cell_wire[360];							inform_L[362][1] = l_cell_wire[361];							inform_L[361][1] = l_cell_wire[362];							inform_L[363][1] = l_cell_wire[363];							inform_L[364][1] = l_cell_wire[364];							inform_L[366][1] = l_cell_wire[365];							inform_L[365][1] = l_cell_wire[366];							inform_L[367][1] = l_cell_wire[367];							inform_L[368][1] = l_cell_wire[368];							inform_L[370][1] = l_cell_wire[369];							inform_L[369][1] = l_cell_wire[370];							inform_L[371][1] = l_cell_wire[371];							inform_L[372][1] = l_cell_wire[372];							inform_L[374][1] = l_cell_wire[373];							inform_L[373][1] = l_cell_wire[374];							inform_L[375][1] = l_cell_wire[375];							inform_L[376][1] = l_cell_wire[376];							inform_L[378][1] = l_cell_wire[377];							inform_L[377][1] = l_cell_wire[378];							inform_L[379][1] = l_cell_wire[379];							inform_L[380][1] = l_cell_wire[380];							inform_L[382][1] = l_cell_wire[381];							inform_L[381][1] = l_cell_wire[382];							inform_L[383][1] = l_cell_wire[383];							inform_L[384][1] = l_cell_wire[384];							inform_L[386][1] = l_cell_wire[385];							inform_L[385][1] = l_cell_wire[386];							inform_L[387][1] = l_cell_wire[387];							inform_L[388][1] = l_cell_wire[388];							inform_L[390][1] = l_cell_wire[389];							inform_L[389][1] = l_cell_wire[390];							inform_L[391][1] = l_cell_wire[391];							inform_L[392][1] = l_cell_wire[392];							inform_L[394][1] = l_cell_wire[393];							inform_L[393][1] = l_cell_wire[394];							inform_L[395][1] = l_cell_wire[395];							inform_L[396][1] = l_cell_wire[396];							inform_L[398][1] = l_cell_wire[397];							inform_L[397][1] = l_cell_wire[398];							inform_L[399][1] = l_cell_wire[399];							inform_L[400][1] = l_cell_wire[400];							inform_L[402][1] = l_cell_wire[401];							inform_L[401][1] = l_cell_wire[402];							inform_L[403][1] = l_cell_wire[403];							inform_L[404][1] = l_cell_wire[404];							inform_L[406][1] = l_cell_wire[405];							inform_L[405][1] = l_cell_wire[406];							inform_L[407][1] = l_cell_wire[407];							inform_L[408][1] = l_cell_wire[408];							inform_L[410][1] = l_cell_wire[409];							inform_L[409][1] = l_cell_wire[410];							inform_L[411][1] = l_cell_wire[411];							inform_L[412][1] = l_cell_wire[412];							inform_L[414][1] = l_cell_wire[413];							inform_L[413][1] = l_cell_wire[414];							inform_L[415][1] = l_cell_wire[415];							inform_L[416][1] = l_cell_wire[416];							inform_L[418][1] = l_cell_wire[417];							inform_L[417][1] = l_cell_wire[418];							inform_L[419][1] = l_cell_wire[419];							inform_L[420][1] = l_cell_wire[420];							inform_L[422][1] = l_cell_wire[421];							inform_L[421][1] = l_cell_wire[422];							inform_L[423][1] = l_cell_wire[423];							inform_L[424][1] = l_cell_wire[424];							inform_L[426][1] = l_cell_wire[425];							inform_L[425][1] = l_cell_wire[426];							inform_L[427][1] = l_cell_wire[427];							inform_L[428][1] = l_cell_wire[428];							inform_L[430][1] = l_cell_wire[429];							inform_L[429][1] = l_cell_wire[430];							inform_L[431][1] = l_cell_wire[431];							inform_L[432][1] = l_cell_wire[432];							inform_L[434][1] = l_cell_wire[433];							inform_L[433][1] = l_cell_wire[434];							inform_L[435][1] = l_cell_wire[435];							inform_L[436][1] = l_cell_wire[436];							inform_L[438][1] = l_cell_wire[437];							inform_L[437][1] = l_cell_wire[438];							inform_L[439][1] = l_cell_wire[439];							inform_L[440][1] = l_cell_wire[440];							inform_L[442][1] = l_cell_wire[441];							inform_L[441][1] = l_cell_wire[442];							inform_L[443][1] = l_cell_wire[443];							inform_L[444][1] = l_cell_wire[444];							inform_L[446][1] = l_cell_wire[445];							inform_L[445][1] = l_cell_wire[446];							inform_L[447][1] = l_cell_wire[447];							inform_L[448][1] = l_cell_wire[448];							inform_L[450][1] = l_cell_wire[449];							inform_L[449][1] = l_cell_wire[450];							inform_L[451][1] = l_cell_wire[451];							inform_L[452][1] = l_cell_wire[452];							inform_L[454][1] = l_cell_wire[453];							inform_L[453][1] = l_cell_wire[454];							inform_L[455][1] = l_cell_wire[455];							inform_L[456][1] = l_cell_wire[456];							inform_L[458][1] = l_cell_wire[457];							inform_L[457][1] = l_cell_wire[458];							inform_L[459][1] = l_cell_wire[459];							inform_L[460][1] = l_cell_wire[460];							inform_L[462][1] = l_cell_wire[461];							inform_L[461][1] = l_cell_wire[462];							inform_L[463][1] = l_cell_wire[463];							inform_L[464][1] = l_cell_wire[464];							inform_L[466][1] = l_cell_wire[465];							inform_L[465][1] = l_cell_wire[466];							inform_L[467][1] = l_cell_wire[467];							inform_L[468][1] = l_cell_wire[468];							inform_L[470][1] = l_cell_wire[469];							inform_L[469][1] = l_cell_wire[470];							inform_L[471][1] = l_cell_wire[471];							inform_L[472][1] = l_cell_wire[472];							inform_L[474][1] = l_cell_wire[473];							inform_L[473][1] = l_cell_wire[474];							inform_L[475][1] = l_cell_wire[475];							inform_L[476][1] = l_cell_wire[476];							inform_L[478][1] = l_cell_wire[477];							inform_L[477][1] = l_cell_wire[478];							inform_L[479][1] = l_cell_wire[479];							inform_L[480][1] = l_cell_wire[480];							inform_L[482][1] = l_cell_wire[481];							inform_L[481][1] = l_cell_wire[482];							inform_L[483][1] = l_cell_wire[483];							inform_L[484][1] = l_cell_wire[484];							inform_L[486][1] = l_cell_wire[485];							inform_L[485][1] = l_cell_wire[486];							inform_L[487][1] = l_cell_wire[487];							inform_L[488][1] = l_cell_wire[488];							inform_L[490][1] = l_cell_wire[489];							inform_L[489][1] = l_cell_wire[490];							inform_L[491][1] = l_cell_wire[491];							inform_L[492][1] = l_cell_wire[492];							inform_L[494][1] = l_cell_wire[493];							inform_L[493][1] = l_cell_wire[494];							inform_L[495][1] = l_cell_wire[495];							inform_L[496][1] = l_cell_wire[496];							inform_L[498][1] = l_cell_wire[497];							inform_L[497][1] = l_cell_wire[498];							inform_L[499][1] = l_cell_wire[499];							inform_L[500][1] = l_cell_wire[500];							inform_L[502][1] = l_cell_wire[501];							inform_L[501][1] = l_cell_wire[502];							inform_L[503][1] = l_cell_wire[503];							inform_L[504][1] = l_cell_wire[504];							inform_L[506][1] = l_cell_wire[505];							inform_L[505][1] = l_cell_wire[506];							inform_L[507][1] = l_cell_wire[507];							inform_L[508][1] = l_cell_wire[508];							inform_L[510][1] = l_cell_wire[509];							inform_L[509][1] = l_cell_wire[510];							inform_L[511][1] = l_cell_wire[511];							inform_L[512][1] = l_cell_wire[512];							inform_L[514][1] = l_cell_wire[513];							inform_L[513][1] = l_cell_wire[514];							inform_L[515][1] = l_cell_wire[515];							inform_L[516][1] = l_cell_wire[516];							inform_L[518][1] = l_cell_wire[517];							inform_L[517][1] = l_cell_wire[518];							inform_L[519][1] = l_cell_wire[519];							inform_L[520][1] = l_cell_wire[520];							inform_L[522][1] = l_cell_wire[521];							inform_L[521][1] = l_cell_wire[522];							inform_L[523][1] = l_cell_wire[523];							inform_L[524][1] = l_cell_wire[524];							inform_L[526][1] = l_cell_wire[525];							inform_L[525][1] = l_cell_wire[526];							inform_L[527][1] = l_cell_wire[527];							inform_L[528][1] = l_cell_wire[528];							inform_L[530][1] = l_cell_wire[529];							inform_L[529][1] = l_cell_wire[530];							inform_L[531][1] = l_cell_wire[531];							inform_L[532][1] = l_cell_wire[532];							inform_L[534][1] = l_cell_wire[533];							inform_L[533][1] = l_cell_wire[534];							inform_L[535][1] = l_cell_wire[535];							inform_L[536][1] = l_cell_wire[536];							inform_L[538][1] = l_cell_wire[537];							inform_L[537][1] = l_cell_wire[538];							inform_L[539][1] = l_cell_wire[539];							inform_L[540][1] = l_cell_wire[540];							inform_L[542][1] = l_cell_wire[541];							inform_L[541][1] = l_cell_wire[542];							inform_L[543][1] = l_cell_wire[543];							inform_L[544][1] = l_cell_wire[544];							inform_L[546][1] = l_cell_wire[545];							inform_L[545][1] = l_cell_wire[546];							inform_L[547][1] = l_cell_wire[547];							inform_L[548][1] = l_cell_wire[548];							inform_L[550][1] = l_cell_wire[549];							inform_L[549][1] = l_cell_wire[550];							inform_L[551][1] = l_cell_wire[551];							inform_L[552][1] = l_cell_wire[552];							inform_L[554][1] = l_cell_wire[553];							inform_L[553][1] = l_cell_wire[554];							inform_L[555][1] = l_cell_wire[555];							inform_L[556][1] = l_cell_wire[556];							inform_L[558][1] = l_cell_wire[557];							inform_L[557][1] = l_cell_wire[558];							inform_L[559][1] = l_cell_wire[559];							inform_L[560][1] = l_cell_wire[560];							inform_L[562][1] = l_cell_wire[561];							inform_L[561][1] = l_cell_wire[562];							inform_L[563][1] = l_cell_wire[563];							inform_L[564][1] = l_cell_wire[564];							inform_L[566][1] = l_cell_wire[565];							inform_L[565][1] = l_cell_wire[566];							inform_L[567][1] = l_cell_wire[567];							inform_L[568][1] = l_cell_wire[568];							inform_L[570][1] = l_cell_wire[569];							inform_L[569][1] = l_cell_wire[570];							inform_L[571][1] = l_cell_wire[571];							inform_L[572][1] = l_cell_wire[572];							inform_L[574][1] = l_cell_wire[573];							inform_L[573][1] = l_cell_wire[574];							inform_L[575][1] = l_cell_wire[575];							inform_L[576][1] = l_cell_wire[576];							inform_L[578][1] = l_cell_wire[577];							inform_L[577][1] = l_cell_wire[578];							inform_L[579][1] = l_cell_wire[579];							inform_L[580][1] = l_cell_wire[580];							inform_L[582][1] = l_cell_wire[581];							inform_L[581][1] = l_cell_wire[582];							inform_L[583][1] = l_cell_wire[583];							inform_L[584][1] = l_cell_wire[584];							inform_L[586][1] = l_cell_wire[585];							inform_L[585][1] = l_cell_wire[586];							inform_L[587][1] = l_cell_wire[587];							inform_L[588][1] = l_cell_wire[588];							inform_L[590][1] = l_cell_wire[589];							inform_L[589][1] = l_cell_wire[590];							inform_L[591][1] = l_cell_wire[591];							inform_L[592][1] = l_cell_wire[592];							inform_L[594][1] = l_cell_wire[593];							inform_L[593][1] = l_cell_wire[594];							inform_L[595][1] = l_cell_wire[595];							inform_L[596][1] = l_cell_wire[596];							inform_L[598][1] = l_cell_wire[597];							inform_L[597][1] = l_cell_wire[598];							inform_L[599][1] = l_cell_wire[599];							inform_L[600][1] = l_cell_wire[600];							inform_L[602][1] = l_cell_wire[601];							inform_L[601][1] = l_cell_wire[602];							inform_L[603][1] = l_cell_wire[603];							inform_L[604][1] = l_cell_wire[604];							inform_L[606][1] = l_cell_wire[605];							inform_L[605][1] = l_cell_wire[606];							inform_L[607][1] = l_cell_wire[607];							inform_L[608][1] = l_cell_wire[608];							inform_L[610][1] = l_cell_wire[609];							inform_L[609][1] = l_cell_wire[610];							inform_L[611][1] = l_cell_wire[611];							inform_L[612][1] = l_cell_wire[612];							inform_L[614][1] = l_cell_wire[613];							inform_L[613][1] = l_cell_wire[614];							inform_L[615][1] = l_cell_wire[615];							inform_L[616][1] = l_cell_wire[616];							inform_L[618][1] = l_cell_wire[617];							inform_L[617][1] = l_cell_wire[618];							inform_L[619][1] = l_cell_wire[619];							inform_L[620][1] = l_cell_wire[620];							inform_L[622][1] = l_cell_wire[621];							inform_L[621][1] = l_cell_wire[622];							inform_L[623][1] = l_cell_wire[623];							inform_L[624][1] = l_cell_wire[624];							inform_L[626][1] = l_cell_wire[625];							inform_L[625][1] = l_cell_wire[626];							inform_L[627][1] = l_cell_wire[627];							inform_L[628][1] = l_cell_wire[628];							inform_L[630][1] = l_cell_wire[629];							inform_L[629][1] = l_cell_wire[630];							inform_L[631][1] = l_cell_wire[631];							inform_L[632][1] = l_cell_wire[632];							inform_L[634][1] = l_cell_wire[633];							inform_L[633][1] = l_cell_wire[634];							inform_L[635][1] = l_cell_wire[635];							inform_L[636][1] = l_cell_wire[636];							inform_L[638][1] = l_cell_wire[637];							inform_L[637][1] = l_cell_wire[638];							inform_L[639][1] = l_cell_wire[639];							inform_L[640][1] = l_cell_wire[640];							inform_L[642][1] = l_cell_wire[641];							inform_L[641][1] = l_cell_wire[642];							inform_L[643][1] = l_cell_wire[643];							inform_L[644][1] = l_cell_wire[644];							inform_L[646][1] = l_cell_wire[645];							inform_L[645][1] = l_cell_wire[646];							inform_L[647][1] = l_cell_wire[647];							inform_L[648][1] = l_cell_wire[648];							inform_L[650][1] = l_cell_wire[649];							inform_L[649][1] = l_cell_wire[650];							inform_L[651][1] = l_cell_wire[651];							inform_L[652][1] = l_cell_wire[652];							inform_L[654][1] = l_cell_wire[653];							inform_L[653][1] = l_cell_wire[654];							inform_L[655][1] = l_cell_wire[655];							inform_L[656][1] = l_cell_wire[656];							inform_L[658][1] = l_cell_wire[657];							inform_L[657][1] = l_cell_wire[658];							inform_L[659][1] = l_cell_wire[659];							inform_L[660][1] = l_cell_wire[660];							inform_L[662][1] = l_cell_wire[661];							inform_L[661][1] = l_cell_wire[662];							inform_L[663][1] = l_cell_wire[663];							inform_L[664][1] = l_cell_wire[664];							inform_L[666][1] = l_cell_wire[665];							inform_L[665][1] = l_cell_wire[666];							inform_L[667][1] = l_cell_wire[667];							inform_L[668][1] = l_cell_wire[668];							inform_L[670][1] = l_cell_wire[669];							inform_L[669][1] = l_cell_wire[670];							inform_L[671][1] = l_cell_wire[671];							inform_L[672][1] = l_cell_wire[672];							inform_L[674][1] = l_cell_wire[673];							inform_L[673][1] = l_cell_wire[674];							inform_L[675][1] = l_cell_wire[675];							inform_L[676][1] = l_cell_wire[676];							inform_L[678][1] = l_cell_wire[677];							inform_L[677][1] = l_cell_wire[678];							inform_L[679][1] = l_cell_wire[679];							inform_L[680][1] = l_cell_wire[680];							inform_L[682][1] = l_cell_wire[681];							inform_L[681][1] = l_cell_wire[682];							inform_L[683][1] = l_cell_wire[683];							inform_L[684][1] = l_cell_wire[684];							inform_L[686][1] = l_cell_wire[685];							inform_L[685][1] = l_cell_wire[686];							inform_L[687][1] = l_cell_wire[687];							inform_L[688][1] = l_cell_wire[688];							inform_L[690][1] = l_cell_wire[689];							inform_L[689][1] = l_cell_wire[690];							inform_L[691][1] = l_cell_wire[691];							inform_L[692][1] = l_cell_wire[692];							inform_L[694][1] = l_cell_wire[693];							inform_L[693][1] = l_cell_wire[694];							inform_L[695][1] = l_cell_wire[695];							inform_L[696][1] = l_cell_wire[696];							inform_L[698][1] = l_cell_wire[697];							inform_L[697][1] = l_cell_wire[698];							inform_L[699][1] = l_cell_wire[699];							inform_L[700][1] = l_cell_wire[700];							inform_L[702][1] = l_cell_wire[701];							inform_L[701][1] = l_cell_wire[702];							inform_L[703][1] = l_cell_wire[703];							inform_L[704][1] = l_cell_wire[704];							inform_L[706][1] = l_cell_wire[705];							inform_L[705][1] = l_cell_wire[706];							inform_L[707][1] = l_cell_wire[707];							inform_L[708][1] = l_cell_wire[708];							inform_L[710][1] = l_cell_wire[709];							inform_L[709][1] = l_cell_wire[710];							inform_L[711][1] = l_cell_wire[711];							inform_L[712][1] = l_cell_wire[712];							inform_L[714][1] = l_cell_wire[713];							inform_L[713][1] = l_cell_wire[714];							inform_L[715][1] = l_cell_wire[715];							inform_L[716][1] = l_cell_wire[716];							inform_L[718][1] = l_cell_wire[717];							inform_L[717][1] = l_cell_wire[718];							inform_L[719][1] = l_cell_wire[719];							inform_L[720][1] = l_cell_wire[720];							inform_L[722][1] = l_cell_wire[721];							inform_L[721][1] = l_cell_wire[722];							inform_L[723][1] = l_cell_wire[723];							inform_L[724][1] = l_cell_wire[724];							inform_L[726][1] = l_cell_wire[725];							inform_L[725][1] = l_cell_wire[726];							inform_L[727][1] = l_cell_wire[727];							inform_L[728][1] = l_cell_wire[728];							inform_L[730][1] = l_cell_wire[729];							inform_L[729][1] = l_cell_wire[730];							inform_L[731][1] = l_cell_wire[731];							inform_L[732][1] = l_cell_wire[732];							inform_L[734][1] = l_cell_wire[733];							inform_L[733][1] = l_cell_wire[734];							inform_L[735][1] = l_cell_wire[735];							inform_L[736][1] = l_cell_wire[736];							inform_L[738][1] = l_cell_wire[737];							inform_L[737][1] = l_cell_wire[738];							inform_L[739][1] = l_cell_wire[739];							inform_L[740][1] = l_cell_wire[740];							inform_L[742][1] = l_cell_wire[741];							inform_L[741][1] = l_cell_wire[742];							inform_L[743][1] = l_cell_wire[743];							inform_L[744][1] = l_cell_wire[744];							inform_L[746][1] = l_cell_wire[745];							inform_L[745][1] = l_cell_wire[746];							inform_L[747][1] = l_cell_wire[747];							inform_L[748][1] = l_cell_wire[748];							inform_L[750][1] = l_cell_wire[749];							inform_L[749][1] = l_cell_wire[750];							inform_L[751][1] = l_cell_wire[751];							inform_L[752][1] = l_cell_wire[752];							inform_L[754][1] = l_cell_wire[753];							inform_L[753][1] = l_cell_wire[754];							inform_L[755][1] = l_cell_wire[755];							inform_L[756][1] = l_cell_wire[756];							inform_L[758][1] = l_cell_wire[757];							inform_L[757][1] = l_cell_wire[758];							inform_L[759][1] = l_cell_wire[759];							inform_L[760][1] = l_cell_wire[760];							inform_L[762][1] = l_cell_wire[761];							inform_L[761][1] = l_cell_wire[762];							inform_L[763][1] = l_cell_wire[763];							inform_L[764][1] = l_cell_wire[764];							inform_L[766][1] = l_cell_wire[765];							inform_L[765][1] = l_cell_wire[766];							inform_L[767][1] = l_cell_wire[767];							inform_L[768][1] = l_cell_wire[768];							inform_L[770][1] = l_cell_wire[769];							inform_L[769][1] = l_cell_wire[770];							inform_L[771][1] = l_cell_wire[771];							inform_L[772][1] = l_cell_wire[772];							inform_L[774][1] = l_cell_wire[773];							inform_L[773][1] = l_cell_wire[774];							inform_L[775][1] = l_cell_wire[775];							inform_L[776][1] = l_cell_wire[776];							inform_L[778][1] = l_cell_wire[777];							inform_L[777][1] = l_cell_wire[778];							inform_L[779][1] = l_cell_wire[779];							inform_L[780][1] = l_cell_wire[780];							inform_L[782][1] = l_cell_wire[781];							inform_L[781][1] = l_cell_wire[782];							inform_L[783][1] = l_cell_wire[783];							inform_L[784][1] = l_cell_wire[784];							inform_L[786][1] = l_cell_wire[785];							inform_L[785][1] = l_cell_wire[786];							inform_L[787][1] = l_cell_wire[787];							inform_L[788][1] = l_cell_wire[788];							inform_L[790][1] = l_cell_wire[789];							inform_L[789][1] = l_cell_wire[790];							inform_L[791][1] = l_cell_wire[791];							inform_L[792][1] = l_cell_wire[792];							inform_L[794][1] = l_cell_wire[793];							inform_L[793][1] = l_cell_wire[794];							inform_L[795][1] = l_cell_wire[795];							inform_L[796][1] = l_cell_wire[796];							inform_L[798][1] = l_cell_wire[797];							inform_L[797][1] = l_cell_wire[798];							inform_L[799][1] = l_cell_wire[799];							inform_L[800][1] = l_cell_wire[800];							inform_L[802][1] = l_cell_wire[801];							inform_L[801][1] = l_cell_wire[802];							inform_L[803][1] = l_cell_wire[803];							inform_L[804][1] = l_cell_wire[804];							inform_L[806][1] = l_cell_wire[805];							inform_L[805][1] = l_cell_wire[806];							inform_L[807][1] = l_cell_wire[807];							inform_L[808][1] = l_cell_wire[808];							inform_L[810][1] = l_cell_wire[809];							inform_L[809][1] = l_cell_wire[810];							inform_L[811][1] = l_cell_wire[811];							inform_L[812][1] = l_cell_wire[812];							inform_L[814][1] = l_cell_wire[813];							inform_L[813][1] = l_cell_wire[814];							inform_L[815][1] = l_cell_wire[815];							inform_L[816][1] = l_cell_wire[816];							inform_L[818][1] = l_cell_wire[817];							inform_L[817][1] = l_cell_wire[818];							inform_L[819][1] = l_cell_wire[819];							inform_L[820][1] = l_cell_wire[820];							inform_L[822][1] = l_cell_wire[821];							inform_L[821][1] = l_cell_wire[822];							inform_L[823][1] = l_cell_wire[823];							inform_L[824][1] = l_cell_wire[824];							inform_L[826][1] = l_cell_wire[825];							inform_L[825][1] = l_cell_wire[826];							inform_L[827][1] = l_cell_wire[827];							inform_L[828][1] = l_cell_wire[828];							inform_L[830][1] = l_cell_wire[829];							inform_L[829][1] = l_cell_wire[830];							inform_L[831][1] = l_cell_wire[831];							inform_L[832][1] = l_cell_wire[832];							inform_L[834][1] = l_cell_wire[833];							inform_L[833][1] = l_cell_wire[834];							inform_L[835][1] = l_cell_wire[835];							inform_L[836][1] = l_cell_wire[836];							inform_L[838][1] = l_cell_wire[837];							inform_L[837][1] = l_cell_wire[838];							inform_L[839][1] = l_cell_wire[839];							inform_L[840][1] = l_cell_wire[840];							inform_L[842][1] = l_cell_wire[841];							inform_L[841][1] = l_cell_wire[842];							inform_L[843][1] = l_cell_wire[843];							inform_L[844][1] = l_cell_wire[844];							inform_L[846][1] = l_cell_wire[845];							inform_L[845][1] = l_cell_wire[846];							inform_L[847][1] = l_cell_wire[847];							inform_L[848][1] = l_cell_wire[848];							inform_L[850][1] = l_cell_wire[849];							inform_L[849][1] = l_cell_wire[850];							inform_L[851][1] = l_cell_wire[851];							inform_L[852][1] = l_cell_wire[852];							inform_L[854][1] = l_cell_wire[853];							inform_L[853][1] = l_cell_wire[854];							inform_L[855][1] = l_cell_wire[855];							inform_L[856][1] = l_cell_wire[856];							inform_L[858][1] = l_cell_wire[857];							inform_L[857][1] = l_cell_wire[858];							inform_L[859][1] = l_cell_wire[859];							inform_L[860][1] = l_cell_wire[860];							inform_L[862][1] = l_cell_wire[861];							inform_L[861][1] = l_cell_wire[862];							inform_L[863][1] = l_cell_wire[863];							inform_L[864][1] = l_cell_wire[864];							inform_L[866][1] = l_cell_wire[865];							inform_L[865][1] = l_cell_wire[866];							inform_L[867][1] = l_cell_wire[867];							inform_L[868][1] = l_cell_wire[868];							inform_L[870][1] = l_cell_wire[869];							inform_L[869][1] = l_cell_wire[870];							inform_L[871][1] = l_cell_wire[871];							inform_L[872][1] = l_cell_wire[872];							inform_L[874][1] = l_cell_wire[873];							inform_L[873][1] = l_cell_wire[874];							inform_L[875][1] = l_cell_wire[875];							inform_L[876][1] = l_cell_wire[876];							inform_L[878][1] = l_cell_wire[877];							inform_L[877][1] = l_cell_wire[878];							inform_L[879][1] = l_cell_wire[879];							inform_L[880][1] = l_cell_wire[880];							inform_L[882][1] = l_cell_wire[881];							inform_L[881][1] = l_cell_wire[882];							inform_L[883][1] = l_cell_wire[883];							inform_L[884][1] = l_cell_wire[884];							inform_L[886][1] = l_cell_wire[885];							inform_L[885][1] = l_cell_wire[886];							inform_L[887][1] = l_cell_wire[887];							inform_L[888][1] = l_cell_wire[888];							inform_L[890][1] = l_cell_wire[889];							inform_L[889][1] = l_cell_wire[890];							inform_L[891][1] = l_cell_wire[891];							inform_L[892][1] = l_cell_wire[892];							inform_L[894][1] = l_cell_wire[893];							inform_L[893][1] = l_cell_wire[894];							inform_L[895][1] = l_cell_wire[895];							inform_L[896][1] = l_cell_wire[896];							inform_L[898][1] = l_cell_wire[897];							inform_L[897][1] = l_cell_wire[898];							inform_L[899][1] = l_cell_wire[899];							inform_L[900][1] = l_cell_wire[900];							inform_L[902][1] = l_cell_wire[901];							inform_L[901][1] = l_cell_wire[902];							inform_L[903][1] = l_cell_wire[903];							inform_L[904][1] = l_cell_wire[904];							inform_L[906][1] = l_cell_wire[905];							inform_L[905][1] = l_cell_wire[906];							inform_L[907][1] = l_cell_wire[907];							inform_L[908][1] = l_cell_wire[908];							inform_L[910][1] = l_cell_wire[909];							inform_L[909][1] = l_cell_wire[910];							inform_L[911][1] = l_cell_wire[911];							inform_L[912][1] = l_cell_wire[912];							inform_L[914][1] = l_cell_wire[913];							inform_L[913][1] = l_cell_wire[914];							inform_L[915][1] = l_cell_wire[915];							inform_L[916][1] = l_cell_wire[916];							inform_L[918][1] = l_cell_wire[917];							inform_L[917][1] = l_cell_wire[918];							inform_L[919][1] = l_cell_wire[919];							inform_L[920][1] = l_cell_wire[920];							inform_L[922][1] = l_cell_wire[921];							inform_L[921][1] = l_cell_wire[922];							inform_L[923][1] = l_cell_wire[923];							inform_L[924][1] = l_cell_wire[924];							inform_L[926][1] = l_cell_wire[925];							inform_L[925][1] = l_cell_wire[926];							inform_L[927][1] = l_cell_wire[927];							inform_L[928][1] = l_cell_wire[928];							inform_L[930][1] = l_cell_wire[929];							inform_L[929][1] = l_cell_wire[930];							inform_L[931][1] = l_cell_wire[931];							inform_L[932][1] = l_cell_wire[932];							inform_L[934][1] = l_cell_wire[933];							inform_L[933][1] = l_cell_wire[934];							inform_L[935][1] = l_cell_wire[935];							inform_L[936][1] = l_cell_wire[936];							inform_L[938][1] = l_cell_wire[937];							inform_L[937][1] = l_cell_wire[938];							inform_L[939][1] = l_cell_wire[939];							inform_L[940][1] = l_cell_wire[940];							inform_L[942][1] = l_cell_wire[941];							inform_L[941][1] = l_cell_wire[942];							inform_L[943][1] = l_cell_wire[943];							inform_L[944][1] = l_cell_wire[944];							inform_L[946][1] = l_cell_wire[945];							inform_L[945][1] = l_cell_wire[946];							inform_L[947][1] = l_cell_wire[947];							inform_L[948][1] = l_cell_wire[948];							inform_L[950][1] = l_cell_wire[949];							inform_L[949][1] = l_cell_wire[950];							inform_L[951][1] = l_cell_wire[951];							inform_L[952][1] = l_cell_wire[952];							inform_L[954][1] = l_cell_wire[953];							inform_L[953][1] = l_cell_wire[954];							inform_L[955][1] = l_cell_wire[955];							inform_L[956][1] = l_cell_wire[956];							inform_L[958][1] = l_cell_wire[957];							inform_L[957][1] = l_cell_wire[958];							inform_L[959][1] = l_cell_wire[959];							inform_L[960][1] = l_cell_wire[960];							inform_L[962][1] = l_cell_wire[961];							inform_L[961][1] = l_cell_wire[962];							inform_L[963][1] = l_cell_wire[963];							inform_L[964][1] = l_cell_wire[964];							inform_L[966][1] = l_cell_wire[965];							inform_L[965][1] = l_cell_wire[966];							inform_L[967][1] = l_cell_wire[967];							inform_L[968][1] = l_cell_wire[968];							inform_L[970][1] = l_cell_wire[969];							inform_L[969][1] = l_cell_wire[970];							inform_L[971][1] = l_cell_wire[971];							inform_L[972][1] = l_cell_wire[972];							inform_L[974][1] = l_cell_wire[973];							inform_L[973][1] = l_cell_wire[974];							inform_L[975][1] = l_cell_wire[975];							inform_L[976][1] = l_cell_wire[976];							inform_L[978][1] = l_cell_wire[977];							inform_L[977][1] = l_cell_wire[978];							inform_L[979][1] = l_cell_wire[979];							inform_L[980][1] = l_cell_wire[980];							inform_L[982][1] = l_cell_wire[981];							inform_L[981][1] = l_cell_wire[982];							inform_L[983][1] = l_cell_wire[983];							inform_L[984][1] = l_cell_wire[984];							inform_L[986][1] = l_cell_wire[985];							inform_L[985][1] = l_cell_wire[986];							inform_L[987][1] = l_cell_wire[987];							inform_L[988][1] = l_cell_wire[988];							inform_L[990][1] = l_cell_wire[989];							inform_L[989][1] = l_cell_wire[990];							inform_L[991][1] = l_cell_wire[991];							inform_L[992][1] = l_cell_wire[992];							inform_L[994][1] = l_cell_wire[993];							inform_L[993][1] = l_cell_wire[994];							inform_L[995][1] = l_cell_wire[995];							inform_L[996][1] = l_cell_wire[996];							inform_L[998][1] = l_cell_wire[997];							inform_L[997][1] = l_cell_wire[998];							inform_L[999][1] = l_cell_wire[999];							inform_L[1000][1] = l_cell_wire[1000];							inform_L[1002][1] = l_cell_wire[1001];							inform_L[1001][1] = l_cell_wire[1002];							inform_L[1003][1] = l_cell_wire[1003];							inform_L[1004][1] = l_cell_wire[1004];							inform_L[1006][1] = l_cell_wire[1005];							inform_L[1005][1] = l_cell_wire[1006];							inform_L[1007][1] = l_cell_wire[1007];							inform_L[1008][1] = l_cell_wire[1008];							inform_L[1010][1] = l_cell_wire[1009];							inform_L[1009][1] = l_cell_wire[1010];							inform_L[1011][1] = l_cell_wire[1011];							inform_L[1012][1] = l_cell_wire[1012];							inform_L[1014][1] = l_cell_wire[1013];							inform_L[1013][1] = l_cell_wire[1014];							inform_L[1015][1] = l_cell_wire[1015];							inform_L[1016][1] = l_cell_wire[1016];							inform_L[1018][1] = l_cell_wire[1017];							inform_L[1017][1] = l_cell_wire[1018];							inform_L[1019][1] = l_cell_wire[1019];							inform_L[1020][1] = l_cell_wire[1020];							inform_L[1022][1] = l_cell_wire[1021];							inform_L[1021][1] = l_cell_wire[1022];							inform_L[1023][1] = l_cell_wire[1023];						end
						3:						begin							inform_R[0][3] = r_cell_wire[0];							inform_R[4][3] = r_cell_wire[1];							inform_R[1][3] = r_cell_wire[2];							inform_R[5][3] = r_cell_wire[3];							inform_R[2][3] = r_cell_wire[4];							inform_R[6][3] = r_cell_wire[5];							inform_R[3][3] = r_cell_wire[6];							inform_R[7][3] = r_cell_wire[7];							inform_R[8][3] = r_cell_wire[8];							inform_R[12][3] = r_cell_wire[9];							inform_R[9][3] = r_cell_wire[10];							inform_R[13][3] = r_cell_wire[11];							inform_R[10][3] = r_cell_wire[12];							inform_R[14][3] = r_cell_wire[13];							inform_R[11][3] = r_cell_wire[14];							inform_R[15][3] = r_cell_wire[15];							inform_R[16][3] = r_cell_wire[16];							inform_R[20][3] = r_cell_wire[17];							inform_R[17][3] = r_cell_wire[18];							inform_R[21][3] = r_cell_wire[19];							inform_R[18][3] = r_cell_wire[20];							inform_R[22][3] = r_cell_wire[21];							inform_R[19][3] = r_cell_wire[22];							inform_R[23][3] = r_cell_wire[23];							inform_R[24][3] = r_cell_wire[24];							inform_R[28][3] = r_cell_wire[25];							inform_R[25][3] = r_cell_wire[26];							inform_R[29][3] = r_cell_wire[27];							inform_R[26][3] = r_cell_wire[28];							inform_R[30][3] = r_cell_wire[29];							inform_R[27][3] = r_cell_wire[30];							inform_R[31][3] = r_cell_wire[31];							inform_R[32][3] = r_cell_wire[32];							inform_R[36][3] = r_cell_wire[33];							inform_R[33][3] = r_cell_wire[34];							inform_R[37][3] = r_cell_wire[35];							inform_R[34][3] = r_cell_wire[36];							inform_R[38][3] = r_cell_wire[37];							inform_R[35][3] = r_cell_wire[38];							inform_R[39][3] = r_cell_wire[39];							inform_R[40][3] = r_cell_wire[40];							inform_R[44][3] = r_cell_wire[41];							inform_R[41][3] = r_cell_wire[42];							inform_R[45][3] = r_cell_wire[43];							inform_R[42][3] = r_cell_wire[44];							inform_R[46][3] = r_cell_wire[45];							inform_R[43][3] = r_cell_wire[46];							inform_R[47][3] = r_cell_wire[47];							inform_R[48][3] = r_cell_wire[48];							inform_R[52][3] = r_cell_wire[49];							inform_R[49][3] = r_cell_wire[50];							inform_R[53][3] = r_cell_wire[51];							inform_R[50][3] = r_cell_wire[52];							inform_R[54][3] = r_cell_wire[53];							inform_R[51][3] = r_cell_wire[54];							inform_R[55][3] = r_cell_wire[55];							inform_R[56][3] = r_cell_wire[56];							inform_R[60][3] = r_cell_wire[57];							inform_R[57][3] = r_cell_wire[58];							inform_R[61][3] = r_cell_wire[59];							inform_R[58][3] = r_cell_wire[60];							inform_R[62][3] = r_cell_wire[61];							inform_R[59][3] = r_cell_wire[62];							inform_R[63][3] = r_cell_wire[63];							inform_R[64][3] = r_cell_wire[64];							inform_R[68][3] = r_cell_wire[65];							inform_R[65][3] = r_cell_wire[66];							inform_R[69][3] = r_cell_wire[67];							inform_R[66][3] = r_cell_wire[68];							inform_R[70][3] = r_cell_wire[69];							inform_R[67][3] = r_cell_wire[70];							inform_R[71][3] = r_cell_wire[71];							inform_R[72][3] = r_cell_wire[72];							inform_R[76][3] = r_cell_wire[73];							inform_R[73][3] = r_cell_wire[74];							inform_R[77][3] = r_cell_wire[75];							inform_R[74][3] = r_cell_wire[76];							inform_R[78][3] = r_cell_wire[77];							inform_R[75][3] = r_cell_wire[78];							inform_R[79][3] = r_cell_wire[79];							inform_R[80][3] = r_cell_wire[80];							inform_R[84][3] = r_cell_wire[81];							inform_R[81][3] = r_cell_wire[82];							inform_R[85][3] = r_cell_wire[83];							inform_R[82][3] = r_cell_wire[84];							inform_R[86][3] = r_cell_wire[85];							inform_R[83][3] = r_cell_wire[86];							inform_R[87][3] = r_cell_wire[87];							inform_R[88][3] = r_cell_wire[88];							inform_R[92][3] = r_cell_wire[89];							inform_R[89][3] = r_cell_wire[90];							inform_R[93][3] = r_cell_wire[91];							inform_R[90][3] = r_cell_wire[92];							inform_R[94][3] = r_cell_wire[93];							inform_R[91][3] = r_cell_wire[94];							inform_R[95][3] = r_cell_wire[95];							inform_R[96][3] = r_cell_wire[96];							inform_R[100][3] = r_cell_wire[97];							inform_R[97][3] = r_cell_wire[98];							inform_R[101][3] = r_cell_wire[99];							inform_R[98][3] = r_cell_wire[100];							inform_R[102][3] = r_cell_wire[101];							inform_R[99][3] = r_cell_wire[102];							inform_R[103][3] = r_cell_wire[103];							inform_R[104][3] = r_cell_wire[104];							inform_R[108][3] = r_cell_wire[105];							inform_R[105][3] = r_cell_wire[106];							inform_R[109][3] = r_cell_wire[107];							inform_R[106][3] = r_cell_wire[108];							inform_R[110][3] = r_cell_wire[109];							inform_R[107][3] = r_cell_wire[110];							inform_R[111][3] = r_cell_wire[111];							inform_R[112][3] = r_cell_wire[112];							inform_R[116][3] = r_cell_wire[113];							inform_R[113][3] = r_cell_wire[114];							inform_R[117][3] = r_cell_wire[115];							inform_R[114][3] = r_cell_wire[116];							inform_R[118][3] = r_cell_wire[117];							inform_R[115][3] = r_cell_wire[118];							inform_R[119][3] = r_cell_wire[119];							inform_R[120][3] = r_cell_wire[120];							inform_R[124][3] = r_cell_wire[121];							inform_R[121][3] = r_cell_wire[122];							inform_R[125][3] = r_cell_wire[123];							inform_R[122][3] = r_cell_wire[124];							inform_R[126][3] = r_cell_wire[125];							inform_R[123][3] = r_cell_wire[126];							inform_R[127][3] = r_cell_wire[127];							inform_R[128][3] = r_cell_wire[128];							inform_R[132][3] = r_cell_wire[129];							inform_R[129][3] = r_cell_wire[130];							inform_R[133][3] = r_cell_wire[131];							inform_R[130][3] = r_cell_wire[132];							inform_R[134][3] = r_cell_wire[133];							inform_R[131][3] = r_cell_wire[134];							inform_R[135][3] = r_cell_wire[135];							inform_R[136][3] = r_cell_wire[136];							inform_R[140][3] = r_cell_wire[137];							inform_R[137][3] = r_cell_wire[138];							inform_R[141][3] = r_cell_wire[139];							inform_R[138][3] = r_cell_wire[140];							inform_R[142][3] = r_cell_wire[141];							inform_R[139][3] = r_cell_wire[142];							inform_R[143][3] = r_cell_wire[143];							inform_R[144][3] = r_cell_wire[144];							inform_R[148][3] = r_cell_wire[145];							inform_R[145][3] = r_cell_wire[146];							inform_R[149][3] = r_cell_wire[147];							inform_R[146][3] = r_cell_wire[148];							inform_R[150][3] = r_cell_wire[149];							inform_R[147][3] = r_cell_wire[150];							inform_R[151][3] = r_cell_wire[151];							inform_R[152][3] = r_cell_wire[152];							inform_R[156][3] = r_cell_wire[153];							inform_R[153][3] = r_cell_wire[154];							inform_R[157][3] = r_cell_wire[155];							inform_R[154][3] = r_cell_wire[156];							inform_R[158][3] = r_cell_wire[157];							inform_R[155][3] = r_cell_wire[158];							inform_R[159][3] = r_cell_wire[159];							inform_R[160][3] = r_cell_wire[160];							inform_R[164][3] = r_cell_wire[161];							inform_R[161][3] = r_cell_wire[162];							inform_R[165][3] = r_cell_wire[163];							inform_R[162][3] = r_cell_wire[164];							inform_R[166][3] = r_cell_wire[165];							inform_R[163][3] = r_cell_wire[166];							inform_R[167][3] = r_cell_wire[167];							inform_R[168][3] = r_cell_wire[168];							inform_R[172][3] = r_cell_wire[169];							inform_R[169][3] = r_cell_wire[170];							inform_R[173][3] = r_cell_wire[171];							inform_R[170][3] = r_cell_wire[172];							inform_R[174][3] = r_cell_wire[173];							inform_R[171][3] = r_cell_wire[174];							inform_R[175][3] = r_cell_wire[175];							inform_R[176][3] = r_cell_wire[176];							inform_R[180][3] = r_cell_wire[177];							inform_R[177][3] = r_cell_wire[178];							inform_R[181][3] = r_cell_wire[179];							inform_R[178][3] = r_cell_wire[180];							inform_R[182][3] = r_cell_wire[181];							inform_R[179][3] = r_cell_wire[182];							inform_R[183][3] = r_cell_wire[183];							inform_R[184][3] = r_cell_wire[184];							inform_R[188][3] = r_cell_wire[185];							inform_R[185][3] = r_cell_wire[186];							inform_R[189][3] = r_cell_wire[187];							inform_R[186][3] = r_cell_wire[188];							inform_R[190][3] = r_cell_wire[189];							inform_R[187][3] = r_cell_wire[190];							inform_R[191][3] = r_cell_wire[191];							inform_R[192][3] = r_cell_wire[192];							inform_R[196][3] = r_cell_wire[193];							inform_R[193][3] = r_cell_wire[194];							inform_R[197][3] = r_cell_wire[195];							inform_R[194][3] = r_cell_wire[196];							inform_R[198][3] = r_cell_wire[197];							inform_R[195][3] = r_cell_wire[198];							inform_R[199][3] = r_cell_wire[199];							inform_R[200][3] = r_cell_wire[200];							inform_R[204][3] = r_cell_wire[201];							inform_R[201][3] = r_cell_wire[202];							inform_R[205][3] = r_cell_wire[203];							inform_R[202][3] = r_cell_wire[204];							inform_R[206][3] = r_cell_wire[205];							inform_R[203][3] = r_cell_wire[206];							inform_R[207][3] = r_cell_wire[207];							inform_R[208][3] = r_cell_wire[208];							inform_R[212][3] = r_cell_wire[209];							inform_R[209][3] = r_cell_wire[210];							inform_R[213][3] = r_cell_wire[211];							inform_R[210][3] = r_cell_wire[212];							inform_R[214][3] = r_cell_wire[213];							inform_R[211][3] = r_cell_wire[214];							inform_R[215][3] = r_cell_wire[215];							inform_R[216][3] = r_cell_wire[216];							inform_R[220][3] = r_cell_wire[217];							inform_R[217][3] = r_cell_wire[218];							inform_R[221][3] = r_cell_wire[219];							inform_R[218][3] = r_cell_wire[220];							inform_R[222][3] = r_cell_wire[221];							inform_R[219][3] = r_cell_wire[222];							inform_R[223][3] = r_cell_wire[223];							inform_R[224][3] = r_cell_wire[224];							inform_R[228][3] = r_cell_wire[225];							inform_R[225][3] = r_cell_wire[226];							inform_R[229][3] = r_cell_wire[227];							inform_R[226][3] = r_cell_wire[228];							inform_R[230][3] = r_cell_wire[229];							inform_R[227][3] = r_cell_wire[230];							inform_R[231][3] = r_cell_wire[231];							inform_R[232][3] = r_cell_wire[232];							inform_R[236][3] = r_cell_wire[233];							inform_R[233][3] = r_cell_wire[234];							inform_R[237][3] = r_cell_wire[235];							inform_R[234][3] = r_cell_wire[236];							inform_R[238][3] = r_cell_wire[237];							inform_R[235][3] = r_cell_wire[238];							inform_R[239][3] = r_cell_wire[239];							inform_R[240][3] = r_cell_wire[240];							inform_R[244][3] = r_cell_wire[241];							inform_R[241][3] = r_cell_wire[242];							inform_R[245][3] = r_cell_wire[243];							inform_R[242][3] = r_cell_wire[244];							inform_R[246][3] = r_cell_wire[245];							inform_R[243][3] = r_cell_wire[246];							inform_R[247][3] = r_cell_wire[247];							inform_R[248][3] = r_cell_wire[248];							inform_R[252][3] = r_cell_wire[249];							inform_R[249][3] = r_cell_wire[250];							inform_R[253][3] = r_cell_wire[251];							inform_R[250][3] = r_cell_wire[252];							inform_R[254][3] = r_cell_wire[253];							inform_R[251][3] = r_cell_wire[254];							inform_R[255][3] = r_cell_wire[255];							inform_R[256][3] = r_cell_wire[256];							inform_R[260][3] = r_cell_wire[257];							inform_R[257][3] = r_cell_wire[258];							inform_R[261][3] = r_cell_wire[259];							inform_R[258][3] = r_cell_wire[260];							inform_R[262][3] = r_cell_wire[261];							inform_R[259][3] = r_cell_wire[262];							inform_R[263][3] = r_cell_wire[263];							inform_R[264][3] = r_cell_wire[264];							inform_R[268][3] = r_cell_wire[265];							inform_R[265][3] = r_cell_wire[266];							inform_R[269][3] = r_cell_wire[267];							inform_R[266][3] = r_cell_wire[268];							inform_R[270][3] = r_cell_wire[269];							inform_R[267][3] = r_cell_wire[270];							inform_R[271][3] = r_cell_wire[271];							inform_R[272][3] = r_cell_wire[272];							inform_R[276][3] = r_cell_wire[273];							inform_R[273][3] = r_cell_wire[274];							inform_R[277][3] = r_cell_wire[275];							inform_R[274][3] = r_cell_wire[276];							inform_R[278][3] = r_cell_wire[277];							inform_R[275][3] = r_cell_wire[278];							inform_R[279][3] = r_cell_wire[279];							inform_R[280][3] = r_cell_wire[280];							inform_R[284][3] = r_cell_wire[281];							inform_R[281][3] = r_cell_wire[282];							inform_R[285][3] = r_cell_wire[283];							inform_R[282][3] = r_cell_wire[284];							inform_R[286][3] = r_cell_wire[285];							inform_R[283][3] = r_cell_wire[286];							inform_R[287][3] = r_cell_wire[287];							inform_R[288][3] = r_cell_wire[288];							inform_R[292][3] = r_cell_wire[289];							inform_R[289][3] = r_cell_wire[290];							inform_R[293][3] = r_cell_wire[291];							inform_R[290][3] = r_cell_wire[292];							inform_R[294][3] = r_cell_wire[293];							inform_R[291][3] = r_cell_wire[294];							inform_R[295][3] = r_cell_wire[295];							inform_R[296][3] = r_cell_wire[296];							inform_R[300][3] = r_cell_wire[297];							inform_R[297][3] = r_cell_wire[298];							inform_R[301][3] = r_cell_wire[299];							inform_R[298][3] = r_cell_wire[300];							inform_R[302][3] = r_cell_wire[301];							inform_R[299][3] = r_cell_wire[302];							inform_R[303][3] = r_cell_wire[303];							inform_R[304][3] = r_cell_wire[304];							inform_R[308][3] = r_cell_wire[305];							inform_R[305][3] = r_cell_wire[306];							inform_R[309][3] = r_cell_wire[307];							inform_R[306][3] = r_cell_wire[308];							inform_R[310][3] = r_cell_wire[309];							inform_R[307][3] = r_cell_wire[310];							inform_R[311][3] = r_cell_wire[311];							inform_R[312][3] = r_cell_wire[312];							inform_R[316][3] = r_cell_wire[313];							inform_R[313][3] = r_cell_wire[314];							inform_R[317][3] = r_cell_wire[315];							inform_R[314][3] = r_cell_wire[316];							inform_R[318][3] = r_cell_wire[317];							inform_R[315][3] = r_cell_wire[318];							inform_R[319][3] = r_cell_wire[319];							inform_R[320][3] = r_cell_wire[320];							inform_R[324][3] = r_cell_wire[321];							inform_R[321][3] = r_cell_wire[322];							inform_R[325][3] = r_cell_wire[323];							inform_R[322][3] = r_cell_wire[324];							inform_R[326][3] = r_cell_wire[325];							inform_R[323][3] = r_cell_wire[326];							inform_R[327][3] = r_cell_wire[327];							inform_R[328][3] = r_cell_wire[328];							inform_R[332][3] = r_cell_wire[329];							inform_R[329][3] = r_cell_wire[330];							inform_R[333][3] = r_cell_wire[331];							inform_R[330][3] = r_cell_wire[332];							inform_R[334][3] = r_cell_wire[333];							inform_R[331][3] = r_cell_wire[334];							inform_R[335][3] = r_cell_wire[335];							inform_R[336][3] = r_cell_wire[336];							inform_R[340][3] = r_cell_wire[337];							inform_R[337][3] = r_cell_wire[338];							inform_R[341][3] = r_cell_wire[339];							inform_R[338][3] = r_cell_wire[340];							inform_R[342][3] = r_cell_wire[341];							inform_R[339][3] = r_cell_wire[342];							inform_R[343][3] = r_cell_wire[343];							inform_R[344][3] = r_cell_wire[344];							inform_R[348][3] = r_cell_wire[345];							inform_R[345][3] = r_cell_wire[346];							inform_R[349][3] = r_cell_wire[347];							inform_R[346][3] = r_cell_wire[348];							inform_R[350][3] = r_cell_wire[349];							inform_R[347][3] = r_cell_wire[350];							inform_R[351][3] = r_cell_wire[351];							inform_R[352][3] = r_cell_wire[352];							inform_R[356][3] = r_cell_wire[353];							inform_R[353][3] = r_cell_wire[354];							inform_R[357][3] = r_cell_wire[355];							inform_R[354][3] = r_cell_wire[356];							inform_R[358][3] = r_cell_wire[357];							inform_R[355][3] = r_cell_wire[358];							inform_R[359][3] = r_cell_wire[359];							inform_R[360][3] = r_cell_wire[360];							inform_R[364][3] = r_cell_wire[361];							inform_R[361][3] = r_cell_wire[362];							inform_R[365][3] = r_cell_wire[363];							inform_R[362][3] = r_cell_wire[364];							inform_R[366][3] = r_cell_wire[365];							inform_R[363][3] = r_cell_wire[366];							inform_R[367][3] = r_cell_wire[367];							inform_R[368][3] = r_cell_wire[368];							inform_R[372][3] = r_cell_wire[369];							inform_R[369][3] = r_cell_wire[370];							inform_R[373][3] = r_cell_wire[371];							inform_R[370][3] = r_cell_wire[372];							inform_R[374][3] = r_cell_wire[373];							inform_R[371][3] = r_cell_wire[374];							inform_R[375][3] = r_cell_wire[375];							inform_R[376][3] = r_cell_wire[376];							inform_R[380][3] = r_cell_wire[377];							inform_R[377][3] = r_cell_wire[378];							inform_R[381][3] = r_cell_wire[379];							inform_R[378][3] = r_cell_wire[380];							inform_R[382][3] = r_cell_wire[381];							inform_R[379][3] = r_cell_wire[382];							inform_R[383][3] = r_cell_wire[383];							inform_R[384][3] = r_cell_wire[384];							inform_R[388][3] = r_cell_wire[385];							inform_R[385][3] = r_cell_wire[386];							inform_R[389][3] = r_cell_wire[387];							inform_R[386][3] = r_cell_wire[388];							inform_R[390][3] = r_cell_wire[389];							inform_R[387][3] = r_cell_wire[390];							inform_R[391][3] = r_cell_wire[391];							inform_R[392][3] = r_cell_wire[392];							inform_R[396][3] = r_cell_wire[393];							inform_R[393][3] = r_cell_wire[394];							inform_R[397][3] = r_cell_wire[395];							inform_R[394][3] = r_cell_wire[396];							inform_R[398][3] = r_cell_wire[397];							inform_R[395][3] = r_cell_wire[398];							inform_R[399][3] = r_cell_wire[399];							inform_R[400][3] = r_cell_wire[400];							inform_R[404][3] = r_cell_wire[401];							inform_R[401][3] = r_cell_wire[402];							inform_R[405][3] = r_cell_wire[403];							inform_R[402][3] = r_cell_wire[404];							inform_R[406][3] = r_cell_wire[405];							inform_R[403][3] = r_cell_wire[406];							inform_R[407][3] = r_cell_wire[407];							inform_R[408][3] = r_cell_wire[408];							inform_R[412][3] = r_cell_wire[409];							inform_R[409][3] = r_cell_wire[410];							inform_R[413][3] = r_cell_wire[411];							inform_R[410][3] = r_cell_wire[412];							inform_R[414][3] = r_cell_wire[413];							inform_R[411][3] = r_cell_wire[414];							inform_R[415][3] = r_cell_wire[415];							inform_R[416][3] = r_cell_wire[416];							inform_R[420][3] = r_cell_wire[417];							inform_R[417][3] = r_cell_wire[418];							inform_R[421][3] = r_cell_wire[419];							inform_R[418][3] = r_cell_wire[420];							inform_R[422][3] = r_cell_wire[421];							inform_R[419][3] = r_cell_wire[422];							inform_R[423][3] = r_cell_wire[423];							inform_R[424][3] = r_cell_wire[424];							inform_R[428][3] = r_cell_wire[425];							inform_R[425][3] = r_cell_wire[426];							inform_R[429][3] = r_cell_wire[427];							inform_R[426][3] = r_cell_wire[428];							inform_R[430][3] = r_cell_wire[429];							inform_R[427][3] = r_cell_wire[430];							inform_R[431][3] = r_cell_wire[431];							inform_R[432][3] = r_cell_wire[432];							inform_R[436][3] = r_cell_wire[433];							inform_R[433][3] = r_cell_wire[434];							inform_R[437][3] = r_cell_wire[435];							inform_R[434][3] = r_cell_wire[436];							inform_R[438][3] = r_cell_wire[437];							inform_R[435][3] = r_cell_wire[438];							inform_R[439][3] = r_cell_wire[439];							inform_R[440][3] = r_cell_wire[440];							inform_R[444][3] = r_cell_wire[441];							inform_R[441][3] = r_cell_wire[442];							inform_R[445][3] = r_cell_wire[443];							inform_R[442][3] = r_cell_wire[444];							inform_R[446][3] = r_cell_wire[445];							inform_R[443][3] = r_cell_wire[446];							inform_R[447][3] = r_cell_wire[447];							inform_R[448][3] = r_cell_wire[448];							inform_R[452][3] = r_cell_wire[449];							inform_R[449][3] = r_cell_wire[450];							inform_R[453][3] = r_cell_wire[451];							inform_R[450][3] = r_cell_wire[452];							inform_R[454][3] = r_cell_wire[453];							inform_R[451][3] = r_cell_wire[454];							inform_R[455][3] = r_cell_wire[455];							inform_R[456][3] = r_cell_wire[456];							inform_R[460][3] = r_cell_wire[457];							inform_R[457][3] = r_cell_wire[458];							inform_R[461][3] = r_cell_wire[459];							inform_R[458][3] = r_cell_wire[460];							inform_R[462][3] = r_cell_wire[461];							inform_R[459][3] = r_cell_wire[462];							inform_R[463][3] = r_cell_wire[463];							inform_R[464][3] = r_cell_wire[464];							inform_R[468][3] = r_cell_wire[465];							inform_R[465][3] = r_cell_wire[466];							inform_R[469][3] = r_cell_wire[467];							inform_R[466][3] = r_cell_wire[468];							inform_R[470][3] = r_cell_wire[469];							inform_R[467][3] = r_cell_wire[470];							inform_R[471][3] = r_cell_wire[471];							inform_R[472][3] = r_cell_wire[472];							inform_R[476][3] = r_cell_wire[473];							inform_R[473][3] = r_cell_wire[474];							inform_R[477][3] = r_cell_wire[475];							inform_R[474][3] = r_cell_wire[476];							inform_R[478][3] = r_cell_wire[477];							inform_R[475][3] = r_cell_wire[478];							inform_R[479][3] = r_cell_wire[479];							inform_R[480][3] = r_cell_wire[480];							inform_R[484][3] = r_cell_wire[481];							inform_R[481][3] = r_cell_wire[482];							inform_R[485][3] = r_cell_wire[483];							inform_R[482][3] = r_cell_wire[484];							inform_R[486][3] = r_cell_wire[485];							inform_R[483][3] = r_cell_wire[486];							inform_R[487][3] = r_cell_wire[487];							inform_R[488][3] = r_cell_wire[488];							inform_R[492][3] = r_cell_wire[489];							inform_R[489][3] = r_cell_wire[490];							inform_R[493][3] = r_cell_wire[491];							inform_R[490][3] = r_cell_wire[492];							inform_R[494][3] = r_cell_wire[493];							inform_R[491][3] = r_cell_wire[494];							inform_R[495][3] = r_cell_wire[495];							inform_R[496][3] = r_cell_wire[496];							inform_R[500][3] = r_cell_wire[497];							inform_R[497][3] = r_cell_wire[498];							inform_R[501][3] = r_cell_wire[499];							inform_R[498][3] = r_cell_wire[500];							inform_R[502][3] = r_cell_wire[501];							inform_R[499][3] = r_cell_wire[502];							inform_R[503][3] = r_cell_wire[503];							inform_R[504][3] = r_cell_wire[504];							inform_R[508][3] = r_cell_wire[505];							inform_R[505][3] = r_cell_wire[506];							inform_R[509][3] = r_cell_wire[507];							inform_R[506][3] = r_cell_wire[508];							inform_R[510][3] = r_cell_wire[509];							inform_R[507][3] = r_cell_wire[510];							inform_R[511][3] = r_cell_wire[511];							inform_R[512][3] = r_cell_wire[512];							inform_R[516][3] = r_cell_wire[513];							inform_R[513][3] = r_cell_wire[514];							inform_R[517][3] = r_cell_wire[515];							inform_R[514][3] = r_cell_wire[516];							inform_R[518][3] = r_cell_wire[517];							inform_R[515][3] = r_cell_wire[518];							inform_R[519][3] = r_cell_wire[519];							inform_R[520][3] = r_cell_wire[520];							inform_R[524][3] = r_cell_wire[521];							inform_R[521][3] = r_cell_wire[522];							inform_R[525][3] = r_cell_wire[523];							inform_R[522][3] = r_cell_wire[524];							inform_R[526][3] = r_cell_wire[525];							inform_R[523][3] = r_cell_wire[526];							inform_R[527][3] = r_cell_wire[527];							inform_R[528][3] = r_cell_wire[528];							inform_R[532][3] = r_cell_wire[529];							inform_R[529][3] = r_cell_wire[530];							inform_R[533][3] = r_cell_wire[531];							inform_R[530][3] = r_cell_wire[532];							inform_R[534][3] = r_cell_wire[533];							inform_R[531][3] = r_cell_wire[534];							inform_R[535][3] = r_cell_wire[535];							inform_R[536][3] = r_cell_wire[536];							inform_R[540][3] = r_cell_wire[537];							inform_R[537][3] = r_cell_wire[538];							inform_R[541][3] = r_cell_wire[539];							inform_R[538][3] = r_cell_wire[540];							inform_R[542][3] = r_cell_wire[541];							inform_R[539][3] = r_cell_wire[542];							inform_R[543][3] = r_cell_wire[543];							inform_R[544][3] = r_cell_wire[544];							inform_R[548][3] = r_cell_wire[545];							inform_R[545][3] = r_cell_wire[546];							inform_R[549][3] = r_cell_wire[547];							inform_R[546][3] = r_cell_wire[548];							inform_R[550][3] = r_cell_wire[549];							inform_R[547][3] = r_cell_wire[550];							inform_R[551][3] = r_cell_wire[551];							inform_R[552][3] = r_cell_wire[552];							inform_R[556][3] = r_cell_wire[553];							inform_R[553][3] = r_cell_wire[554];							inform_R[557][3] = r_cell_wire[555];							inform_R[554][3] = r_cell_wire[556];							inform_R[558][3] = r_cell_wire[557];							inform_R[555][3] = r_cell_wire[558];							inform_R[559][3] = r_cell_wire[559];							inform_R[560][3] = r_cell_wire[560];							inform_R[564][3] = r_cell_wire[561];							inform_R[561][3] = r_cell_wire[562];							inform_R[565][3] = r_cell_wire[563];							inform_R[562][3] = r_cell_wire[564];							inform_R[566][3] = r_cell_wire[565];							inform_R[563][3] = r_cell_wire[566];							inform_R[567][3] = r_cell_wire[567];							inform_R[568][3] = r_cell_wire[568];							inform_R[572][3] = r_cell_wire[569];							inform_R[569][3] = r_cell_wire[570];							inform_R[573][3] = r_cell_wire[571];							inform_R[570][3] = r_cell_wire[572];							inform_R[574][3] = r_cell_wire[573];							inform_R[571][3] = r_cell_wire[574];							inform_R[575][3] = r_cell_wire[575];							inform_R[576][3] = r_cell_wire[576];							inform_R[580][3] = r_cell_wire[577];							inform_R[577][3] = r_cell_wire[578];							inform_R[581][3] = r_cell_wire[579];							inform_R[578][3] = r_cell_wire[580];							inform_R[582][3] = r_cell_wire[581];							inform_R[579][3] = r_cell_wire[582];							inform_R[583][3] = r_cell_wire[583];							inform_R[584][3] = r_cell_wire[584];							inform_R[588][3] = r_cell_wire[585];							inform_R[585][3] = r_cell_wire[586];							inform_R[589][3] = r_cell_wire[587];							inform_R[586][3] = r_cell_wire[588];							inform_R[590][3] = r_cell_wire[589];							inform_R[587][3] = r_cell_wire[590];							inform_R[591][3] = r_cell_wire[591];							inform_R[592][3] = r_cell_wire[592];							inform_R[596][3] = r_cell_wire[593];							inform_R[593][3] = r_cell_wire[594];							inform_R[597][3] = r_cell_wire[595];							inform_R[594][3] = r_cell_wire[596];							inform_R[598][3] = r_cell_wire[597];							inform_R[595][3] = r_cell_wire[598];							inform_R[599][3] = r_cell_wire[599];							inform_R[600][3] = r_cell_wire[600];							inform_R[604][3] = r_cell_wire[601];							inform_R[601][3] = r_cell_wire[602];							inform_R[605][3] = r_cell_wire[603];							inform_R[602][3] = r_cell_wire[604];							inform_R[606][3] = r_cell_wire[605];							inform_R[603][3] = r_cell_wire[606];							inform_R[607][3] = r_cell_wire[607];							inform_R[608][3] = r_cell_wire[608];							inform_R[612][3] = r_cell_wire[609];							inform_R[609][3] = r_cell_wire[610];							inform_R[613][3] = r_cell_wire[611];							inform_R[610][3] = r_cell_wire[612];							inform_R[614][3] = r_cell_wire[613];							inform_R[611][3] = r_cell_wire[614];							inform_R[615][3] = r_cell_wire[615];							inform_R[616][3] = r_cell_wire[616];							inform_R[620][3] = r_cell_wire[617];							inform_R[617][3] = r_cell_wire[618];							inform_R[621][3] = r_cell_wire[619];							inform_R[618][3] = r_cell_wire[620];							inform_R[622][3] = r_cell_wire[621];							inform_R[619][3] = r_cell_wire[622];							inform_R[623][3] = r_cell_wire[623];							inform_R[624][3] = r_cell_wire[624];							inform_R[628][3] = r_cell_wire[625];							inform_R[625][3] = r_cell_wire[626];							inform_R[629][3] = r_cell_wire[627];							inform_R[626][3] = r_cell_wire[628];							inform_R[630][3] = r_cell_wire[629];							inform_R[627][3] = r_cell_wire[630];							inform_R[631][3] = r_cell_wire[631];							inform_R[632][3] = r_cell_wire[632];							inform_R[636][3] = r_cell_wire[633];							inform_R[633][3] = r_cell_wire[634];							inform_R[637][3] = r_cell_wire[635];							inform_R[634][3] = r_cell_wire[636];							inform_R[638][3] = r_cell_wire[637];							inform_R[635][3] = r_cell_wire[638];							inform_R[639][3] = r_cell_wire[639];							inform_R[640][3] = r_cell_wire[640];							inform_R[644][3] = r_cell_wire[641];							inform_R[641][3] = r_cell_wire[642];							inform_R[645][3] = r_cell_wire[643];							inform_R[642][3] = r_cell_wire[644];							inform_R[646][3] = r_cell_wire[645];							inform_R[643][3] = r_cell_wire[646];							inform_R[647][3] = r_cell_wire[647];							inform_R[648][3] = r_cell_wire[648];							inform_R[652][3] = r_cell_wire[649];							inform_R[649][3] = r_cell_wire[650];							inform_R[653][3] = r_cell_wire[651];							inform_R[650][3] = r_cell_wire[652];							inform_R[654][3] = r_cell_wire[653];							inform_R[651][3] = r_cell_wire[654];							inform_R[655][3] = r_cell_wire[655];							inform_R[656][3] = r_cell_wire[656];							inform_R[660][3] = r_cell_wire[657];							inform_R[657][3] = r_cell_wire[658];							inform_R[661][3] = r_cell_wire[659];							inform_R[658][3] = r_cell_wire[660];							inform_R[662][3] = r_cell_wire[661];							inform_R[659][3] = r_cell_wire[662];							inform_R[663][3] = r_cell_wire[663];							inform_R[664][3] = r_cell_wire[664];							inform_R[668][3] = r_cell_wire[665];							inform_R[665][3] = r_cell_wire[666];							inform_R[669][3] = r_cell_wire[667];							inform_R[666][3] = r_cell_wire[668];							inform_R[670][3] = r_cell_wire[669];							inform_R[667][3] = r_cell_wire[670];							inform_R[671][3] = r_cell_wire[671];							inform_R[672][3] = r_cell_wire[672];							inform_R[676][3] = r_cell_wire[673];							inform_R[673][3] = r_cell_wire[674];							inform_R[677][3] = r_cell_wire[675];							inform_R[674][3] = r_cell_wire[676];							inform_R[678][3] = r_cell_wire[677];							inform_R[675][3] = r_cell_wire[678];							inform_R[679][3] = r_cell_wire[679];							inform_R[680][3] = r_cell_wire[680];							inform_R[684][3] = r_cell_wire[681];							inform_R[681][3] = r_cell_wire[682];							inform_R[685][3] = r_cell_wire[683];							inform_R[682][3] = r_cell_wire[684];							inform_R[686][3] = r_cell_wire[685];							inform_R[683][3] = r_cell_wire[686];							inform_R[687][3] = r_cell_wire[687];							inform_R[688][3] = r_cell_wire[688];							inform_R[692][3] = r_cell_wire[689];							inform_R[689][3] = r_cell_wire[690];							inform_R[693][3] = r_cell_wire[691];							inform_R[690][3] = r_cell_wire[692];							inform_R[694][3] = r_cell_wire[693];							inform_R[691][3] = r_cell_wire[694];							inform_R[695][3] = r_cell_wire[695];							inform_R[696][3] = r_cell_wire[696];							inform_R[700][3] = r_cell_wire[697];							inform_R[697][3] = r_cell_wire[698];							inform_R[701][3] = r_cell_wire[699];							inform_R[698][3] = r_cell_wire[700];							inform_R[702][3] = r_cell_wire[701];							inform_R[699][3] = r_cell_wire[702];							inform_R[703][3] = r_cell_wire[703];							inform_R[704][3] = r_cell_wire[704];							inform_R[708][3] = r_cell_wire[705];							inform_R[705][3] = r_cell_wire[706];							inform_R[709][3] = r_cell_wire[707];							inform_R[706][3] = r_cell_wire[708];							inform_R[710][3] = r_cell_wire[709];							inform_R[707][3] = r_cell_wire[710];							inform_R[711][3] = r_cell_wire[711];							inform_R[712][3] = r_cell_wire[712];							inform_R[716][3] = r_cell_wire[713];							inform_R[713][3] = r_cell_wire[714];							inform_R[717][3] = r_cell_wire[715];							inform_R[714][3] = r_cell_wire[716];							inform_R[718][3] = r_cell_wire[717];							inform_R[715][3] = r_cell_wire[718];							inform_R[719][3] = r_cell_wire[719];							inform_R[720][3] = r_cell_wire[720];							inform_R[724][3] = r_cell_wire[721];							inform_R[721][3] = r_cell_wire[722];							inform_R[725][3] = r_cell_wire[723];							inform_R[722][3] = r_cell_wire[724];							inform_R[726][3] = r_cell_wire[725];							inform_R[723][3] = r_cell_wire[726];							inform_R[727][3] = r_cell_wire[727];							inform_R[728][3] = r_cell_wire[728];							inform_R[732][3] = r_cell_wire[729];							inform_R[729][3] = r_cell_wire[730];							inform_R[733][3] = r_cell_wire[731];							inform_R[730][3] = r_cell_wire[732];							inform_R[734][3] = r_cell_wire[733];							inform_R[731][3] = r_cell_wire[734];							inform_R[735][3] = r_cell_wire[735];							inform_R[736][3] = r_cell_wire[736];							inform_R[740][3] = r_cell_wire[737];							inform_R[737][3] = r_cell_wire[738];							inform_R[741][3] = r_cell_wire[739];							inform_R[738][3] = r_cell_wire[740];							inform_R[742][3] = r_cell_wire[741];							inform_R[739][3] = r_cell_wire[742];							inform_R[743][3] = r_cell_wire[743];							inform_R[744][3] = r_cell_wire[744];							inform_R[748][3] = r_cell_wire[745];							inform_R[745][3] = r_cell_wire[746];							inform_R[749][3] = r_cell_wire[747];							inform_R[746][3] = r_cell_wire[748];							inform_R[750][3] = r_cell_wire[749];							inform_R[747][3] = r_cell_wire[750];							inform_R[751][3] = r_cell_wire[751];							inform_R[752][3] = r_cell_wire[752];							inform_R[756][3] = r_cell_wire[753];							inform_R[753][3] = r_cell_wire[754];							inform_R[757][3] = r_cell_wire[755];							inform_R[754][3] = r_cell_wire[756];							inform_R[758][3] = r_cell_wire[757];							inform_R[755][3] = r_cell_wire[758];							inform_R[759][3] = r_cell_wire[759];							inform_R[760][3] = r_cell_wire[760];							inform_R[764][3] = r_cell_wire[761];							inform_R[761][3] = r_cell_wire[762];							inform_R[765][3] = r_cell_wire[763];							inform_R[762][3] = r_cell_wire[764];							inform_R[766][3] = r_cell_wire[765];							inform_R[763][3] = r_cell_wire[766];							inform_R[767][3] = r_cell_wire[767];							inform_R[768][3] = r_cell_wire[768];							inform_R[772][3] = r_cell_wire[769];							inform_R[769][3] = r_cell_wire[770];							inform_R[773][3] = r_cell_wire[771];							inform_R[770][3] = r_cell_wire[772];							inform_R[774][3] = r_cell_wire[773];							inform_R[771][3] = r_cell_wire[774];							inform_R[775][3] = r_cell_wire[775];							inform_R[776][3] = r_cell_wire[776];							inform_R[780][3] = r_cell_wire[777];							inform_R[777][3] = r_cell_wire[778];							inform_R[781][3] = r_cell_wire[779];							inform_R[778][3] = r_cell_wire[780];							inform_R[782][3] = r_cell_wire[781];							inform_R[779][3] = r_cell_wire[782];							inform_R[783][3] = r_cell_wire[783];							inform_R[784][3] = r_cell_wire[784];							inform_R[788][3] = r_cell_wire[785];							inform_R[785][3] = r_cell_wire[786];							inform_R[789][3] = r_cell_wire[787];							inform_R[786][3] = r_cell_wire[788];							inform_R[790][3] = r_cell_wire[789];							inform_R[787][3] = r_cell_wire[790];							inform_R[791][3] = r_cell_wire[791];							inform_R[792][3] = r_cell_wire[792];							inform_R[796][3] = r_cell_wire[793];							inform_R[793][3] = r_cell_wire[794];							inform_R[797][3] = r_cell_wire[795];							inform_R[794][3] = r_cell_wire[796];							inform_R[798][3] = r_cell_wire[797];							inform_R[795][3] = r_cell_wire[798];							inform_R[799][3] = r_cell_wire[799];							inform_R[800][3] = r_cell_wire[800];							inform_R[804][3] = r_cell_wire[801];							inform_R[801][3] = r_cell_wire[802];							inform_R[805][3] = r_cell_wire[803];							inform_R[802][3] = r_cell_wire[804];							inform_R[806][3] = r_cell_wire[805];							inform_R[803][3] = r_cell_wire[806];							inform_R[807][3] = r_cell_wire[807];							inform_R[808][3] = r_cell_wire[808];							inform_R[812][3] = r_cell_wire[809];							inform_R[809][3] = r_cell_wire[810];							inform_R[813][3] = r_cell_wire[811];							inform_R[810][3] = r_cell_wire[812];							inform_R[814][3] = r_cell_wire[813];							inform_R[811][3] = r_cell_wire[814];							inform_R[815][3] = r_cell_wire[815];							inform_R[816][3] = r_cell_wire[816];							inform_R[820][3] = r_cell_wire[817];							inform_R[817][3] = r_cell_wire[818];							inform_R[821][3] = r_cell_wire[819];							inform_R[818][3] = r_cell_wire[820];							inform_R[822][3] = r_cell_wire[821];							inform_R[819][3] = r_cell_wire[822];							inform_R[823][3] = r_cell_wire[823];							inform_R[824][3] = r_cell_wire[824];							inform_R[828][3] = r_cell_wire[825];							inform_R[825][3] = r_cell_wire[826];							inform_R[829][3] = r_cell_wire[827];							inform_R[826][3] = r_cell_wire[828];							inform_R[830][3] = r_cell_wire[829];							inform_R[827][3] = r_cell_wire[830];							inform_R[831][3] = r_cell_wire[831];							inform_R[832][3] = r_cell_wire[832];							inform_R[836][3] = r_cell_wire[833];							inform_R[833][3] = r_cell_wire[834];							inform_R[837][3] = r_cell_wire[835];							inform_R[834][3] = r_cell_wire[836];							inform_R[838][3] = r_cell_wire[837];							inform_R[835][3] = r_cell_wire[838];							inform_R[839][3] = r_cell_wire[839];							inform_R[840][3] = r_cell_wire[840];							inform_R[844][3] = r_cell_wire[841];							inform_R[841][3] = r_cell_wire[842];							inform_R[845][3] = r_cell_wire[843];							inform_R[842][3] = r_cell_wire[844];							inform_R[846][3] = r_cell_wire[845];							inform_R[843][3] = r_cell_wire[846];							inform_R[847][3] = r_cell_wire[847];							inform_R[848][3] = r_cell_wire[848];							inform_R[852][3] = r_cell_wire[849];							inform_R[849][3] = r_cell_wire[850];							inform_R[853][3] = r_cell_wire[851];							inform_R[850][3] = r_cell_wire[852];							inform_R[854][3] = r_cell_wire[853];							inform_R[851][3] = r_cell_wire[854];							inform_R[855][3] = r_cell_wire[855];							inform_R[856][3] = r_cell_wire[856];							inform_R[860][3] = r_cell_wire[857];							inform_R[857][3] = r_cell_wire[858];							inform_R[861][3] = r_cell_wire[859];							inform_R[858][3] = r_cell_wire[860];							inform_R[862][3] = r_cell_wire[861];							inform_R[859][3] = r_cell_wire[862];							inform_R[863][3] = r_cell_wire[863];							inform_R[864][3] = r_cell_wire[864];							inform_R[868][3] = r_cell_wire[865];							inform_R[865][3] = r_cell_wire[866];							inform_R[869][3] = r_cell_wire[867];							inform_R[866][3] = r_cell_wire[868];							inform_R[870][3] = r_cell_wire[869];							inform_R[867][3] = r_cell_wire[870];							inform_R[871][3] = r_cell_wire[871];							inform_R[872][3] = r_cell_wire[872];							inform_R[876][3] = r_cell_wire[873];							inform_R[873][3] = r_cell_wire[874];							inform_R[877][3] = r_cell_wire[875];							inform_R[874][3] = r_cell_wire[876];							inform_R[878][3] = r_cell_wire[877];							inform_R[875][3] = r_cell_wire[878];							inform_R[879][3] = r_cell_wire[879];							inform_R[880][3] = r_cell_wire[880];							inform_R[884][3] = r_cell_wire[881];							inform_R[881][3] = r_cell_wire[882];							inform_R[885][3] = r_cell_wire[883];							inform_R[882][3] = r_cell_wire[884];							inform_R[886][3] = r_cell_wire[885];							inform_R[883][3] = r_cell_wire[886];							inform_R[887][3] = r_cell_wire[887];							inform_R[888][3] = r_cell_wire[888];							inform_R[892][3] = r_cell_wire[889];							inform_R[889][3] = r_cell_wire[890];							inform_R[893][3] = r_cell_wire[891];							inform_R[890][3] = r_cell_wire[892];							inform_R[894][3] = r_cell_wire[893];							inform_R[891][3] = r_cell_wire[894];							inform_R[895][3] = r_cell_wire[895];							inform_R[896][3] = r_cell_wire[896];							inform_R[900][3] = r_cell_wire[897];							inform_R[897][3] = r_cell_wire[898];							inform_R[901][3] = r_cell_wire[899];							inform_R[898][3] = r_cell_wire[900];							inform_R[902][3] = r_cell_wire[901];							inform_R[899][3] = r_cell_wire[902];							inform_R[903][3] = r_cell_wire[903];							inform_R[904][3] = r_cell_wire[904];							inform_R[908][3] = r_cell_wire[905];							inform_R[905][3] = r_cell_wire[906];							inform_R[909][3] = r_cell_wire[907];							inform_R[906][3] = r_cell_wire[908];							inform_R[910][3] = r_cell_wire[909];							inform_R[907][3] = r_cell_wire[910];							inform_R[911][3] = r_cell_wire[911];							inform_R[912][3] = r_cell_wire[912];							inform_R[916][3] = r_cell_wire[913];							inform_R[913][3] = r_cell_wire[914];							inform_R[917][3] = r_cell_wire[915];							inform_R[914][3] = r_cell_wire[916];							inform_R[918][3] = r_cell_wire[917];							inform_R[915][3] = r_cell_wire[918];							inform_R[919][3] = r_cell_wire[919];							inform_R[920][3] = r_cell_wire[920];							inform_R[924][3] = r_cell_wire[921];							inform_R[921][3] = r_cell_wire[922];							inform_R[925][3] = r_cell_wire[923];							inform_R[922][3] = r_cell_wire[924];							inform_R[926][3] = r_cell_wire[925];							inform_R[923][3] = r_cell_wire[926];							inform_R[927][3] = r_cell_wire[927];							inform_R[928][3] = r_cell_wire[928];							inform_R[932][3] = r_cell_wire[929];							inform_R[929][3] = r_cell_wire[930];							inform_R[933][3] = r_cell_wire[931];							inform_R[930][3] = r_cell_wire[932];							inform_R[934][3] = r_cell_wire[933];							inform_R[931][3] = r_cell_wire[934];							inform_R[935][3] = r_cell_wire[935];							inform_R[936][3] = r_cell_wire[936];							inform_R[940][3] = r_cell_wire[937];							inform_R[937][3] = r_cell_wire[938];							inform_R[941][3] = r_cell_wire[939];							inform_R[938][3] = r_cell_wire[940];							inform_R[942][3] = r_cell_wire[941];							inform_R[939][3] = r_cell_wire[942];							inform_R[943][3] = r_cell_wire[943];							inform_R[944][3] = r_cell_wire[944];							inform_R[948][3] = r_cell_wire[945];							inform_R[945][3] = r_cell_wire[946];							inform_R[949][3] = r_cell_wire[947];							inform_R[946][3] = r_cell_wire[948];							inform_R[950][3] = r_cell_wire[949];							inform_R[947][3] = r_cell_wire[950];							inform_R[951][3] = r_cell_wire[951];							inform_R[952][3] = r_cell_wire[952];							inform_R[956][3] = r_cell_wire[953];							inform_R[953][3] = r_cell_wire[954];							inform_R[957][3] = r_cell_wire[955];							inform_R[954][3] = r_cell_wire[956];							inform_R[958][3] = r_cell_wire[957];							inform_R[955][3] = r_cell_wire[958];							inform_R[959][3] = r_cell_wire[959];							inform_R[960][3] = r_cell_wire[960];							inform_R[964][3] = r_cell_wire[961];							inform_R[961][3] = r_cell_wire[962];							inform_R[965][3] = r_cell_wire[963];							inform_R[962][3] = r_cell_wire[964];							inform_R[966][3] = r_cell_wire[965];							inform_R[963][3] = r_cell_wire[966];							inform_R[967][3] = r_cell_wire[967];							inform_R[968][3] = r_cell_wire[968];							inform_R[972][3] = r_cell_wire[969];							inform_R[969][3] = r_cell_wire[970];							inform_R[973][3] = r_cell_wire[971];							inform_R[970][3] = r_cell_wire[972];							inform_R[974][3] = r_cell_wire[973];							inform_R[971][3] = r_cell_wire[974];							inform_R[975][3] = r_cell_wire[975];							inform_R[976][3] = r_cell_wire[976];							inform_R[980][3] = r_cell_wire[977];							inform_R[977][3] = r_cell_wire[978];							inform_R[981][3] = r_cell_wire[979];							inform_R[978][3] = r_cell_wire[980];							inform_R[982][3] = r_cell_wire[981];							inform_R[979][3] = r_cell_wire[982];							inform_R[983][3] = r_cell_wire[983];							inform_R[984][3] = r_cell_wire[984];							inform_R[988][3] = r_cell_wire[985];							inform_R[985][3] = r_cell_wire[986];							inform_R[989][3] = r_cell_wire[987];							inform_R[986][3] = r_cell_wire[988];							inform_R[990][3] = r_cell_wire[989];							inform_R[987][3] = r_cell_wire[990];							inform_R[991][3] = r_cell_wire[991];							inform_R[992][3] = r_cell_wire[992];							inform_R[996][3] = r_cell_wire[993];							inform_R[993][3] = r_cell_wire[994];							inform_R[997][3] = r_cell_wire[995];							inform_R[994][3] = r_cell_wire[996];							inform_R[998][3] = r_cell_wire[997];							inform_R[995][3] = r_cell_wire[998];							inform_R[999][3] = r_cell_wire[999];							inform_R[1000][3] = r_cell_wire[1000];							inform_R[1004][3] = r_cell_wire[1001];							inform_R[1001][3] = r_cell_wire[1002];							inform_R[1005][3] = r_cell_wire[1003];							inform_R[1002][3] = r_cell_wire[1004];							inform_R[1006][3] = r_cell_wire[1005];							inform_R[1003][3] = r_cell_wire[1006];							inform_R[1007][3] = r_cell_wire[1007];							inform_R[1008][3] = r_cell_wire[1008];							inform_R[1012][3] = r_cell_wire[1009];							inform_R[1009][3] = r_cell_wire[1010];							inform_R[1013][3] = r_cell_wire[1011];							inform_R[1010][3] = r_cell_wire[1012];							inform_R[1014][3] = r_cell_wire[1013];							inform_R[1011][3] = r_cell_wire[1014];							inform_R[1015][3] = r_cell_wire[1015];							inform_R[1016][3] = r_cell_wire[1016];							inform_R[1020][3] = r_cell_wire[1017];							inform_R[1017][3] = r_cell_wire[1018];							inform_R[1021][3] = r_cell_wire[1019];							inform_R[1018][3] = r_cell_wire[1020];							inform_R[1022][3] = r_cell_wire[1021];							inform_R[1019][3] = r_cell_wire[1022];							inform_R[1023][3] = r_cell_wire[1023];							inform_L[0][2] = l_cell_wire[0];							inform_L[4][2] = l_cell_wire[1];							inform_L[1][2] = l_cell_wire[2];							inform_L[5][2] = l_cell_wire[3];							inform_L[2][2] = l_cell_wire[4];							inform_L[6][2] = l_cell_wire[5];							inform_L[3][2] = l_cell_wire[6];							inform_L[7][2] = l_cell_wire[7];							inform_L[8][2] = l_cell_wire[8];							inform_L[12][2] = l_cell_wire[9];							inform_L[9][2] = l_cell_wire[10];							inform_L[13][2] = l_cell_wire[11];							inform_L[10][2] = l_cell_wire[12];							inform_L[14][2] = l_cell_wire[13];							inform_L[11][2] = l_cell_wire[14];							inform_L[15][2] = l_cell_wire[15];							inform_L[16][2] = l_cell_wire[16];							inform_L[20][2] = l_cell_wire[17];							inform_L[17][2] = l_cell_wire[18];							inform_L[21][2] = l_cell_wire[19];							inform_L[18][2] = l_cell_wire[20];							inform_L[22][2] = l_cell_wire[21];							inform_L[19][2] = l_cell_wire[22];							inform_L[23][2] = l_cell_wire[23];							inform_L[24][2] = l_cell_wire[24];							inform_L[28][2] = l_cell_wire[25];							inform_L[25][2] = l_cell_wire[26];							inform_L[29][2] = l_cell_wire[27];							inform_L[26][2] = l_cell_wire[28];							inform_L[30][2] = l_cell_wire[29];							inform_L[27][2] = l_cell_wire[30];							inform_L[31][2] = l_cell_wire[31];							inform_L[32][2] = l_cell_wire[32];							inform_L[36][2] = l_cell_wire[33];							inform_L[33][2] = l_cell_wire[34];							inform_L[37][2] = l_cell_wire[35];							inform_L[34][2] = l_cell_wire[36];							inform_L[38][2] = l_cell_wire[37];							inform_L[35][2] = l_cell_wire[38];							inform_L[39][2] = l_cell_wire[39];							inform_L[40][2] = l_cell_wire[40];							inform_L[44][2] = l_cell_wire[41];							inform_L[41][2] = l_cell_wire[42];							inform_L[45][2] = l_cell_wire[43];							inform_L[42][2] = l_cell_wire[44];							inform_L[46][2] = l_cell_wire[45];							inform_L[43][2] = l_cell_wire[46];							inform_L[47][2] = l_cell_wire[47];							inform_L[48][2] = l_cell_wire[48];							inform_L[52][2] = l_cell_wire[49];							inform_L[49][2] = l_cell_wire[50];							inform_L[53][2] = l_cell_wire[51];							inform_L[50][2] = l_cell_wire[52];							inform_L[54][2] = l_cell_wire[53];							inform_L[51][2] = l_cell_wire[54];							inform_L[55][2] = l_cell_wire[55];							inform_L[56][2] = l_cell_wire[56];							inform_L[60][2] = l_cell_wire[57];							inform_L[57][2] = l_cell_wire[58];							inform_L[61][2] = l_cell_wire[59];							inform_L[58][2] = l_cell_wire[60];							inform_L[62][2] = l_cell_wire[61];							inform_L[59][2] = l_cell_wire[62];							inform_L[63][2] = l_cell_wire[63];							inform_L[64][2] = l_cell_wire[64];							inform_L[68][2] = l_cell_wire[65];							inform_L[65][2] = l_cell_wire[66];							inform_L[69][2] = l_cell_wire[67];							inform_L[66][2] = l_cell_wire[68];							inform_L[70][2] = l_cell_wire[69];							inform_L[67][2] = l_cell_wire[70];							inform_L[71][2] = l_cell_wire[71];							inform_L[72][2] = l_cell_wire[72];							inform_L[76][2] = l_cell_wire[73];							inform_L[73][2] = l_cell_wire[74];							inform_L[77][2] = l_cell_wire[75];							inform_L[74][2] = l_cell_wire[76];							inform_L[78][2] = l_cell_wire[77];							inform_L[75][2] = l_cell_wire[78];							inform_L[79][2] = l_cell_wire[79];							inform_L[80][2] = l_cell_wire[80];							inform_L[84][2] = l_cell_wire[81];							inform_L[81][2] = l_cell_wire[82];							inform_L[85][2] = l_cell_wire[83];							inform_L[82][2] = l_cell_wire[84];							inform_L[86][2] = l_cell_wire[85];							inform_L[83][2] = l_cell_wire[86];							inform_L[87][2] = l_cell_wire[87];							inform_L[88][2] = l_cell_wire[88];							inform_L[92][2] = l_cell_wire[89];							inform_L[89][2] = l_cell_wire[90];							inform_L[93][2] = l_cell_wire[91];							inform_L[90][2] = l_cell_wire[92];							inform_L[94][2] = l_cell_wire[93];							inform_L[91][2] = l_cell_wire[94];							inform_L[95][2] = l_cell_wire[95];							inform_L[96][2] = l_cell_wire[96];							inform_L[100][2] = l_cell_wire[97];							inform_L[97][2] = l_cell_wire[98];							inform_L[101][2] = l_cell_wire[99];							inform_L[98][2] = l_cell_wire[100];							inform_L[102][2] = l_cell_wire[101];							inform_L[99][2] = l_cell_wire[102];							inform_L[103][2] = l_cell_wire[103];							inform_L[104][2] = l_cell_wire[104];							inform_L[108][2] = l_cell_wire[105];							inform_L[105][2] = l_cell_wire[106];							inform_L[109][2] = l_cell_wire[107];							inform_L[106][2] = l_cell_wire[108];							inform_L[110][2] = l_cell_wire[109];							inform_L[107][2] = l_cell_wire[110];							inform_L[111][2] = l_cell_wire[111];							inform_L[112][2] = l_cell_wire[112];							inform_L[116][2] = l_cell_wire[113];							inform_L[113][2] = l_cell_wire[114];							inform_L[117][2] = l_cell_wire[115];							inform_L[114][2] = l_cell_wire[116];							inform_L[118][2] = l_cell_wire[117];							inform_L[115][2] = l_cell_wire[118];							inform_L[119][2] = l_cell_wire[119];							inform_L[120][2] = l_cell_wire[120];							inform_L[124][2] = l_cell_wire[121];							inform_L[121][2] = l_cell_wire[122];							inform_L[125][2] = l_cell_wire[123];							inform_L[122][2] = l_cell_wire[124];							inform_L[126][2] = l_cell_wire[125];							inform_L[123][2] = l_cell_wire[126];							inform_L[127][2] = l_cell_wire[127];							inform_L[128][2] = l_cell_wire[128];							inform_L[132][2] = l_cell_wire[129];							inform_L[129][2] = l_cell_wire[130];							inform_L[133][2] = l_cell_wire[131];							inform_L[130][2] = l_cell_wire[132];							inform_L[134][2] = l_cell_wire[133];							inform_L[131][2] = l_cell_wire[134];							inform_L[135][2] = l_cell_wire[135];							inform_L[136][2] = l_cell_wire[136];							inform_L[140][2] = l_cell_wire[137];							inform_L[137][2] = l_cell_wire[138];							inform_L[141][2] = l_cell_wire[139];							inform_L[138][2] = l_cell_wire[140];							inform_L[142][2] = l_cell_wire[141];							inform_L[139][2] = l_cell_wire[142];							inform_L[143][2] = l_cell_wire[143];							inform_L[144][2] = l_cell_wire[144];							inform_L[148][2] = l_cell_wire[145];							inform_L[145][2] = l_cell_wire[146];							inform_L[149][2] = l_cell_wire[147];							inform_L[146][2] = l_cell_wire[148];							inform_L[150][2] = l_cell_wire[149];							inform_L[147][2] = l_cell_wire[150];							inform_L[151][2] = l_cell_wire[151];							inform_L[152][2] = l_cell_wire[152];							inform_L[156][2] = l_cell_wire[153];							inform_L[153][2] = l_cell_wire[154];							inform_L[157][2] = l_cell_wire[155];							inform_L[154][2] = l_cell_wire[156];							inform_L[158][2] = l_cell_wire[157];							inform_L[155][2] = l_cell_wire[158];							inform_L[159][2] = l_cell_wire[159];							inform_L[160][2] = l_cell_wire[160];							inform_L[164][2] = l_cell_wire[161];							inform_L[161][2] = l_cell_wire[162];							inform_L[165][2] = l_cell_wire[163];							inform_L[162][2] = l_cell_wire[164];							inform_L[166][2] = l_cell_wire[165];							inform_L[163][2] = l_cell_wire[166];							inform_L[167][2] = l_cell_wire[167];							inform_L[168][2] = l_cell_wire[168];							inform_L[172][2] = l_cell_wire[169];							inform_L[169][2] = l_cell_wire[170];							inform_L[173][2] = l_cell_wire[171];							inform_L[170][2] = l_cell_wire[172];							inform_L[174][2] = l_cell_wire[173];							inform_L[171][2] = l_cell_wire[174];							inform_L[175][2] = l_cell_wire[175];							inform_L[176][2] = l_cell_wire[176];							inform_L[180][2] = l_cell_wire[177];							inform_L[177][2] = l_cell_wire[178];							inform_L[181][2] = l_cell_wire[179];							inform_L[178][2] = l_cell_wire[180];							inform_L[182][2] = l_cell_wire[181];							inform_L[179][2] = l_cell_wire[182];							inform_L[183][2] = l_cell_wire[183];							inform_L[184][2] = l_cell_wire[184];							inform_L[188][2] = l_cell_wire[185];							inform_L[185][2] = l_cell_wire[186];							inform_L[189][2] = l_cell_wire[187];							inform_L[186][2] = l_cell_wire[188];							inform_L[190][2] = l_cell_wire[189];							inform_L[187][2] = l_cell_wire[190];							inform_L[191][2] = l_cell_wire[191];							inform_L[192][2] = l_cell_wire[192];							inform_L[196][2] = l_cell_wire[193];							inform_L[193][2] = l_cell_wire[194];							inform_L[197][2] = l_cell_wire[195];							inform_L[194][2] = l_cell_wire[196];							inform_L[198][2] = l_cell_wire[197];							inform_L[195][2] = l_cell_wire[198];							inform_L[199][2] = l_cell_wire[199];							inform_L[200][2] = l_cell_wire[200];							inform_L[204][2] = l_cell_wire[201];							inform_L[201][2] = l_cell_wire[202];							inform_L[205][2] = l_cell_wire[203];							inform_L[202][2] = l_cell_wire[204];							inform_L[206][2] = l_cell_wire[205];							inform_L[203][2] = l_cell_wire[206];							inform_L[207][2] = l_cell_wire[207];							inform_L[208][2] = l_cell_wire[208];							inform_L[212][2] = l_cell_wire[209];							inform_L[209][2] = l_cell_wire[210];							inform_L[213][2] = l_cell_wire[211];							inform_L[210][2] = l_cell_wire[212];							inform_L[214][2] = l_cell_wire[213];							inform_L[211][2] = l_cell_wire[214];							inform_L[215][2] = l_cell_wire[215];							inform_L[216][2] = l_cell_wire[216];							inform_L[220][2] = l_cell_wire[217];							inform_L[217][2] = l_cell_wire[218];							inform_L[221][2] = l_cell_wire[219];							inform_L[218][2] = l_cell_wire[220];							inform_L[222][2] = l_cell_wire[221];							inform_L[219][2] = l_cell_wire[222];							inform_L[223][2] = l_cell_wire[223];							inform_L[224][2] = l_cell_wire[224];							inform_L[228][2] = l_cell_wire[225];							inform_L[225][2] = l_cell_wire[226];							inform_L[229][2] = l_cell_wire[227];							inform_L[226][2] = l_cell_wire[228];							inform_L[230][2] = l_cell_wire[229];							inform_L[227][2] = l_cell_wire[230];							inform_L[231][2] = l_cell_wire[231];							inform_L[232][2] = l_cell_wire[232];							inform_L[236][2] = l_cell_wire[233];							inform_L[233][2] = l_cell_wire[234];							inform_L[237][2] = l_cell_wire[235];							inform_L[234][2] = l_cell_wire[236];							inform_L[238][2] = l_cell_wire[237];							inform_L[235][2] = l_cell_wire[238];							inform_L[239][2] = l_cell_wire[239];							inform_L[240][2] = l_cell_wire[240];							inform_L[244][2] = l_cell_wire[241];							inform_L[241][2] = l_cell_wire[242];							inform_L[245][2] = l_cell_wire[243];							inform_L[242][2] = l_cell_wire[244];							inform_L[246][2] = l_cell_wire[245];							inform_L[243][2] = l_cell_wire[246];							inform_L[247][2] = l_cell_wire[247];							inform_L[248][2] = l_cell_wire[248];							inform_L[252][2] = l_cell_wire[249];							inform_L[249][2] = l_cell_wire[250];							inform_L[253][2] = l_cell_wire[251];							inform_L[250][2] = l_cell_wire[252];							inform_L[254][2] = l_cell_wire[253];							inform_L[251][2] = l_cell_wire[254];							inform_L[255][2] = l_cell_wire[255];							inform_L[256][2] = l_cell_wire[256];							inform_L[260][2] = l_cell_wire[257];							inform_L[257][2] = l_cell_wire[258];							inform_L[261][2] = l_cell_wire[259];							inform_L[258][2] = l_cell_wire[260];							inform_L[262][2] = l_cell_wire[261];							inform_L[259][2] = l_cell_wire[262];							inform_L[263][2] = l_cell_wire[263];							inform_L[264][2] = l_cell_wire[264];							inform_L[268][2] = l_cell_wire[265];							inform_L[265][2] = l_cell_wire[266];							inform_L[269][2] = l_cell_wire[267];							inform_L[266][2] = l_cell_wire[268];							inform_L[270][2] = l_cell_wire[269];							inform_L[267][2] = l_cell_wire[270];							inform_L[271][2] = l_cell_wire[271];							inform_L[272][2] = l_cell_wire[272];							inform_L[276][2] = l_cell_wire[273];							inform_L[273][2] = l_cell_wire[274];							inform_L[277][2] = l_cell_wire[275];							inform_L[274][2] = l_cell_wire[276];							inform_L[278][2] = l_cell_wire[277];							inform_L[275][2] = l_cell_wire[278];							inform_L[279][2] = l_cell_wire[279];							inform_L[280][2] = l_cell_wire[280];							inform_L[284][2] = l_cell_wire[281];							inform_L[281][2] = l_cell_wire[282];							inform_L[285][2] = l_cell_wire[283];							inform_L[282][2] = l_cell_wire[284];							inform_L[286][2] = l_cell_wire[285];							inform_L[283][2] = l_cell_wire[286];							inform_L[287][2] = l_cell_wire[287];							inform_L[288][2] = l_cell_wire[288];							inform_L[292][2] = l_cell_wire[289];							inform_L[289][2] = l_cell_wire[290];							inform_L[293][2] = l_cell_wire[291];							inform_L[290][2] = l_cell_wire[292];							inform_L[294][2] = l_cell_wire[293];							inform_L[291][2] = l_cell_wire[294];							inform_L[295][2] = l_cell_wire[295];							inform_L[296][2] = l_cell_wire[296];							inform_L[300][2] = l_cell_wire[297];							inform_L[297][2] = l_cell_wire[298];							inform_L[301][2] = l_cell_wire[299];							inform_L[298][2] = l_cell_wire[300];							inform_L[302][2] = l_cell_wire[301];							inform_L[299][2] = l_cell_wire[302];							inform_L[303][2] = l_cell_wire[303];							inform_L[304][2] = l_cell_wire[304];							inform_L[308][2] = l_cell_wire[305];							inform_L[305][2] = l_cell_wire[306];							inform_L[309][2] = l_cell_wire[307];							inform_L[306][2] = l_cell_wire[308];							inform_L[310][2] = l_cell_wire[309];							inform_L[307][2] = l_cell_wire[310];							inform_L[311][2] = l_cell_wire[311];							inform_L[312][2] = l_cell_wire[312];							inform_L[316][2] = l_cell_wire[313];							inform_L[313][2] = l_cell_wire[314];							inform_L[317][2] = l_cell_wire[315];							inform_L[314][2] = l_cell_wire[316];							inform_L[318][2] = l_cell_wire[317];							inform_L[315][2] = l_cell_wire[318];							inform_L[319][2] = l_cell_wire[319];							inform_L[320][2] = l_cell_wire[320];							inform_L[324][2] = l_cell_wire[321];							inform_L[321][2] = l_cell_wire[322];							inform_L[325][2] = l_cell_wire[323];							inform_L[322][2] = l_cell_wire[324];							inform_L[326][2] = l_cell_wire[325];							inform_L[323][2] = l_cell_wire[326];							inform_L[327][2] = l_cell_wire[327];							inform_L[328][2] = l_cell_wire[328];							inform_L[332][2] = l_cell_wire[329];							inform_L[329][2] = l_cell_wire[330];							inform_L[333][2] = l_cell_wire[331];							inform_L[330][2] = l_cell_wire[332];							inform_L[334][2] = l_cell_wire[333];							inform_L[331][2] = l_cell_wire[334];							inform_L[335][2] = l_cell_wire[335];							inform_L[336][2] = l_cell_wire[336];							inform_L[340][2] = l_cell_wire[337];							inform_L[337][2] = l_cell_wire[338];							inform_L[341][2] = l_cell_wire[339];							inform_L[338][2] = l_cell_wire[340];							inform_L[342][2] = l_cell_wire[341];							inform_L[339][2] = l_cell_wire[342];							inform_L[343][2] = l_cell_wire[343];							inform_L[344][2] = l_cell_wire[344];							inform_L[348][2] = l_cell_wire[345];							inform_L[345][2] = l_cell_wire[346];							inform_L[349][2] = l_cell_wire[347];							inform_L[346][2] = l_cell_wire[348];							inform_L[350][2] = l_cell_wire[349];							inform_L[347][2] = l_cell_wire[350];							inform_L[351][2] = l_cell_wire[351];							inform_L[352][2] = l_cell_wire[352];							inform_L[356][2] = l_cell_wire[353];							inform_L[353][2] = l_cell_wire[354];							inform_L[357][2] = l_cell_wire[355];							inform_L[354][2] = l_cell_wire[356];							inform_L[358][2] = l_cell_wire[357];							inform_L[355][2] = l_cell_wire[358];							inform_L[359][2] = l_cell_wire[359];							inform_L[360][2] = l_cell_wire[360];							inform_L[364][2] = l_cell_wire[361];							inform_L[361][2] = l_cell_wire[362];							inform_L[365][2] = l_cell_wire[363];							inform_L[362][2] = l_cell_wire[364];							inform_L[366][2] = l_cell_wire[365];							inform_L[363][2] = l_cell_wire[366];							inform_L[367][2] = l_cell_wire[367];							inform_L[368][2] = l_cell_wire[368];							inform_L[372][2] = l_cell_wire[369];							inform_L[369][2] = l_cell_wire[370];							inform_L[373][2] = l_cell_wire[371];							inform_L[370][2] = l_cell_wire[372];							inform_L[374][2] = l_cell_wire[373];							inform_L[371][2] = l_cell_wire[374];							inform_L[375][2] = l_cell_wire[375];							inform_L[376][2] = l_cell_wire[376];							inform_L[380][2] = l_cell_wire[377];							inform_L[377][2] = l_cell_wire[378];							inform_L[381][2] = l_cell_wire[379];							inform_L[378][2] = l_cell_wire[380];							inform_L[382][2] = l_cell_wire[381];							inform_L[379][2] = l_cell_wire[382];							inform_L[383][2] = l_cell_wire[383];							inform_L[384][2] = l_cell_wire[384];							inform_L[388][2] = l_cell_wire[385];							inform_L[385][2] = l_cell_wire[386];							inform_L[389][2] = l_cell_wire[387];							inform_L[386][2] = l_cell_wire[388];							inform_L[390][2] = l_cell_wire[389];							inform_L[387][2] = l_cell_wire[390];							inform_L[391][2] = l_cell_wire[391];							inform_L[392][2] = l_cell_wire[392];							inform_L[396][2] = l_cell_wire[393];							inform_L[393][2] = l_cell_wire[394];							inform_L[397][2] = l_cell_wire[395];							inform_L[394][2] = l_cell_wire[396];							inform_L[398][2] = l_cell_wire[397];							inform_L[395][2] = l_cell_wire[398];							inform_L[399][2] = l_cell_wire[399];							inform_L[400][2] = l_cell_wire[400];							inform_L[404][2] = l_cell_wire[401];							inform_L[401][2] = l_cell_wire[402];							inform_L[405][2] = l_cell_wire[403];							inform_L[402][2] = l_cell_wire[404];							inform_L[406][2] = l_cell_wire[405];							inform_L[403][2] = l_cell_wire[406];							inform_L[407][2] = l_cell_wire[407];							inform_L[408][2] = l_cell_wire[408];							inform_L[412][2] = l_cell_wire[409];							inform_L[409][2] = l_cell_wire[410];							inform_L[413][2] = l_cell_wire[411];							inform_L[410][2] = l_cell_wire[412];							inform_L[414][2] = l_cell_wire[413];							inform_L[411][2] = l_cell_wire[414];							inform_L[415][2] = l_cell_wire[415];							inform_L[416][2] = l_cell_wire[416];							inform_L[420][2] = l_cell_wire[417];							inform_L[417][2] = l_cell_wire[418];							inform_L[421][2] = l_cell_wire[419];							inform_L[418][2] = l_cell_wire[420];							inform_L[422][2] = l_cell_wire[421];							inform_L[419][2] = l_cell_wire[422];							inform_L[423][2] = l_cell_wire[423];							inform_L[424][2] = l_cell_wire[424];							inform_L[428][2] = l_cell_wire[425];							inform_L[425][2] = l_cell_wire[426];							inform_L[429][2] = l_cell_wire[427];							inform_L[426][2] = l_cell_wire[428];							inform_L[430][2] = l_cell_wire[429];							inform_L[427][2] = l_cell_wire[430];							inform_L[431][2] = l_cell_wire[431];							inform_L[432][2] = l_cell_wire[432];							inform_L[436][2] = l_cell_wire[433];							inform_L[433][2] = l_cell_wire[434];							inform_L[437][2] = l_cell_wire[435];							inform_L[434][2] = l_cell_wire[436];							inform_L[438][2] = l_cell_wire[437];							inform_L[435][2] = l_cell_wire[438];							inform_L[439][2] = l_cell_wire[439];							inform_L[440][2] = l_cell_wire[440];							inform_L[444][2] = l_cell_wire[441];							inform_L[441][2] = l_cell_wire[442];							inform_L[445][2] = l_cell_wire[443];							inform_L[442][2] = l_cell_wire[444];							inform_L[446][2] = l_cell_wire[445];							inform_L[443][2] = l_cell_wire[446];							inform_L[447][2] = l_cell_wire[447];							inform_L[448][2] = l_cell_wire[448];							inform_L[452][2] = l_cell_wire[449];							inform_L[449][2] = l_cell_wire[450];							inform_L[453][2] = l_cell_wire[451];							inform_L[450][2] = l_cell_wire[452];							inform_L[454][2] = l_cell_wire[453];							inform_L[451][2] = l_cell_wire[454];							inform_L[455][2] = l_cell_wire[455];							inform_L[456][2] = l_cell_wire[456];							inform_L[460][2] = l_cell_wire[457];							inform_L[457][2] = l_cell_wire[458];							inform_L[461][2] = l_cell_wire[459];							inform_L[458][2] = l_cell_wire[460];							inform_L[462][2] = l_cell_wire[461];							inform_L[459][2] = l_cell_wire[462];							inform_L[463][2] = l_cell_wire[463];							inform_L[464][2] = l_cell_wire[464];							inform_L[468][2] = l_cell_wire[465];							inform_L[465][2] = l_cell_wire[466];							inform_L[469][2] = l_cell_wire[467];							inform_L[466][2] = l_cell_wire[468];							inform_L[470][2] = l_cell_wire[469];							inform_L[467][2] = l_cell_wire[470];							inform_L[471][2] = l_cell_wire[471];							inform_L[472][2] = l_cell_wire[472];							inform_L[476][2] = l_cell_wire[473];							inform_L[473][2] = l_cell_wire[474];							inform_L[477][2] = l_cell_wire[475];							inform_L[474][2] = l_cell_wire[476];							inform_L[478][2] = l_cell_wire[477];							inform_L[475][2] = l_cell_wire[478];							inform_L[479][2] = l_cell_wire[479];							inform_L[480][2] = l_cell_wire[480];							inform_L[484][2] = l_cell_wire[481];							inform_L[481][2] = l_cell_wire[482];							inform_L[485][2] = l_cell_wire[483];							inform_L[482][2] = l_cell_wire[484];							inform_L[486][2] = l_cell_wire[485];							inform_L[483][2] = l_cell_wire[486];							inform_L[487][2] = l_cell_wire[487];							inform_L[488][2] = l_cell_wire[488];							inform_L[492][2] = l_cell_wire[489];							inform_L[489][2] = l_cell_wire[490];							inform_L[493][2] = l_cell_wire[491];							inform_L[490][2] = l_cell_wire[492];							inform_L[494][2] = l_cell_wire[493];							inform_L[491][2] = l_cell_wire[494];							inform_L[495][2] = l_cell_wire[495];							inform_L[496][2] = l_cell_wire[496];							inform_L[500][2] = l_cell_wire[497];							inform_L[497][2] = l_cell_wire[498];							inform_L[501][2] = l_cell_wire[499];							inform_L[498][2] = l_cell_wire[500];							inform_L[502][2] = l_cell_wire[501];							inform_L[499][2] = l_cell_wire[502];							inform_L[503][2] = l_cell_wire[503];							inform_L[504][2] = l_cell_wire[504];							inform_L[508][2] = l_cell_wire[505];							inform_L[505][2] = l_cell_wire[506];							inform_L[509][2] = l_cell_wire[507];							inform_L[506][2] = l_cell_wire[508];							inform_L[510][2] = l_cell_wire[509];							inform_L[507][2] = l_cell_wire[510];							inform_L[511][2] = l_cell_wire[511];							inform_L[512][2] = l_cell_wire[512];							inform_L[516][2] = l_cell_wire[513];							inform_L[513][2] = l_cell_wire[514];							inform_L[517][2] = l_cell_wire[515];							inform_L[514][2] = l_cell_wire[516];							inform_L[518][2] = l_cell_wire[517];							inform_L[515][2] = l_cell_wire[518];							inform_L[519][2] = l_cell_wire[519];							inform_L[520][2] = l_cell_wire[520];							inform_L[524][2] = l_cell_wire[521];							inform_L[521][2] = l_cell_wire[522];							inform_L[525][2] = l_cell_wire[523];							inform_L[522][2] = l_cell_wire[524];							inform_L[526][2] = l_cell_wire[525];							inform_L[523][2] = l_cell_wire[526];							inform_L[527][2] = l_cell_wire[527];							inform_L[528][2] = l_cell_wire[528];							inform_L[532][2] = l_cell_wire[529];							inform_L[529][2] = l_cell_wire[530];							inform_L[533][2] = l_cell_wire[531];							inform_L[530][2] = l_cell_wire[532];							inform_L[534][2] = l_cell_wire[533];							inform_L[531][2] = l_cell_wire[534];							inform_L[535][2] = l_cell_wire[535];							inform_L[536][2] = l_cell_wire[536];							inform_L[540][2] = l_cell_wire[537];							inform_L[537][2] = l_cell_wire[538];							inform_L[541][2] = l_cell_wire[539];							inform_L[538][2] = l_cell_wire[540];							inform_L[542][2] = l_cell_wire[541];							inform_L[539][2] = l_cell_wire[542];							inform_L[543][2] = l_cell_wire[543];							inform_L[544][2] = l_cell_wire[544];							inform_L[548][2] = l_cell_wire[545];							inform_L[545][2] = l_cell_wire[546];							inform_L[549][2] = l_cell_wire[547];							inform_L[546][2] = l_cell_wire[548];							inform_L[550][2] = l_cell_wire[549];							inform_L[547][2] = l_cell_wire[550];							inform_L[551][2] = l_cell_wire[551];							inform_L[552][2] = l_cell_wire[552];							inform_L[556][2] = l_cell_wire[553];							inform_L[553][2] = l_cell_wire[554];							inform_L[557][2] = l_cell_wire[555];							inform_L[554][2] = l_cell_wire[556];							inform_L[558][2] = l_cell_wire[557];							inform_L[555][2] = l_cell_wire[558];							inform_L[559][2] = l_cell_wire[559];							inform_L[560][2] = l_cell_wire[560];							inform_L[564][2] = l_cell_wire[561];							inform_L[561][2] = l_cell_wire[562];							inform_L[565][2] = l_cell_wire[563];							inform_L[562][2] = l_cell_wire[564];							inform_L[566][2] = l_cell_wire[565];							inform_L[563][2] = l_cell_wire[566];							inform_L[567][2] = l_cell_wire[567];							inform_L[568][2] = l_cell_wire[568];							inform_L[572][2] = l_cell_wire[569];							inform_L[569][2] = l_cell_wire[570];							inform_L[573][2] = l_cell_wire[571];							inform_L[570][2] = l_cell_wire[572];							inform_L[574][2] = l_cell_wire[573];							inform_L[571][2] = l_cell_wire[574];							inform_L[575][2] = l_cell_wire[575];							inform_L[576][2] = l_cell_wire[576];							inform_L[580][2] = l_cell_wire[577];							inform_L[577][2] = l_cell_wire[578];							inform_L[581][2] = l_cell_wire[579];							inform_L[578][2] = l_cell_wire[580];							inform_L[582][2] = l_cell_wire[581];							inform_L[579][2] = l_cell_wire[582];							inform_L[583][2] = l_cell_wire[583];							inform_L[584][2] = l_cell_wire[584];							inform_L[588][2] = l_cell_wire[585];							inform_L[585][2] = l_cell_wire[586];							inform_L[589][2] = l_cell_wire[587];							inform_L[586][2] = l_cell_wire[588];							inform_L[590][2] = l_cell_wire[589];							inform_L[587][2] = l_cell_wire[590];							inform_L[591][2] = l_cell_wire[591];							inform_L[592][2] = l_cell_wire[592];							inform_L[596][2] = l_cell_wire[593];							inform_L[593][2] = l_cell_wire[594];							inform_L[597][2] = l_cell_wire[595];							inform_L[594][2] = l_cell_wire[596];							inform_L[598][2] = l_cell_wire[597];							inform_L[595][2] = l_cell_wire[598];							inform_L[599][2] = l_cell_wire[599];							inform_L[600][2] = l_cell_wire[600];							inform_L[604][2] = l_cell_wire[601];							inform_L[601][2] = l_cell_wire[602];							inform_L[605][2] = l_cell_wire[603];							inform_L[602][2] = l_cell_wire[604];							inform_L[606][2] = l_cell_wire[605];							inform_L[603][2] = l_cell_wire[606];							inform_L[607][2] = l_cell_wire[607];							inform_L[608][2] = l_cell_wire[608];							inform_L[612][2] = l_cell_wire[609];							inform_L[609][2] = l_cell_wire[610];							inform_L[613][2] = l_cell_wire[611];							inform_L[610][2] = l_cell_wire[612];							inform_L[614][2] = l_cell_wire[613];							inform_L[611][2] = l_cell_wire[614];							inform_L[615][2] = l_cell_wire[615];							inform_L[616][2] = l_cell_wire[616];							inform_L[620][2] = l_cell_wire[617];							inform_L[617][2] = l_cell_wire[618];							inform_L[621][2] = l_cell_wire[619];							inform_L[618][2] = l_cell_wire[620];							inform_L[622][2] = l_cell_wire[621];							inform_L[619][2] = l_cell_wire[622];							inform_L[623][2] = l_cell_wire[623];							inform_L[624][2] = l_cell_wire[624];							inform_L[628][2] = l_cell_wire[625];							inform_L[625][2] = l_cell_wire[626];							inform_L[629][2] = l_cell_wire[627];							inform_L[626][2] = l_cell_wire[628];							inform_L[630][2] = l_cell_wire[629];							inform_L[627][2] = l_cell_wire[630];							inform_L[631][2] = l_cell_wire[631];							inform_L[632][2] = l_cell_wire[632];							inform_L[636][2] = l_cell_wire[633];							inform_L[633][2] = l_cell_wire[634];							inform_L[637][2] = l_cell_wire[635];							inform_L[634][2] = l_cell_wire[636];							inform_L[638][2] = l_cell_wire[637];							inform_L[635][2] = l_cell_wire[638];							inform_L[639][2] = l_cell_wire[639];							inform_L[640][2] = l_cell_wire[640];							inform_L[644][2] = l_cell_wire[641];							inform_L[641][2] = l_cell_wire[642];							inform_L[645][2] = l_cell_wire[643];							inform_L[642][2] = l_cell_wire[644];							inform_L[646][2] = l_cell_wire[645];							inform_L[643][2] = l_cell_wire[646];							inform_L[647][2] = l_cell_wire[647];							inform_L[648][2] = l_cell_wire[648];							inform_L[652][2] = l_cell_wire[649];							inform_L[649][2] = l_cell_wire[650];							inform_L[653][2] = l_cell_wire[651];							inform_L[650][2] = l_cell_wire[652];							inform_L[654][2] = l_cell_wire[653];							inform_L[651][2] = l_cell_wire[654];							inform_L[655][2] = l_cell_wire[655];							inform_L[656][2] = l_cell_wire[656];							inform_L[660][2] = l_cell_wire[657];							inform_L[657][2] = l_cell_wire[658];							inform_L[661][2] = l_cell_wire[659];							inform_L[658][2] = l_cell_wire[660];							inform_L[662][2] = l_cell_wire[661];							inform_L[659][2] = l_cell_wire[662];							inform_L[663][2] = l_cell_wire[663];							inform_L[664][2] = l_cell_wire[664];							inform_L[668][2] = l_cell_wire[665];							inform_L[665][2] = l_cell_wire[666];							inform_L[669][2] = l_cell_wire[667];							inform_L[666][2] = l_cell_wire[668];							inform_L[670][2] = l_cell_wire[669];							inform_L[667][2] = l_cell_wire[670];							inform_L[671][2] = l_cell_wire[671];							inform_L[672][2] = l_cell_wire[672];							inform_L[676][2] = l_cell_wire[673];							inform_L[673][2] = l_cell_wire[674];							inform_L[677][2] = l_cell_wire[675];							inform_L[674][2] = l_cell_wire[676];							inform_L[678][2] = l_cell_wire[677];							inform_L[675][2] = l_cell_wire[678];							inform_L[679][2] = l_cell_wire[679];							inform_L[680][2] = l_cell_wire[680];							inform_L[684][2] = l_cell_wire[681];							inform_L[681][2] = l_cell_wire[682];							inform_L[685][2] = l_cell_wire[683];							inform_L[682][2] = l_cell_wire[684];							inform_L[686][2] = l_cell_wire[685];							inform_L[683][2] = l_cell_wire[686];							inform_L[687][2] = l_cell_wire[687];							inform_L[688][2] = l_cell_wire[688];							inform_L[692][2] = l_cell_wire[689];							inform_L[689][2] = l_cell_wire[690];							inform_L[693][2] = l_cell_wire[691];							inform_L[690][2] = l_cell_wire[692];							inform_L[694][2] = l_cell_wire[693];							inform_L[691][2] = l_cell_wire[694];							inform_L[695][2] = l_cell_wire[695];							inform_L[696][2] = l_cell_wire[696];							inform_L[700][2] = l_cell_wire[697];							inform_L[697][2] = l_cell_wire[698];							inform_L[701][2] = l_cell_wire[699];							inform_L[698][2] = l_cell_wire[700];							inform_L[702][2] = l_cell_wire[701];							inform_L[699][2] = l_cell_wire[702];							inform_L[703][2] = l_cell_wire[703];							inform_L[704][2] = l_cell_wire[704];							inform_L[708][2] = l_cell_wire[705];							inform_L[705][2] = l_cell_wire[706];							inform_L[709][2] = l_cell_wire[707];							inform_L[706][2] = l_cell_wire[708];							inform_L[710][2] = l_cell_wire[709];							inform_L[707][2] = l_cell_wire[710];							inform_L[711][2] = l_cell_wire[711];							inform_L[712][2] = l_cell_wire[712];							inform_L[716][2] = l_cell_wire[713];							inform_L[713][2] = l_cell_wire[714];							inform_L[717][2] = l_cell_wire[715];							inform_L[714][2] = l_cell_wire[716];							inform_L[718][2] = l_cell_wire[717];							inform_L[715][2] = l_cell_wire[718];							inform_L[719][2] = l_cell_wire[719];							inform_L[720][2] = l_cell_wire[720];							inform_L[724][2] = l_cell_wire[721];							inform_L[721][2] = l_cell_wire[722];							inform_L[725][2] = l_cell_wire[723];							inform_L[722][2] = l_cell_wire[724];							inform_L[726][2] = l_cell_wire[725];							inform_L[723][2] = l_cell_wire[726];							inform_L[727][2] = l_cell_wire[727];							inform_L[728][2] = l_cell_wire[728];							inform_L[732][2] = l_cell_wire[729];							inform_L[729][2] = l_cell_wire[730];							inform_L[733][2] = l_cell_wire[731];							inform_L[730][2] = l_cell_wire[732];							inform_L[734][2] = l_cell_wire[733];							inform_L[731][2] = l_cell_wire[734];							inform_L[735][2] = l_cell_wire[735];							inform_L[736][2] = l_cell_wire[736];							inform_L[740][2] = l_cell_wire[737];							inform_L[737][2] = l_cell_wire[738];							inform_L[741][2] = l_cell_wire[739];							inform_L[738][2] = l_cell_wire[740];							inform_L[742][2] = l_cell_wire[741];							inform_L[739][2] = l_cell_wire[742];							inform_L[743][2] = l_cell_wire[743];							inform_L[744][2] = l_cell_wire[744];							inform_L[748][2] = l_cell_wire[745];							inform_L[745][2] = l_cell_wire[746];							inform_L[749][2] = l_cell_wire[747];							inform_L[746][2] = l_cell_wire[748];							inform_L[750][2] = l_cell_wire[749];							inform_L[747][2] = l_cell_wire[750];							inform_L[751][2] = l_cell_wire[751];							inform_L[752][2] = l_cell_wire[752];							inform_L[756][2] = l_cell_wire[753];							inform_L[753][2] = l_cell_wire[754];							inform_L[757][2] = l_cell_wire[755];							inform_L[754][2] = l_cell_wire[756];							inform_L[758][2] = l_cell_wire[757];							inform_L[755][2] = l_cell_wire[758];							inform_L[759][2] = l_cell_wire[759];							inform_L[760][2] = l_cell_wire[760];							inform_L[764][2] = l_cell_wire[761];							inform_L[761][2] = l_cell_wire[762];							inform_L[765][2] = l_cell_wire[763];							inform_L[762][2] = l_cell_wire[764];							inform_L[766][2] = l_cell_wire[765];							inform_L[763][2] = l_cell_wire[766];							inform_L[767][2] = l_cell_wire[767];							inform_L[768][2] = l_cell_wire[768];							inform_L[772][2] = l_cell_wire[769];							inform_L[769][2] = l_cell_wire[770];							inform_L[773][2] = l_cell_wire[771];							inform_L[770][2] = l_cell_wire[772];							inform_L[774][2] = l_cell_wire[773];							inform_L[771][2] = l_cell_wire[774];							inform_L[775][2] = l_cell_wire[775];							inform_L[776][2] = l_cell_wire[776];							inform_L[780][2] = l_cell_wire[777];							inform_L[777][2] = l_cell_wire[778];							inform_L[781][2] = l_cell_wire[779];							inform_L[778][2] = l_cell_wire[780];							inform_L[782][2] = l_cell_wire[781];							inform_L[779][2] = l_cell_wire[782];							inform_L[783][2] = l_cell_wire[783];							inform_L[784][2] = l_cell_wire[784];							inform_L[788][2] = l_cell_wire[785];							inform_L[785][2] = l_cell_wire[786];							inform_L[789][2] = l_cell_wire[787];							inform_L[786][2] = l_cell_wire[788];							inform_L[790][2] = l_cell_wire[789];							inform_L[787][2] = l_cell_wire[790];							inform_L[791][2] = l_cell_wire[791];							inform_L[792][2] = l_cell_wire[792];							inform_L[796][2] = l_cell_wire[793];							inform_L[793][2] = l_cell_wire[794];							inform_L[797][2] = l_cell_wire[795];							inform_L[794][2] = l_cell_wire[796];							inform_L[798][2] = l_cell_wire[797];							inform_L[795][2] = l_cell_wire[798];							inform_L[799][2] = l_cell_wire[799];							inform_L[800][2] = l_cell_wire[800];							inform_L[804][2] = l_cell_wire[801];							inform_L[801][2] = l_cell_wire[802];							inform_L[805][2] = l_cell_wire[803];							inform_L[802][2] = l_cell_wire[804];							inform_L[806][2] = l_cell_wire[805];							inform_L[803][2] = l_cell_wire[806];							inform_L[807][2] = l_cell_wire[807];							inform_L[808][2] = l_cell_wire[808];							inform_L[812][2] = l_cell_wire[809];							inform_L[809][2] = l_cell_wire[810];							inform_L[813][2] = l_cell_wire[811];							inform_L[810][2] = l_cell_wire[812];							inform_L[814][2] = l_cell_wire[813];							inform_L[811][2] = l_cell_wire[814];							inform_L[815][2] = l_cell_wire[815];							inform_L[816][2] = l_cell_wire[816];							inform_L[820][2] = l_cell_wire[817];							inform_L[817][2] = l_cell_wire[818];							inform_L[821][2] = l_cell_wire[819];							inform_L[818][2] = l_cell_wire[820];							inform_L[822][2] = l_cell_wire[821];							inform_L[819][2] = l_cell_wire[822];							inform_L[823][2] = l_cell_wire[823];							inform_L[824][2] = l_cell_wire[824];							inform_L[828][2] = l_cell_wire[825];							inform_L[825][2] = l_cell_wire[826];							inform_L[829][2] = l_cell_wire[827];							inform_L[826][2] = l_cell_wire[828];							inform_L[830][2] = l_cell_wire[829];							inform_L[827][2] = l_cell_wire[830];							inform_L[831][2] = l_cell_wire[831];							inform_L[832][2] = l_cell_wire[832];							inform_L[836][2] = l_cell_wire[833];							inform_L[833][2] = l_cell_wire[834];							inform_L[837][2] = l_cell_wire[835];							inform_L[834][2] = l_cell_wire[836];							inform_L[838][2] = l_cell_wire[837];							inform_L[835][2] = l_cell_wire[838];							inform_L[839][2] = l_cell_wire[839];							inform_L[840][2] = l_cell_wire[840];							inform_L[844][2] = l_cell_wire[841];							inform_L[841][2] = l_cell_wire[842];							inform_L[845][2] = l_cell_wire[843];							inform_L[842][2] = l_cell_wire[844];							inform_L[846][2] = l_cell_wire[845];							inform_L[843][2] = l_cell_wire[846];							inform_L[847][2] = l_cell_wire[847];							inform_L[848][2] = l_cell_wire[848];							inform_L[852][2] = l_cell_wire[849];							inform_L[849][2] = l_cell_wire[850];							inform_L[853][2] = l_cell_wire[851];							inform_L[850][2] = l_cell_wire[852];							inform_L[854][2] = l_cell_wire[853];							inform_L[851][2] = l_cell_wire[854];							inform_L[855][2] = l_cell_wire[855];							inform_L[856][2] = l_cell_wire[856];							inform_L[860][2] = l_cell_wire[857];							inform_L[857][2] = l_cell_wire[858];							inform_L[861][2] = l_cell_wire[859];							inform_L[858][2] = l_cell_wire[860];							inform_L[862][2] = l_cell_wire[861];							inform_L[859][2] = l_cell_wire[862];							inform_L[863][2] = l_cell_wire[863];							inform_L[864][2] = l_cell_wire[864];							inform_L[868][2] = l_cell_wire[865];							inform_L[865][2] = l_cell_wire[866];							inform_L[869][2] = l_cell_wire[867];							inform_L[866][2] = l_cell_wire[868];							inform_L[870][2] = l_cell_wire[869];							inform_L[867][2] = l_cell_wire[870];							inform_L[871][2] = l_cell_wire[871];							inform_L[872][2] = l_cell_wire[872];							inform_L[876][2] = l_cell_wire[873];							inform_L[873][2] = l_cell_wire[874];							inform_L[877][2] = l_cell_wire[875];							inform_L[874][2] = l_cell_wire[876];							inform_L[878][2] = l_cell_wire[877];							inform_L[875][2] = l_cell_wire[878];							inform_L[879][2] = l_cell_wire[879];							inform_L[880][2] = l_cell_wire[880];							inform_L[884][2] = l_cell_wire[881];							inform_L[881][2] = l_cell_wire[882];							inform_L[885][2] = l_cell_wire[883];							inform_L[882][2] = l_cell_wire[884];							inform_L[886][2] = l_cell_wire[885];							inform_L[883][2] = l_cell_wire[886];							inform_L[887][2] = l_cell_wire[887];							inform_L[888][2] = l_cell_wire[888];							inform_L[892][2] = l_cell_wire[889];							inform_L[889][2] = l_cell_wire[890];							inform_L[893][2] = l_cell_wire[891];							inform_L[890][2] = l_cell_wire[892];							inform_L[894][2] = l_cell_wire[893];							inform_L[891][2] = l_cell_wire[894];							inform_L[895][2] = l_cell_wire[895];							inform_L[896][2] = l_cell_wire[896];							inform_L[900][2] = l_cell_wire[897];							inform_L[897][2] = l_cell_wire[898];							inform_L[901][2] = l_cell_wire[899];							inform_L[898][2] = l_cell_wire[900];							inform_L[902][2] = l_cell_wire[901];							inform_L[899][2] = l_cell_wire[902];							inform_L[903][2] = l_cell_wire[903];							inform_L[904][2] = l_cell_wire[904];							inform_L[908][2] = l_cell_wire[905];							inform_L[905][2] = l_cell_wire[906];							inform_L[909][2] = l_cell_wire[907];							inform_L[906][2] = l_cell_wire[908];							inform_L[910][2] = l_cell_wire[909];							inform_L[907][2] = l_cell_wire[910];							inform_L[911][2] = l_cell_wire[911];							inform_L[912][2] = l_cell_wire[912];							inform_L[916][2] = l_cell_wire[913];							inform_L[913][2] = l_cell_wire[914];							inform_L[917][2] = l_cell_wire[915];							inform_L[914][2] = l_cell_wire[916];							inform_L[918][2] = l_cell_wire[917];							inform_L[915][2] = l_cell_wire[918];							inform_L[919][2] = l_cell_wire[919];							inform_L[920][2] = l_cell_wire[920];							inform_L[924][2] = l_cell_wire[921];							inform_L[921][2] = l_cell_wire[922];							inform_L[925][2] = l_cell_wire[923];							inform_L[922][2] = l_cell_wire[924];							inform_L[926][2] = l_cell_wire[925];							inform_L[923][2] = l_cell_wire[926];							inform_L[927][2] = l_cell_wire[927];							inform_L[928][2] = l_cell_wire[928];							inform_L[932][2] = l_cell_wire[929];							inform_L[929][2] = l_cell_wire[930];							inform_L[933][2] = l_cell_wire[931];							inform_L[930][2] = l_cell_wire[932];							inform_L[934][2] = l_cell_wire[933];							inform_L[931][2] = l_cell_wire[934];							inform_L[935][2] = l_cell_wire[935];							inform_L[936][2] = l_cell_wire[936];							inform_L[940][2] = l_cell_wire[937];							inform_L[937][2] = l_cell_wire[938];							inform_L[941][2] = l_cell_wire[939];							inform_L[938][2] = l_cell_wire[940];							inform_L[942][2] = l_cell_wire[941];							inform_L[939][2] = l_cell_wire[942];							inform_L[943][2] = l_cell_wire[943];							inform_L[944][2] = l_cell_wire[944];							inform_L[948][2] = l_cell_wire[945];							inform_L[945][2] = l_cell_wire[946];							inform_L[949][2] = l_cell_wire[947];							inform_L[946][2] = l_cell_wire[948];							inform_L[950][2] = l_cell_wire[949];							inform_L[947][2] = l_cell_wire[950];							inform_L[951][2] = l_cell_wire[951];							inform_L[952][2] = l_cell_wire[952];							inform_L[956][2] = l_cell_wire[953];							inform_L[953][2] = l_cell_wire[954];							inform_L[957][2] = l_cell_wire[955];							inform_L[954][2] = l_cell_wire[956];							inform_L[958][2] = l_cell_wire[957];							inform_L[955][2] = l_cell_wire[958];							inform_L[959][2] = l_cell_wire[959];							inform_L[960][2] = l_cell_wire[960];							inform_L[964][2] = l_cell_wire[961];							inform_L[961][2] = l_cell_wire[962];							inform_L[965][2] = l_cell_wire[963];							inform_L[962][2] = l_cell_wire[964];							inform_L[966][2] = l_cell_wire[965];							inform_L[963][2] = l_cell_wire[966];							inform_L[967][2] = l_cell_wire[967];							inform_L[968][2] = l_cell_wire[968];							inform_L[972][2] = l_cell_wire[969];							inform_L[969][2] = l_cell_wire[970];							inform_L[973][2] = l_cell_wire[971];							inform_L[970][2] = l_cell_wire[972];							inform_L[974][2] = l_cell_wire[973];							inform_L[971][2] = l_cell_wire[974];							inform_L[975][2] = l_cell_wire[975];							inform_L[976][2] = l_cell_wire[976];							inform_L[980][2] = l_cell_wire[977];							inform_L[977][2] = l_cell_wire[978];							inform_L[981][2] = l_cell_wire[979];							inform_L[978][2] = l_cell_wire[980];							inform_L[982][2] = l_cell_wire[981];							inform_L[979][2] = l_cell_wire[982];							inform_L[983][2] = l_cell_wire[983];							inform_L[984][2] = l_cell_wire[984];							inform_L[988][2] = l_cell_wire[985];							inform_L[985][2] = l_cell_wire[986];							inform_L[989][2] = l_cell_wire[987];							inform_L[986][2] = l_cell_wire[988];							inform_L[990][2] = l_cell_wire[989];							inform_L[987][2] = l_cell_wire[990];							inform_L[991][2] = l_cell_wire[991];							inform_L[992][2] = l_cell_wire[992];							inform_L[996][2] = l_cell_wire[993];							inform_L[993][2] = l_cell_wire[994];							inform_L[997][2] = l_cell_wire[995];							inform_L[994][2] = l_cell_wire[996];							inform_L[998][2] = l_cell_wire[997];							inform_L[995][2] = l_cell_wire[998];							inform_L[999][2] = l_cell_wire[999];							inform_L[1000][2] = l_cell_wire[1000];							inform_L[1004][2] = l_cell_wire[1001];							inform_L[1001][2] = l_cell_wire[1002];							inform_L[1005][2] = l_cell_wire[1003];							inform_L[1002][2] = l_cell_wire[1004];							inform_L[1006][2] = l_cell_wire[1005];							inform_L[1003][2] = l_cell_wire[1006];							inform_L[1007][2] = l_cell_wire[1007];							inform_L[1008][2] = l_cell_wire[1008];							inform_L[1012][2] = l_cell_wire[1009];							inform_L[1009][2] = l_cell_wire[1010];							inform_L[1013][2] = l_cell_wire[1011];							inform_L[1010][2] = l_cell_wire[1012];							inform_L[1014][2] = l_cell_wire[1013];							inform_L[1011][2] = l_cell_wire[1014];							inform_L[1015][2] = l_cell_wire[1015];							inform_L[1016][2] = l_cell_wire[1016];							inform_L[1020][2] = l_cell_wire[1017];							inform_L[1017][2] = l_cell_wire[1018];							inform_L[1021][2] = l_cell_wire[1019];							inform_L[1018][2] = l_cell_wire[1020];							inform_L[1022][2] = l_cell_wire[1021];							inform_L[1019][2] = l_cell_wire[1022];							inform_L[1023][2] = l_cell_wire[1023];						end
						4:						begin							inform_R[0][4] = r_cell_wire[0];							inform_R[8][4] = r_cell_wire[1];							inform_R[1][4] = r_cell_wire[2];							inform_R[9][4] = r_cell_wire[3];							inform_R[2][4] = r_cell_wire[4];							inform_R[10][4] = r_cell_wire[5];							inform_R[3][4] = r_cell_wire[6];							inform_R[11][4] = r_cell_wire[7];							inform_R[4][4] = r_cell_wire[8];							inform_R[12][4] = r_cell_wire[9];							inform_R[5][4] = r_cell_wire[10];							inform_R[13][4] = r_cell_wire[11];							inform_R[6][4] = r_cell_wire[12];							inform_R[14][4] = r_cell_wire[13];							inform_R[7][4] = r_cell_wire[14];							inform_R[15][4] = r_cell_wire[15];							inform_R[16][4] = r_cell_wire[16];							inform_R[24][4] = r_cell_wire[17];							inform_R[17][4] = r_cell_wire[18];							inform_R[25][4] = r_cell_wire[19];							inform_R[18][4] = r_cell_wire[20];							inform_R[26][4] = r_cell_wire[21];							inform_R[19][4] = r_cell_wire[22];							inform_R[27][4] = r_cell_wire[23];							inform_R[20][4] = r_cell_wire[24];							inform_R[28][4] = r_cell_wire[25];							inform_R[21][4] = r_cell_wire[26];							inform_R[29][4] = r_cell_wire[27];							inform_R[22][4] = r_cell_wire[28];							inform_R[30][4] = r_cell_wire[29];							inform_R[23][4] = r_cell_wire[30];							inform_R[31][4] = r_cell_wire[31];							inform_R[32][4] = r_cell_wire[32];							inform_R[40][4] = r_cell_wire[33];							inform_R[33][4] = r_cell_wire[34];							inform_R[41][4] = r_cell_wire[35];							inform_R[34][4] = r_cell_wire[36];							inform_R[42][4] = r_cell_wire[37];							inform_R[35][4] = r_cell_wire[38];							inform_R[43][4] = r_cell_wire[39];							inform_R[36][4] = r_cell_wire[40];							inform_R[44][4] = r_cell_wire[41];							inform_R[37][4] = r_cell_wire[42];							inform_R[45][4] = r_cell_wire[43];							inform_R[38][4] = r_cell_wire[44];							inform_R[46][4] = r_cell_wire[45];							inform_R[39][4] = r_cell_wire[46];							inform_R[47][4] = r_cell_wire[47];							inform_R[48][4] = r_cell_wire[48];							inform_R[56][4] = r_cell_wire[49];							inform_R[49][4] = r_cell_wire[50];							inform_R[57][4] = r_cell_wire[51];							inform_R[50][4] = r_cell_wire[52];							inform_R[58][4] = r_cell_wire[53];							inform_R[51][4] = r_cell_wire[54];							inform_R[59][4] = r_cell_wire[55];							inform_R[52][4] = r_cell_wire[56];							inform_R[60][4] = r_cell_wire[57];							inform_R[53][4] = r_cell_wire[58];							inform_R[61][4] = r_cell_wire[59];							inform_R[54][4] = r_cell_wire[60];							inform_R[62][4] = r_cell_wire[61];							inform_R[55][4] = r_cell_wire[62];							inform_R[63][4] = r_cell_wire[63];							inform_R[64][4] = r_cell_wire[64];							inform_R[72][4] = r_cell_wire[65];							inform_R[65][4] = r_cell_wire[66];							inform_R[73][4] = r_cell_wire[67];							inform_R[66][4] = r_cell_wire[68];							inform_R[74][4] = r_cell_wire[69];							inform_R[67][4] = r_cell_wire[70];							inform_R[75][4] = r_cell_wire[71];							inform_R[68][4] = r_cell_wire[72];							inform_R[76][4] = r_cell_wire[73];							inform_R[69][4] = r_cell_wire[74];							inform_R[77][4] = r_cell_wire[75];							inform_R[70][4] = r_cell_wire[76];							inform_R[78][4] = r_cell_wire[77];							inform_R[71][4] = r_cell_wire[78];							inform_R[79][4] = r_cell_wire[79];							inform_R[80][4] = r_cell_wire[80];							inform_R[88][4] = r_cell_wire[81];							inform_R[81][4] = r_cell_wire[82];							inform_R[89][4] = r_cell_wire[83];							inform_R[82][4] = r_cell_wire[84];							inform_R[90][4] = r_cell_wire[85];							inform_R[83][4] = r_cell_wire[86];							inform_R[91][4] = r_cell_wire[87];							inform_R[84][4] = r_cell_wire[88];							inform_R[92][4] = r_cell_wire[89];							inform_R[85][4] = r_cell_wire[90];							inform_R[93][4] = r_cell_wire[91];							inform_R[86][4] = r_cell_wire[92];							inform_R[94][4] = r_cell_wire[93];							inform_R[87][4] = r_cell_wire[94];							inform_R[95][4] = r_cell_wire[95];							inform_R[96][4] = r_cell_wire[96];							inform_R[104][4] = r_cell_wire[97];							inform_R[97][4] = r_cell_wire[98];							inform_R[105][4] = r_cell_wire[99];							inform_R[98][4] = r_cell_wire[100];							inform_R[106][4] = r_cell_wire[101];							inform_R[99][4] = r_cell_wire[102];							inform_R[107][4] = r_cell_wire[103];							inform_R[100][4] = r_cell_wire[104];							inform_R[108][4] = r_cell_wire[105];							inform_R[101][4] = r_cell_wire[106];							inform_R[109][4] = r_cell_wire[107];							inform_R[102][4] = r_cell_wire[108];							inform_R[110][4] = r_cell_wire[109];							inform_R[103][4] = r_cell_wire[110];							inform_R[111][4] = r_cell_wire[111];							inform_R[112][4] = r_cell_wire[112];							inform_R[120][4] = r_cell_wire[113];							inform_R[113][4] = r_cell_wire[114];							inform_R[121][4] = r_cell_wire[115];							inform_R[114][4] = r_cell_wire[116];							inform_R[122][4] = r_cell_wire[117];							inform_R[115][4] = r_cell_wire[118];							inform_R[123][4] = r_cell_wire[119];							inform_R[116][4] = r_cell_wire[120];							inform_R[124][4] = r_cell_wire[121];							inform_R[117][4] = r_cell_wire[122];							inform_R[125][4] = r_cell_wire[123];							inform_R[118][4] = r_cell_wire[124];							inform_R[126][4] = r_cell_wire[125];							inform_R[119][4] = r_cell_wire[126];							inform_R[127][4] = r_cell_wire[127];							inform_R[128][4] = r_cell_wire[128];							inform_R[136][4] = r_cell_wire[129];							inform_R[129][4] = r_cell_wire[130];							inform_R[137][4] = r_cell_wire[131];							inform_R[130][4] = r_cell_wire[132];							inform_R[138][4] = r_cell_wire[133];							inform_R[131][4] = r_cell_wire[134];							inform_R[139][4] = r_cell_wire[135];							inform_R[132][4] = r_cell_wire[136];							inform_R[140][4] = r_cell_wire[137];							inform_R[133][4] = r_cell_wire[138];							inform_R[141][4] = r_cell_wire[139];							inform_R[134][4] = r_cell_wire[140];							inform_R[142][4] = r_cell_wire[141];							inform_R[135][4] = r_cell_wire[142];							inform_R[143][4] = r_cell_wire[143];							inform_R[144][4] = r_cell_wire[144];							inform_R[152][4] = r_cell_wire[145];							inform_R[145][4] = r_cell_wire[146];							inform_R[153][4] = r_cell_wire[147];							inform_R[146][4] = r_cell_wire[148];							inform_R[154][4] = r_cell_wire[149];							inform_R[147][4] = r_cell_wire[150];							inform_R[155][4] = r_cell_wire[151];							inform_R[148][4] = r_cell_wire[152];							inform_R[156][4] = r_cell_wire[153];							inform_R[149][4] = r_cell_wire[154];							inform_R[157][4] = r_cell_wire[155];							inform_R[150][4] = r_cell_wire[156];							inform_R[158][4] = r_cell_wire[157];							inform_R[151][4] = r_cell_wire[158];							inform_R[159][4] = r_cell_wire[159];							inform_R[160][4] = r_cell_wire[160];							inform_R[168][4] = r_cell_wire[161];							inform_R[161][4] = r_cell_wire[162];							inform_R[169][4] = r_cell_wire[163];							inform_R[162][4] = r_cell_wire[164];							inform_R[170][4] = r_cell_wire[165];							inform_R[163][4] = r_cell_wire[166];							inform_R[171][4] = r_cell_wire[167];							inform_R[164][4] = r_cell_wire[168];							inform_R[172][4] = r_cell_wire[169];							inform_R[165][4] = r_cell_wire[170];							inform_R[173][4] = r_cell_wire[171];							inform_R[166][4] = r_cell_wire[172];							inform_R[174][4] = r_cell_wire[173];							inform_R[167][4] = r_cell_wire[174];							inform_R[175][4] = r_cell_wire[175];							inform_R[176][4] = r_cell_wire[176];							inform_R[184][4] = r_cell_wire[177];							inform_R[177][4] = r_cell_wire[178];							inform_R[185][4] = r_cell_wire[179];							inform_R[178][4] = r_cell_wire[180];							inform_R[186][4] = r_cell_wire[181];							inform_R[179][4] = r_cell_wire[182];							inform_R[187][4] = r_cell_wire[183];							inform_R[180][4] = r_cell_wire[184];							inform_R[188][4] = r_cell_wire[185];							inform_R[181][4] = r_cell_wire[186];							inform_R[189][4] = r_cell_wire[187];							inform_R[182][4] = r_cell_wire[188];							inform_R[190][4] = r_cell_wire[189];							inform_R[183][4] = r_cell_wire[190];							inform_R[191][4] = r_cell_wire[191];							inform_R[192][4] = r_cell_wire[192];							inform_R[200][4] = r_cell_wire[193];							inform_R[193][4] = r_cell_wire[194];							inform_R[201][4] = r_cell_wire[195];							inform_R[194][4] = r_cell_wire[196];							inform_R[202][4] = r_cell_wire[197];							inform_R[195][4] = r_cell_wire[198];							inform_R[203][4] = r_cell_wire[199];							inform_R[196][4] = r_cell_wire[200];							inform_R[204][4] = r_cell_wire[201];							inform_R[197][4] = r_cell_wire[202];							inform_R[205][4] = r_cell_wire[203];							inform_R[198][4] = r_cell_wire[204];							inform_R[206][4] = r_cell_wire[205];							inform_R[199][4] = r_cell_wire[206];							inform_R[207][4] = r_cell_wire[207];							inform_R[208][4] = r_cell_wire[208];							inform_R[216][4] = r_cell_wire[209];							inform_R[209][4] = r_cell_wire[210];							inform_R[217][4] = r_cell_wire[211];							inform_R[210][4] = r_cell_wire[212];							inform_R[218][4] = r_cell_wire[213];							inform_R[211][4] = r_cell_wire[214];							inform_R[219][4] = r_cell_wire[215];							inform_R[212][4] = r_cell_wire[216];							inform_R[220][4] = r_cell_wire[217];							inform_R[213][4] = r_cell_wire[218];							inform_R[221][4] = r_cell_wire[219];							inform_R[214][4] = r_cell_wire[220];							inform_R[222][4] = r_cell_wire[221];							inform_R[215][4] = r_cell_wire[222];							inform_R[223][4] = r_cell_wire[223];							inform_R[224][4] = r_cell_wire[224];							inform_R[232][4] = r_cell_wire[225];							inform_R[225][4] = r_cell_wire[226];							inform_R[233][4] = r_cell_wire[227];							inform_R[226][4] = r_cell_wire[228];							inform_R[234][4] = r_cell_wire[229];							inform_R[227][4] = r_cell_wire[230];							inform_R[235][4] = r_cell_wire[231];							inform_R[228][4] = r_cell_wire[232];							inform_R[236][4] = r_cell_wire[233];							inform_R[229][4] = r_cell_wire[234];							inform_R[237][4] = r_cell_wire[235];							inform_R[230][4] = r_cell_wire[236];							inform_R[238][4] = r_cell_wire[237];							inform_R[231][4] = r_cell_wire[238];							inform_R[239][4] = r_cell_wire[239];							inform_R[240][4] = r_cell_wire[240];							inform_R[248][4] = r_cell_wire[241];							inform_R[241][4] = r_cell_wire[242];							inform_R[249][4] = r_cell_wire[243];							inform_R[242][4] = r_cell_wire[244];							inform_R[250][4] = r_cell_wire[245];							inform_R[243][4] = r_cell_wire[246];							inform_R[251][4] = r_cell_wire[247];							inform_R[244][4] = r_cell_wire[248];							inform_R[252][4] = r_cell_wire[249];							inform_R[245][4] = r_cell_wire[250];							inform_R[253][4] = r_cell_wire[251];							inform_R[246][4] = r_cell_wire[252];							inform_R[254][4] = r_cell_wire[253];							inform_R[247][4] = r_cell_wire[254];							inform_R[255][4] = r_cell_wire[255];							inform_R[256][4] = r_cell_wire[256];							inform_R[264][4] = r_cell_wire[257];							inform_R[257][4] = r_cell_wire[258];							inform_R[265][4] = r_cell_wire[259];							inform_R[258][4] = r_cell_wire[260];							inform_R[266][4] = r_cell_wire[261];							inform_R[259][4] = r_cell_wire[262];							inform_R[267][4] = r_cell_wire[263];							inform_R[260][4] = r_cell_wire[264];							inform_R[268][4] = r_cell_wire[265];							inform_R[261][4] = r_cell_wire[266];							inform_R[269][4] = r_cell_wire[267];							inform_R[262][4] = r_cell_wire[268];							inform_R[270][4] = r_cell_wire[269];							inform_R[263][4] = r_cell_wire[270];							inform_R[271][4] = r_cell_wire[271];							inform_R[272][4] = r_cell_wire[272];							inform_R[280][4] = r_cell_wire[273];							inform_R[273][4] = r_cell_wire[274];							inform_R[281][4] = r_cell_wire[275];							inform_R[274][4] = r_cell_wire[276];							inform_R[282][4] = r_cell_wire[277];							inform_R[275][4] = r_cell_wire[278];							inform_R[283][4] = r_cell_wire[279];							inform_R[276][4] = r_cell_wire[280];							inform_R[284][4] = r_cell_wire[281];							inform_R[277][4] = r_cell_wire[282];							inform_R[285][4] = r_cell_wire[283];							inform_R[278][4] = r_cell_wire[284];							inform_R[286][4] = r_cell_wire[285];							inform_R[279][4] = r_cell_wire[286];							inform_R[287][4] = r_cell_wire[287];							inform_R[288][4] = r_cell_wire[288];							inform_R[296][4] = r_cell_wire[289];							inform_R[289][4] = r_cell_wire[290];							inform_R[297][4] = r_cell_wire[291];							inform_R[290][4] = r_cell_wire[292];							inform_R[298][4] = r_cell_wire[293];							inform_R[291][4] = r_cell_wire[294];							inform_R[299][4] = r_cell_wire[295];							inform_R[292][4] = r_cell_wire[296];							inform_R[300][4] = r_cell_wire[297];							inform_R[293][4] = r_cell_wire[298];							inform_R[301][4] = r_cell_wire[299];							inform_R[294][4] = r_cell_wire[300];							inform_R[302][4] = r_cell_wire[301];							inform_R[295][4] = r_cell_wire[302];							inform_R[303][4] = r_cell_wire[303];							inform_R[304][4] = r_cell_wire[304];							inform_R[312][4] = r_cell_wire[305];							inform_R[305][4] = r_cell_wire[306];							inform_R[313][4] = r_cell_wire[307];							inform_R[306][4] = r_cell_wire[308];							inform_R[314][4] = r_cell_wire[309];							inform_R[307][4] = r_cell_wire[310];							inform_R[315][4] = r_cell_wire[311];							inform_R[308][4] = r_cell_wire[312];							inform_R[316][4] = r_cell_wire[313];							inform_R[309][4] = r_cell_wire[314];							inform_R[317][4] = r_cell_wire[315];							inform_R[310][4] = r_cell_wire[316];							inform_R[318][4] = r_cell_wire[317];							inform_R[311][4] = r_cell_wire[318];							inform_R[319][4] = r_cell_wire[319];							inform_R[320][4] = r_cell_wire[320];							inform_R[328][4] = r_cell_wire[321];							inform_R[321][4] = r_cell_wire[322];							inform_R[329][4] = r_cell_wire[323];							inform_R[322][4] = r_cell_wire[324];							inform_R[330][4] = r_cell_wire[325];							inform_R[323][4] = r_cell_wire[326];							inform_R[331][4] = r_cell_wire[327];							inform_R[324][4] = r_cell_wire[328];							inform_R[332][4] = r_cell_wire[329];							inform_R[325][4] = r_cell_wire[330];							inform_R[333][4] = r_cell_wire[331];							inform_R[326][4] = r_cell_wire[332];							inform_R[334][4] = r_cell_wire[333];							inform_R[327][4] = r_cell_wire[334];							inform_R[335][4] = r_cell_wire[335];							inform_R[336][4] = r_cell_wire[336];							inform_R[344][4] = r_cell_wire[337];							inform_R[337][4] = r_cell_wire[338];							inform_R[345][4] = r_cell_wire[339];							inform_R[338][4] = r_cell_wire[340];							inform_R[346][4] = r_cell_wire[341];							inform_R[339][4] = r_cell_wire[342];							inform_R[347][4] = r_cell_wire[343];							inform_R[340][4] = r_cell_wire[344];							inform_R[348][4] = r_cell_wire[345];							inform_R[341][4] = r_cell_wire[346];							inform_R[349][4] = r_cell_wire[347];							inform_R[342][4] = r_cell_wire[348];							inform_R[350][4] = r_cell_wire[349];							inform_R[343][4] = r_cell_wire[350];							inform_R[351][4] = r_cell_wire[351];							inform_R[352][4] = r_cell_wire[352];							inform_R[360][4] = r_cell_wire[353];							inform_R[353][4] = r_cell_wire[354];							inform_R[361][4] = r_cell_wire[355];							inform_R[354][4] = r_cell_wire[356];							inform_R[362][4] = r_cell_wire[357];							inform_R[355][4] = r_cell_wire[358];							inform_R[363][4] = r_cell_wire[359];							inform_R[356][4] = r_cell_wire[360];							inform_R[364][4] = r_cell_wire[361];							inform_R[357][4] = r_cell_wire[362];							inform_R[365][4] = r_cell_wire[363];							inform_R[358][4] = r_cell_wire[364];							inform_R[366][4] = r_cell_wire[365];							inform_R[359][4] = r_cell_wire[366];							inform_R[367][4] = r_cell_wire[367];							inform_R[368][4] = r_cell_wire[368];							inform_R[376][4] = r_cell_wire[369];							inform_R[369][4] = r_cell_wire[370];							inform_R[377][4] = r_cell_wire[371];							inform_R[370][4] = r_cell_wire[372];							inform_R[378][4] = r_cell_wire[373];							inform_R[371][4] = r_cell_wire[374];							inform_R[379][4] = r_cell_wire[375];							inform_R[372][4] = r_cell_wire[376];							inform_R[380][4] = r_cell_wire[377];							inform_R[373][4] = r_cell_wire[378];							inform_R[381][4] = r_cell_wire[379];							inform_R[374][4] = r_cell_wire[380];							inform_R[382][4] = r_cell_wire[381];							inform_R[375][4] = r_cell_wire[382];							inform_R[383][4] = r_cell_wire[383];							inform_R[384][4] = r_cell_wire[384];							inform_R[392][4] = r_cell_wire[385];							inform_R[385][4] = r_cell_wire[386];							inform_R[393][4] = r_cell_wire[387];							inform_R[386][4] = r_cell_wire[388];							inform_R[394][4] = r_cell_wire[389];							inform_R[387][4] = r_cell_wire[390];							inform_R[395][4] = r_cell_wire[391];							inform_R[388][4] = r_cell_wire[392];							inform_R[396][4] = r_cell_wire[393];							inform_R[389][4] = r_cell_wire[394];							inform_R[397][4] = r_cell_wire[395];							inform_R[390][4] = r_cell_wire[396];							inform_R[398][4] = r_cell_wire[397];							inform_R[391][4] = r_cell_wire[398];							inform_R[399][4] = r_cell_wire[399];							inform_R[400][4] = r_cell_wire[400];							inform_R[408][4] = r_cell_wire[401];							inform_R[401][4] = r_cell_wire[402];							inform_R[409][4] = r_cell_wire[403];							inform_R[402][4] = r_cell_wire[404];							inform_R[410][4] = r_cell_wire[405];							inform_R[403][4] = r_cell_wire[406];							inform_R[411][4] = r_cell_wire[407];							inform_R[404][4] = r_cell_wire[408];							inform_R[412][4] = r_cell_wire[409];							inform_R[405][4] = r_cell_wire[410];							inform_R[413][4] = r_cell_wire[411];							inform_R[406][4] = r_cell_wire[412];							inform_R[414][4] = r_cell_wire[413];							inform_R[407][4] = r_cell_wire[414];							inform_R[415][4] = r_cell_wire[415];							inform_R[416][4] = r_cell_wire[416];							inform_R[424][4] = r_cell_wire[417];							inform_R[417][4] = r_cell_wire[418];							inform_R[425][4] = r_cell_wire[419];							inform_R[418][4] = r_cell_wire[420];							inform_R[426][4] = r_cell_wire[421];							inform_R[419][4] = r_cell_wire[422];							inform_R[427][4] = r_cell_wire[423];							inform_R[420][4] = r_cell_wire[424];							inform_R[428][4] = r_cell_wire[425];							inform_R[421][4] = r_cell_wire[426];							inform_R[429][4] = r_cell_wire[427];							inform_R[422][4] = r_cell_wire[428];							inform_R[430][4] = r_cell_wire[429];							inform_R[423][4] = r_cell_wire[430];							inform_R[431][4] = r_cell_wire[431];							inform_R[432][4] = r_cell_wire[432];							inform_R[440][4] = r_cell_wire[433];							inform_R[433][4] = r_cell_wire[434];							inform_R[441][4] = r_cell_wire[435];							inform_R[434][4] = r_cell_wire[436];							inform_R[442][4] = r_cell_wire[437];							inform_R[435][4] = r_cell_wire[438];							inform_R[443][4] = r_cell_wire[439];							inform_R[436][4] = r_cell_wire[440];							inform_R[444][4] = r_cell_wire[441];							inform_R[437][4] = r_cell_wire[442];							inform_R[445][4] = r_cell_wire[443];							inform_R[438][4] = r_cell_wire[444];							inform_R[446][4] = r_cell_wire[445];							inform_R[439][4] = r_cell_wire[446];							inform_R[447][4] = r_cell_wire[447];							inform_R[448][4] = r_cell_wire[448];							inform_R[456][4] = r_cell_wire[449];							inform_R[449][4] = r_cell_wire[450];							inform_R[457][4] = r_cell_wire[451];							inform_R[450][4] = r_cell_wire[452];							inform_R[458][4] = r_cell_wire[453];							inform_R[451][4] = r_cell_wire[454];							inform_R[459][4] = r_cell_wire[455];							inform_R[452][4] = r_cell_wire[456];							inform_R[460][4] = r_cell_wire[457];							inform_R[453][4] = r_cell_wire[458];							inform_R[461][4] = r_cell_wire[459];							inform_R[454][4] = r_cell_wire[460];							inform_R[462][4] = r_cell_wire[461];							inform_R[455][4] = r_cell_wire[462];							inform_R[463][4] = r_cell_wire[463];							inform_R[464][4] = r_cell_wire[464];							inform_R[472][4] = r_cell_wire[465];							inform_R[465][4] = r_cell_wire[466];							inform_R[473][4] = r_cell_wire[467];							inform_R[466][4] = r_cell_wire[468];							inform_R[474][4] = r_cell_wire[469];							inform_R[467][4] = r_cell_wire[470];							inform_R[475][4] = r_cell_wire[471];							inform_R[468][4] = r_cell_wire[472];							inform_R[476][4] = r_cell_wire[473];							inform_R[469][4] = r_cell_wire[474];							inform_R[477][4] = r_cell_wire[475];							inform_R[470][4] = r_cell_wire[476];							inform_R[478][4] = r_cell_wire[477];							inform_R[471][4] = r_cell_wire[478];							inform_R[479][4] = r_cell_wire[479];							inform_R[480][4] = r_cell_wire[480];							inform_R[488][4] = r_cell_wire[481];							inform_R[481][4] = r_cell_wire[482];							inform_R[489][4] = r_cell_wire[483];							inform_R[482][4] = r_cell_wire[484];							inform_R[490][4] = r_cell_wire[485];							inform_R[483][4] = r_cell_wire[486];							inform_R[491][4] = r_cell_wire[487];							inform_R[484][4] = r_cell_wire[488];							inform_R[492][4] = r_cell_wire[489];							inform_R[485][4] = r_cell_wire[490];							inform_R[493][4] = r_cell_wire[491];							inform_R[486][4] = r_cell_wire[492];							inform_R[494][4] = r_cell_wire[493];							inform_R[487][4] = r_cell_wire[494];							inform_R[495][4] = r_cell_wire[495];							inform_R[496][4] = r_cell_wire[496];							inform_R[504][4] = r_cell_wire[497];							inform_R[497][4] = r_cell_wire[498];							inform_R[505][4] = r_cell_wire[499];							inform_R[498][4] = r_cell_wire[500];							inform_R[506][4] = r_cell_wire[501];							inform_R[499][4] = r_cell_wire[502];							inform_R[507][4] = r_cell_wire[503];							inform_R[500][4] = r_cell_wire[504];							inform_R[508][4] = r_cell_wire[505];							inform_R[501][4] = r_cell_wire[506];							inform_R[509][4] = r_cell_wire[507];							inform_R[502][4] = r_cell_wire[508];							inform_R[510][4] = r_cell_wire[509];							inform_R[503][4] = r_cell_wire[510];							inform_R[511][4] = r_cell_wire[511];							inform_R[512][4] = r_cell_wire[512];							inform_R[520][4] = r_cell_wire[513];							inform_R[513][4] = r_cell_wire[514];							inform_R[521][4] = r_cell_wire[515];							inform_R[514][4] = r_cell_wire[516];							inform_R[522][4] = r_cell_wire[517];							inform_R[515][4] = r_cell_wire[518];							inform_R[523][4] = r_cell_wire[519];							inform_R[516][4] = r_cell_wire[520];							inform_R[524][4] = r_cell_wire[521];							inform_R[517][4] = r_cell_wire[522];							inform_R[525][4] = r_cell_wire[523];							inform_R[518][4] = r_cell_wire[524];							inform_R[526][4] = r_cell_wire[525];							inform_R[519][4] = r_cell_wire[526];							inform_R[527][4] = r_cell_wire[527];							inform_R[528][4] = r_cell_wire[528];							inform_R[536][4] = r_cell_wire[529];							inform_R[529][4] = r_cell_wire[530];							inform_R[537][4] = r_cell_wire[531];							inform_R[530][4] = r_cell_wire[532];							inform_R[538][4] = r_cell_wire[533];							inform_R[531][4] = r_cell_wire[534];							inform_R[539][4] = r_cell_wire[535];							inform_R[532][4] = r_cell_wire[536];							inform_R[540][4] = r_cell_wire[537];							inform_R[533][4] = r_cell_wire[538];							inform_R[541][4] = r_cell_wire[539];							inform_R[534][4] = r_cell_wire[540];							inform_R[542][4] = r_cell_wire[541];							inform_R[535][4] = r_cell_wire[542];							inform_R[543][4] = r_cell_wire[543];							inform_R[544][4] = r_cell_wire[544];							inform_R[552][4] = r_cell_wire[545];							inform_R[545][4] = r_cell_wire[546];							inform_R[553][4] = r_cell_wire[547];							inform_R[546][4] = r_cell_wire[548];							inform_R[554][4] = r_cell_wire[549];							inform_R[547][4] = r_cell_wire[550];							inform_R[555][4] = r_cell_wire[551];							inform_R[548][4] = r_cell_wire[552];							inform_R[556][4] = r_cell_wire[553];							inform_R[549][4] = r_cell_wire[554];							inform_R[557][4] = r_cell_wire[555];							inform_R[550][4] = r_cell_wire[556];							inform_R[558][4] = r_cell_wire[557];							inform_R[551][4] = r_cell_wire[558];							inform_R[559][4] = r_cell_wire[559];							inform_R[560][4] = r_cell_wire[560];							inform_R[568][4] = r_cell_wire[561];							inform_R[561][4] = r_cell_wire[562];							inform_R[569][4] = r_cell_wire[563];							inform_R[562][4] = r_cell_wire[564];							inform_R[570][4] = r_cell_wire[565];							inform_R[563][4] = r_cell_wire[566];							inform_R[571][4] = r_cell_wire[567];							inform_R[564][4] = r_cell_wire[568];							inform_R[572][4] = r_cell_wire[569];							inform_R[565][4] = r_cell_wire[570];							inform_R[573][4] = r_cell_wire[571];							inform_R[566][4] = r_cell_wire[572];							inform_R[574][4] = r_cell_wire[573];							inform_R[567][4] = r_cell_wire[574];							inform_R[575][4] = r_cell_wire[575];							inform_R[576][4] = r_cell_wire[576];							inform_R[584][4] = r_cell_wire[577];							inform_R[577][4] = r_cell_wire[578];							inform_R[585][4] = r_cell_wire[579];							inform_R[578][4] = r_cell_wire[580];							inform_R[586][4] = r_cell_wire[581];							inform_R[579][4] = r_cell_wire[582];							inform_R[587][4] = r_cell_wire[583];							inform_R[580][4] = r_cell_wire[584];							inform_R[588][4] = r_cell_wire[585];							inform_R[581][4] = r_cell_wire[586];							inform_R[589][4] = r_cell_wire[587];							inform_R[582][4] = r_cell_wire[588];							inform_R[590][4] = r_cell_wire[589];							inform_R[583][4] = r_cell_wire[590];							inform_R[591][4] = r_cell_wire[591];							inform_R[592][4] = r_cell_wire[592];							inform_R[600][4] = r_cell_wire[593];							inform_R[593][4] = r_cell_wire[594];							inform_R[601][4] = r_cell_wire[595];							inform_R[594][4] = r_cell_wire[596];							inform_R[602][4] = r_cell_wire[597];							inform_R[595][4] = r_cell_wire[598];							inform_R[603][4] = r_cell_wire[599];							inform_R[596][4] = r_cell_wire[600];							inform_R[604][4] = r_cell_wire[601];							inform_R[597][4] = r_cell_wire[602];							inform_R[605][4] = r_cell_wire[603];							inform_R[598][4] = r_cell_wire[604];							inform_R[606][4] = r_cell_wire[605];							inform_R[599][4] = r_cell_wire[606];							inform_R[607][4] = r_cell_wire[607];							inform_R[608][4] = r_cell_wire[608];							inform_R[616][4] = r_cell_wire[609];							inform_R[609][4] = r_cell_wire[610];							inform_R[617][4] = r_cell_wire[611];							inform_R[610][4] = r_cell_wire[612];							inform_R[618][4] = r_cell_wire[613];							inform_R[611][4] = r_cell_wire[614];							inform_R[619][4] = r_cell_wire[615];							inform_R[612][4] = r_cell_wire[616];							inform_R[620][4] = r_cell_wire[617];							inform_R[613][4] = r_cell_wire[618];							inform_R[621][4] = r_cell_wire[619];							inform_R[614][4] = r_cell_wire[620];							inform_R[622][4] = r_cell_wire[621];							inform_R[615][4] = r_cell_wire[622];							inform_R[623][4] = r_cell_wire[623];							inform_R[624][4] = r_cell_wire[624];							inform_R[632][4] = r_cell_wire[625];							inform_R[625][4] = r_cell_wire[626];							inform_R[633][4] = r_cell_wire[627];							inform_R[626][4] = r_cell_wire[628];							inform_R[634][4] = r_cell_wire[629];							inform_R[627][4] = r_cell_wire[630];							inform_R[635][4] = r_cell_wire[631];							inform_R[628][4] = r_cell_wire[632];							inform_R[636][4] = r_cell_wire[633];							inform_R[629][4] = r_cell_wire[634];							inform_R[637][4] = r_cell_wire[635];							inform_R[630][4] = r_cell_wire[636];							inform_R[638][4] = r_cell_wire[637];							inform_R[631][4] = r_cell_wire[638];							inform_R[639][4] = r_cell_wire[639];							inform_R[640][4] = r_cell_wire[640];							inform_R[648][4] = r_cell_wire[641];							inform_R[641][4] = r_cell_wire[642];							inform_R[649][4] = r_cell_wire[643];							inform_R[642][4] = r_cell_wire[644];							inform_R[650][4] = r_cell_wire[645];							inform_R[643][4] = r_cell_wire[646];							inform_R[651][4] = r_cell_wire[647];							inform_R[644][4] = r_cell_wire[648];							inform_R[652][4] = r_cell_wire[649];							inform_R[645][4] = r_cell_wire[650];							inform_R[653][4] = r_cell_wire[651];							inform_R[646][4] = r_cell_wire[652];							inform_R[654][4] = r_cell_wire[653];							inform_R[647][4] = r_cell_wire[654];							inform_R[655][4] = r_cell_wire[655];							inform_R[656][4] = r_cell_wire[656];							inform_R[664][4] = r_cell_wire[657];							inform_R[657][4] = r_cell_wire[658];							inform_R[665][4] = r_cell_wire[659];							inform_R[658][4] = r_cell_wire[660];							inform_R[666][4] = r_cell_wire[661];							inform_R[659][4] = r_cell_wire[662];							inform_R[667][4] = r_cell_wire[663];							inform_R[660][4] = r_cell_wire[664];							inform_R[668][4] = r_cell_wire[665];							inform_R[661][4] = r_cell_wire[666];							inform_R[669][4] = r_cell_wire[667];							inform_R[662][4] = r_cell_wire[668];							inform_R[670][4] = r_cell_wire[669];							inform_R[663][4] = r_cell_wire[670];							inform_R[671][4] = r_cell_wire[671];							inform_R[672][4] = r_cell_wire[672];							inform_R[680][4] = r_cell_wire[673];							inform_R[673][4] = r_cell_wire[674];							inform_R[681][4] = r_cell_wire[675];							inform_R[674][4] = r_cell_wire[676];							inform_R[682][4] = r_cell_wire[677];							inform_R[675][4] = r_cell_wire[678];							inform_R[683][4] = r_cell_wire[679];							inform_R[676][4] = r_cell_wire[680];							inform_R[684][4] = r_cell_wire[681];							inform_R[677][4] = r_cell_wire[682];							inform_R[685][4] = r_cell_wire[683];							inform_R[678][4] = r_cell_wire[684];							inform_R[686][4] = r_cell_wire[685];							inform_R[679][4] = r_cell_wire[686];							inform_R[687][4] = r_cell_wire[687];							inform_R[688][4] = r_cell_wire[688];							inform_R[696][4] = r_cell_wire[689];							inform_R[689][4] = r_cell_wire[690];							inform_R[697][4] = r_cell_wire[691];							inform_R[690][4] = r_cell_wire[692];							inform_R[698][4] = r_cell_wire[693];							inform_R[691][4] = r_cell_wire[694];							inform_R[699][4] = r_cell_wire[695];							inform_R[692][4] = r_cell_wire[696];							inform_R[700][4] = r_cell_wire[697];							inform_R[693][4] = r_cell_wire[698];							inform_R[701][4] = r_cell_wire[699];							inform_R[694][4] = r_cell_wire[700];							inform_R[702][4] = r_cell_wire[701];							inform_R[695][4] = r_cell_wire[702];							inform_R[703][4] = r_cell_wire[703];							inform_R[704][4] = r_cell_wire[704];							inform_R[712][4] = r_cell_wire[705];							inform_R[705][4] = r_cell_wire[706];							inform_R[713][4] = r_cell_wire[707];							inform_R[706][4] = r_cell_wire[708];							inform_R[714][4] = r_cell_wire[709];							inform_R[707][4] = r_cell_wire[710];							inform_R[715][4] = r_cell_wire[711];							inform_R[708][4] = r_cell_wire[712];							inform_R[716][4] = r_cell_wire[713];							inform_R[709][4] = r_cell_wire[714];							inform_R[717][4] = r_cell_wire[715];							inform_R[710][4] = r_cell_wire[716];							inform_R[718][4] = r_cell_wire[717];							inform_R[711][4] = r_cell_wire[718];							inform_R[719][4] = r_cell_wire[719];							inform_R[720][4] = r_cell_wire[720];							inform_R[728][4] = r_cell_wire[721];							inform_R[721][4] = r_cell_wire[722];							inform_R[729][4] = r_cell_wire[723];							inform_R[722][4] = r_cell_wire[724];							inform_R[730][4] = r_cell_wire[725];							inform_R[723][4] = r_cell_wire[726];							inform_R[731][4] = r_cell_wire[727];							inform_R[724][4] = r_cell_wire[728];							inform_R[732][4] = r_cell_wire[729];							inform_R[725][4] = r_cell_wire[730];							inform_R[733][4] = r_cell_wire[731];							inform_R[726][4] = r_cell_wire[732];							inform_R[734][4] = r_cell_wire[733];							inform_R[727][4] = r_cell_wire[734];							inform_R[735][4] = r_cell_wire[735];							inform_R[736][4] = r_cell_wire[736];							inform_R[744][4] = r_cell_wire[737];							inform_R[737][4] = r_cell_wire[738];							inform_R[745][4] = r_cell_wire[739];							inform_R[738][4] = r_cell_wire[740];							inform_R[746][4] = r_cell_wire[741];							inform_R[739][4] = r_cell_wire[742];							inform_R[747][4] = r_cell_wire[743];							inform_R[740][4] = r_cell_wire[744];							inform_R[748][4] = r_cell_wire[745];							inform_R[741][4] = r_cell_wire[746];							inform_R[749][4] = r_cell_wire[747];							inform_R[742][4] = r_cell_wire[748];							inform_R[750][4] = r_cell_wire[749];							inform_R[743][4] = r_cell_wire[750];							inform_R[751][4] = r_cell_wire[751];							inform_R[752][4] = r_cell_wire[752];							inform_R[760][4] = r_cell_wire[753];							inform_R[753][4] = r_cell_wire[754];							inform_R[761][4] = r_cell_wire[755];							inform_R[754][4] = r_cell_wire[756];							inform_R[762][4] = r_cell_wire[757];							inform_R[755][4] = r_cell_wire[758];							inform_R[763][4] = r_cell_wire[759];							inform_R[756][4] = r_cell_wire[760];							inform_R[764][4] = r_cell_wire[761];							inform_R[757][4] = r_cell_wire[762];							inform_R[765][4] = r_cell_wire[763];							inform_R[758][4] = r_cell_wire[764];							inform_R[766][4] = r_cell_wire[765];							inform_R[759][4] = r_cell_wire[766];							inform_R[767][4] = r_cell_wire[767];							inform_R[768][4] = r_cell_wire[768];							inform_R[776][4] = r_cell_wire[769];							inform_R[769][4] = r_cell_wire[770];							inform_R[777][4] = r_cell_wire[771];							inform_R[770][4] = r_cell_wire[772];							inform_R[778][4] = r_cell_wire[773];							inform_R[771][4] = r_cell_wire[774];							inform_R[779][4] = r_cell_wire[775];							inform_R[772][4] = r_cell_wire[776];							inform_R[780][4] = r_cell_wire[777];							inform_R[773][4] = r_cell_wire[778];							inform_R[781][4] = r_cell_wire[779];							inform_R[774][4] = r_cell_wire[780];							inform_R[782][4] = r_cell_wire[781];							inform_R[775][4] = r_cell_wire[782];							inform_R[783][4] = r_cell_wire[783];							inform_R[784][4] = r_cell_wire[784];							inform_R[792][4] = r_cell_wire[785];							inform_R[785][4] = r_cell_wire[786];							inform_R[793][4] = r_cell_wire[787];							inform_R[786][4] = r_cell_wire[788];							inform_R[794][4] = r_cell_wire[789];							inform_R[787][4] = r_cell_wire[790];							inform_R[795][4] = r_cell_wire[791];							inform_R[788][4] = r_cell_wire[792];							inform_R[796][4] = r_cell_wire[793];							inform_R[789][4] = r_cell_wire[794];							inform_R[797][4] = r_cell_wire[795];							inform_R[790][4] = r_cell_wire[796];							inform_R[798][4] = r_cell_wire[797];							inform_R[791][4] = r_cell_wire[798];							inform_R[799][4] = r_cell_wire[799];							inform_R[800][4] = r_cell_wire[800];							inform_R[808][4] = r_cell_wire[801];							inform_R[801][4] = r_cell_wire[802];							inform_R[809][4] = r_cell_wire[803];							inform_R[802][4] = r_cell_wire[804];							inform_R[810][4] = r_cell_wire[805];							inform_R[803][4] = r_cell_wire[806];							inform_R[811][4] = r_cell_wire[807];							inform_R[804][4] = r_cell_wire[808];							inform_R[812][4] = r_cell_wire[809];							inform_R[805][4] = r_cell_wire[810];							inform_R[813][4] = r_cell_wire[811];							inform_R[806][4] = r_cell_wire[812];							inform_R[814][4] = r_cell_wire[813];							inform_R[807][4] = r_cell_wire[814];							inform_R[815][4] = r_cell_wire[815];							inform_R[816][4] = r_cell_wire[816];							inform_R[824][4] = r_cell_wire[817];							inform_R[817][4] = r_cell_wire[818];							inform_R[825][4] = r_cell_wire[819];							inform_R[818][4] = r_cell_wire[820];							inform_R[826][4] = r_cell_wire[821];							inform_R[819][4] = r_cell_wire[822];							inform_R[827][4] = r_cell_wire[823];							inform_R[820][4] = r_cell_wire[824];							inform_R[828][4] = r_cell_wire[825];							inform_R[821][4] = r_cell_wire[826];							inform_R[829][4] = r_cell_wire[827];							inform_R[822][4] = r_cell_wire[828];							inform_R[830][4] = r_cell_wire[829];							inform_R[823][4] = r_cell_wire[830];							inform_R[831][4] = r_cell_wire[831];							inform_R[832][4] = r_cell_wire[832];							inform_R[840][4] = r_cell_wire[833];							inform_R[833][4] = r_cell_wire[834];							inform_R[841][4] = r_cell_wire[835];							inform_R[834][4] = r_cell_wire[836];							inform_R[842][4] = r_cell_wire[837];							inform_R[835][4] = r_cell_wire[838];							inform_R[843][4] = r_cell_wire[839];							inform_R[836][4] = r_cell_wire[840];							inform_R[844][4] = r_cell_wire[841];							inform_R[837][4] = r_cell_wire[842];							inform_R[845][4] = r_cell_wire[843];							inform_R[838][4] = r_cell_wire[844];							inform_R[846][4] = r_cell_wire[845];							inform_R[839][4] = r_cell_wire[846];							inform_R[847][4] = r_cell_wire[847];							inform_R[848][4] = r_cell_wire[848];							inform_R[856][4] = r_cell_wire[849];							inform_R[849][4] = r_cell_wire[850];							inform_R[857][4] = r_cell_wire[851];							inform_R[850][4] = r_cell_wire[852];							inform_R[858][4] = r_cell_wire[853];							inform_R[851][4] = r_cell_wire[854];							inform_R[859][4] = r_cell_wire[855];							inform_R[852][4] = r_cell_wire[856];							inform_R[860][4] = r_cell_wire[857];							inform_R[853][4] = r_cell_wire[858];							inform_R[861][4] = r_cell_wire[859];							inform_R[854][4] = r_cell_wire[860];							inform_R[862][4] = r_cell_wire[861];							inform_R[855][4] = r_cell_wire[862];							inform_R[863][4] = r_cell_wire[863];							inform_R[864][4] = r_cell_wire[864];							inform_R[872][4] = r_cell_wire[865];							inform_R[865][4] = r_cell_wire[866];							inform_R[873][4] = r_cell_wire[867];							inform_R[866][4] = r_cell_wire[868];							inform_R[874][4] = r_cell_wire[869];							inform_R[867][4] = r_cell_wire[870];							inform_R[875][4] = r_cell_wire[871];							inform_R[868][4] = r_cell_wire[872];							inform_R[876][4] = r_cell_wire[873];							inform_R[869][4] = r_cell_wire[874];							inform_R[877][4] = r_cell_wire[875];							inform_R[870][4] = r_cell_wire[876];							inform_R[878][4] = r_cell_wire[877];							inform_R[871][4] = r_cell_wire[878];							inform_R[879][4] = r_cell_wire[879];							inform_R[880][4] = r_cell_wire[880];							inform_R[888][4] = r_cell_wire[881];							inform_R[881][4] = r_cell_wire[882];							inform_R[889][4] = r_cell_wire[883];							inform_R[882][4] = r_cell_wire[884];							inform_R[890][4] = r_cell_wire[885];							inform_R[883][4] = r_cell_wire[886];							inform_R[891][4] = r_cell_wire[887];							inform_R[884][4] = r_cell_wire[888];							inform_R[892][4] = r_cell_wire[889];							inform_R[885][4] = r_cell_wire[890];							inform_R[893][4] = r_cell_wire[891];							inform_R[886][4] = r_cell_wire[892];							inform_R[894][4] = r_cell_wire[893];							inform_R[887][4] = r_cell_wire[894];							inform_R[895][4] = r_cell_wire[895];							inform_R[896][4] = r_cell_wire[896];							inform_R[904][4] = r_cell_wire[897];							inform_R[897][4] = r_cell_wire[898];							inform_R[905][4] = r_cell_wire[899];							inform_R[898][4] = r_cell_wire[900];							inform_R[906][4] = r_cell_wire[901];							inform_R[899][4] = r_cell_wire[902];							inform_R[907][4] = r_cell_wire[903];							inform_R[900][4] = r_cell_wire[904];							inform_R[908][4] = r_cell_wire[905];							inform_R[901][4] = r_cell_wire[906];							inform_R[909][4] = r_cell_wire[907];							inform_R[902][4] = r_cell_wire[908];							inform_R[910][4] = r_cell_wire[909];							inform_R[903][4] = r_cell_wire[910];							inform_R[911][4] = r_cell_wire[911];							inform_R[912][4] = r_cell_wire[912];							inform_R[920][4] = r_cell_wire[913];							inform_R[913][4] = r_cell_wire[914];							inform_R[921][4] = r_cell_wire[915];							inform_R[914][4] = r_cell_wire[916];							inform_R[922][4] = r_cell_wire[917];							inform_R[915][4] = r_cell_wire[918];							inform_R[923][4] = r_cell_wire[919];							inform_R[916][4] = r_cell_wire[920];							inform_R[924][4] = r_cell_wire[921];							inform_R[917][4] = r_cell_wire[922];							inform_R[925][4] = r_cell_wire[923];							inform_R[918][4] = r_cell_wire[924];							inform_R[926][4] = r_cell_wire[925];							inform_R[919][4] = r_cell_wire[926];							inform_R[927][4] = r_cell_wire[927];							inform_R[928][4] = r_cell_wire[928];							inform_R[936][4] = r_cell_wire[929];							inform_R[929][4] = r_cell_wire[930];							inform_R[937][4] = r_cell_wire[931];							inform_R[930][4] = r_cell_wire[932];							inform_R[938][4] = r_cell_wire[933];							inform_R[931][4] = r_cell_wire[934];							inform_R[939][4] = r_cell_wire[935];							inform_R[932][4] = r_cell_wire[936];							inform_R[940][4] = r_cell_wire[937];							inform_R[933][4] = r_cell_wire[938];							inform_R[941][4] = r_cell_wire[939];							inform_R[934][4] = r_cell_wire[940];							inform_R[942][4] = r_cell_wire[941];							inform_R[935][4] = r_cell_wire[942];							inform_R[943][4] = r_cell_wire[943];							inform_R[944][4] = r_cell_wire[944];							inform_R[952][4] = r_cell_wire[945];							inform_R[945][4] = r_cell_wire[946];							inform_R[953][4] = r_cell_wire[947];							inform_R[946][4] = r_cell_wire[948];							inform_R[954][4] = r_cell_wire[949];							inform_R[947][4] = r_cell_wire[950];							inform_R[955][4] = r_cell_wire[951];							inform_R[948][4] = r_cell_wire[952];							inform_R[956][4] = r_cell_wire[953];							inform_R[949][4] = r_cell_wire[954];							inform_R[957][4] = r_cell_wire[955];							inform_R[950][4] = r_cell_wire[956];							inform_R[958][4] = r_cell_wire[957];							inform_R[951][4] = r_cell_wire[958];							inform_R[959][4] = r_cell_wire[959];							inform_R[960][4] = r_cell_wire[960];							inform_R[968][4] = r_cell_wire[961];							inform_R[961][4] = r_cell_wire[962];							inform_R[969][4] = r_cell_wire[963];							inform_R[962][4] = r_cell_wire[964];							inform_R[970][4] = r_cell_wire[965];							inform_R[963][4] = r_cell_wire[966];							inform_R[971][4] = r_cell_wire[967];							inform_R[964][4] = r_cell_wire[968];							inform_R[972][4] = r_cell_wire[969];							inform_R[965][4] = r_cell_wire[970];							inform_R[973][4] = r_cell_wire[971];							inform_R[966][4] = r_cell_wire[972];							inform_R[974][4] = r_cell_wire[973];							inform_R[967][4] = r_cell_wire[974];							inform_R[975][4] = r_cell_wire[975];							inform_R[976][4] = r_cell_wire[976];							inform_R[984][4] = r_cell_wire[977];							inform_R[977][4] = r_cell_wire[978];							inform_R[985][4] = r_cell_wire[979];							inform_R[978][4] = r_cell_wire[980];							inform_R[986][4] = r_cell_wire[981];							inform_R[979][4] = r_cell_wire[982];							inform_R[987][4] = r_cell_wire[983];							inform_R[980][4] = r_cell_wire[984];							inform_R[988][4] = r_cell_wire[985];							inform_R[981][4] = r_cell_wire[986];							inform_R[989][4] = r_cell_wire[987];							inform_R[982][4] = r_cell_wire[988];							inform_R[990][4] = r_cell_wire[989];							inform_R[983][4] = r_cell_wire[990];							inform_R[991][4] = r_cell_wire[991];							inform_R[992][4] = r_cell_wire[992];							inform_R[1000][4] = r_cell_wire[993];							inform_R[993][4] = r_cell_wire[994];							inform_R[1001][4] = r_cell_wire[995];							inform_R[994][4] = r_cell_wire[996];							inform_R[1002][4] = r_cell_wire[997];							inform_R[995][4] = r_cell_wire[998];							inform_R[1003][4] = r_cell_wire[999];							inform_R[996][4] = r_cell_wire[1000];							inform_R[1004][4] = r_cell_wire[1001];							inform_R[997][4] = r_cell_wire[1002];							inform_R[1005][4] = r_cell_wire[1003];							inform_R[998][4] = r_cell_wire[1004];							inform_R[1006][4] = r_cell_wire[1005];							inform_R[999][4] = r_cell_wire[1006];							inform_R[1007][4] = r_cell_wire[1007];							inform_R[1008][4] = r_cell_wire[1008];							inform_R[1016][4] = r_cell_wire[1009];							inform_R[1009][4] = r_cell_wire[1010];							inform_R[1017][4] = r_cell_wire[1011];							inform_R[1010][4] = r_cell_wire[1012];							inform_R[1018][4] = r_cell_wire[1013];							inform_R[1011][4] = r_cell_wire[1014];							inform_R[1019][4] = r_cell_wire[1015];							inform_R[1012][4] = r_cell_wire[1016];							inform_R[1020][4] = r_cell_wire[1017];							inform_R[1013][4] = r_cell_wire[1018];							inform_R[1021][4] = r_cell_wire[1019];							inform_R[1014][4] = r_cell_wire[1020];							inform_R[1022][4] = r_cell_wire[1021];							inform_R[1015][4] = r_cell_wire[1022];							inform_R[1023][4] = r_cell_wire[1023];							inform_L[0][3] = l_cell_wire[0];							inform_L[8][3] = l_cell_wire[1];							inform_L[1][3] = l_cell_wire[2];							inform_L[9][3] = l_cell_wire[3];							inform_L[2][3] = l_cell_wire[4];							inform_L[10][3] = l_cell_wire[5];							inform_L[3][3] = l_cell_wire[6];							inform_L[11][3] = l_cell_wire[7];							inform_L[4][3] = l_cell_wire[8];							inform_L[12][3] = l_cell_wire[9];							inform_L[5][3] = l_cell_wire[10];							inform_L[13][3] = l_cell_wire[11];							inform_L[6][3] = l_cell_wire[12];							inform_L[14][3] = l_cell_wire[13];							inform_L[7][3] = l_cell_wire[14];							inform_L[15][3] = l_cell_wire[15];							inform_L[16][3] = l_cell_wire[16];							inform_L[24][3] = l_cell_wire[17];							inform_L[17][3] = l_cell_wire[18];							inform_L[25][3] = l_cell_wire[19];							inform_L[18][3] = l_cell_wire[20];							inform_L[26][3] = l_cell_wire[21];							inform_L[19][3] = l_cell_wire[22];							inform_L[27][3] = l_cell_wire[23];							inform_L[20][3] = l_cell_wire[24];							inform_L[28][3] = l_cell_wire[25];							inform_L[21][3] = l_cell_wire[26];							inform_L[29][3] = l_cell_wire[27];							inform_L[22][3] = l_cell_wire[28];							inform_L[30][3] = l_cell_wire[29];							inform_L[23][3] = l_cell_wire[30];							inform_L[31][3] = l_cell_wire[31];							inform_L[32][3] = l_cell_wire[32];							inform_L[40][3] = l_cell_wire[33];							inform_L[33][3] = l_cell_wire[34];							inform_L[41][3] = l_cell_wire[35];							inform_L[34][3] = l_cell_wire[36];							inform_L[42][3] = l_cell_wire[37];							inform_L[35][3] = l_cell_wire[38];							inform_L[43][3] = l_cell_wire[39];							inform_L[36][3] = l_cell_wire[40];							inform_L[44][3] = l_cell_wire[41];							inform_L[37][3] = l_cell_wire[42];							inform_L[45][3] = l_cell_wire[43];							inform_L[38][3] = l_cell_wire[44];							inform_L[46][3] = l_cell_wire[45];							inform_L[39][3] = l_cell_wire[46];							inform_L[47][3] = l_cell_wire[47];							inform_L[48][3] = l_cell_wire[48];							inform_L[56][3] = l_cell_wire[49];							inform_L[49][3] = l_cell_wire[50];							inform_L[57][3] = l_cell_wire[51];							inform_L[50][3] = l_cell_wire[52];							inform_L[58][3] = l_cell_wire[53];							inform_L[51][3] = l_cell_wire[54];							inform_L[59][3] = l_cell_wire[55];							inform_L[52][3] = l_cell_wire[56];							inform_L[60][3] = l_cell_wire[57];							inform_L[53][3] = l_cell_wire[58];							inform_L[61][3] = l_cell_wire[59];							inform_L[54][3] = l_cell_wire[60];							inform_L[62][3] = l_cell_wire[61];							inform_L[55][3] = l_cell_wire[62];							inform_L[63][3] = l_cell_wire[63];							inform_L[64][3] = l_cell_wire[64];							inform_L[72][3] = l_cell_wire[65];							inform_L[65][3] = l_cell_wire[66];							inform_L[73][3] = l_cell_wire[67];							inform_L[66][3] = l_cell_wire[68];							inform_L[74][3] = l_cell_wire[69];							inform_L[67][3] = l_cell_wire[70];							inform_L[75][3] = l_cell_wire[71];							inform_L[68][3] = l_cell_wire[72];							inform_L[76][3] = l_cell_wire[73];							inform_L[69][3] = l_cell_wire[74];							inform_L[77][3] = l_cell_wire[75];							inform_L[70][3] = l_cell_wire[76];							inform_L[78][3] = l_cell_wire[77];							inform_L[71][3] = l_cell_wire[78];							inform_L[79][3] = l_cell_wire[79];							inform_L[80][3] = l_cell_wire[80];							inform_L[88][3] = l_cell_wire[81];							inform_L[81][3] = l_cell_wire[82];							inform_L[89][3] = l_cell_wire[83];							inform_L[82][3] = l_cell_wire[84];							inform_L[90][3] = l_cell_wire[85];							inform_L[83][3] = l_cell_wire[86];							inform_L[91][3] = l_cell_wire[87];							inform_L[84][3] = l_cell_wire[88];							inform_L[92][3] = l_cell_wire[89];							inform_L[85][3] = l_cell_wire[90];							inform_L[93][3] = l_cell_wire[91];							inform_L[86][3] = l_cell_wire[92];							inform_L[94][3] = l_cell_wire[93];							inform_L[87][3] = l_cell_wire[94];							inform_L[95][3] = l_cell_wire[95];							inform_L[96][3] = l_cell_wire[96];							inform_L[104][3] = l_cell_wire[97];							inform_L[97][3] = l_cell_wire[98];							inform_L[105][3] = l_cell_wire[99];							inform_L[98][3] = l_cell_wire[100];							inform_L[106][3] = l_cell_wire[101];							inform_L[99][3] = l_cell_wire[102];							inform_L[107][3] = l_cell_wire[103];							inform_L[100][3] = l_cell_wire[104];							inform_L[108][3] = l_cell_wire[105];							inform_L[101][3] = l_cell_wire[106];							inform_L[109][3] = l_cell_wire[107];							inform_L[102][3] = l_cell_wire[108];							inform_L[110][3] = l_cell_wire[109];							inform_L[103][3] = l_cell_wire[110];							inform_L[111][3] = l_cell_wire[111];							inform_L[112][3] = l_cell_wire[112];							inform_L[120][3] = l_cell_wire[113];							inform_L[113][3] = l_cell_wire[114];							inform_L[121][3] = l_cell_wire[115];							inform_L[114][3] = l_cell_wire[116];							inform_L[122][3] = l_cell_wire[117];							inform_L[115][3] = l_cell_wire[118];							inform_L[123][3] = l_cell_wire[119];							inform_L[116][3] = l_cell_wire[120];							inform_L[124][3] = l_cell_wire[121];							inform_L[117][3] = l_cell_wire[122];							inform_L[125][3] = l_cell_wire[123];							inform_L[118][3] = l_cell_wire[124];							inform_L[126][3] = l_cell_wire[125];							inform_L[119][3] = l_cell_wire[126];							inform_L[127][3] = l_cell_wire[127];							inform_L[128][3] = l_cell_wire[128];							inform_L[136][3] = l_cell_wire[129];							inform_L[129][3] = l_cell_wire[130];							inform_L[137][3] = l_cell_wire[131];							inform_L[130][3] = l_cell_wire[132];							inform_L[138][3] = l_cell_wire[133];							inform_L[131][3] = l_cell_wire[134];							inform_L[139][3] = l_cell_wire[135];							inform_L[132][3] = l_cell_wire[136];							inform_L[140][3] = l_cell_wire[137];							inform_L[133][3] = l_cell_wire[138];							inform_L[141][3] = l_cell_wire[139];							inform_L[134][3] = l_cell_wire[140];							inform_L[142][3] = l_cell_wire[141];							inform_L[135][3] = l_cell_wire[142];							inform_L[143][3] = l_cell_wire[143];							inform_L[144][3] = l_cell_wire[144];							inform_L[152][3] = l_cell_wire[145];							inform_L[145][3] = l_cell_wire[146];							inform_L[153][3] = l_cell_wire[147];							inform_L[146][3] = l_cell_wire[148];							inform_L[154][3] = l_cell_wire[149];							inform_L[147][3] = l_cell_wire[150];							inform_L[155][3] = l_cell_wire[151];							inform_L[148][3] = l_cell_wire[152];							inform_L[156][3] = l_cell_wire[153];							inform_L[149][3] = l_cell_wire[154];							inform_L[157][3] = l_cell_wire[155];							inform_L[150][3] = l_cell_wire[156];							inform_L[158][3] = l_cell_wire[157];							inform_L[151][3] = l_cell_wire[158];							inform_L[159][3] = l_cell_wire[159];							inform_L[160][3] = l_cell_wire[160];							inform_L[168][3] = l_cell_wire[161];							inform_L[161][3] = l_cell_wire[162];							inform_L[169][3] = l_cell_wire[163];							inform_L[162][3] = l_cell_wire[164];							inform_L[170][3] = l_cell_wire[165];							inform_L[163][3] = l_cell_wire[166];							inform_L[171][3] = l_cell_wire[167];							inform_L[164][3] = l_cell_wire[168];							inform_L[172][3] = l_cell_wire[169];							inform_L[165][3] = l_cell_wire[170];							inform_L[173][3] = l_cell_wire[171];							inform_L[166][3] = l_cell_wire[172];							inform_L[174][3] = l_cell_wire[173];							inform_L[167][3] = l_cell_wire[174];							inform_L[175][3] = l_cell_wire[175];							inform_L[176][3] = l_cell_wire[176];							inform_L[184][3] = l_cell_wire[177];							inform_L[177][3] = l_cell_wire[178];							inform_L[185][3] = l_cell_wire[179];							inform_L[178][3] = l_cell_wire[180];							inform_L[186][3] = l_cell_wire[181];							inform_L[179][3] = l_cell_wire[182];							inform_L[187][3] = l_cell_wire[183];							inform_L[180][3] = l_cell_wire[184];							inform_L[188][3] = l_cell_wire[185];							inform_L[181][3] = l_cell_wire[186];							inform_L[189][3] = l_cell_wire[187];							inform_L[182][3] = l_cell_wire[188];							inform_L[190][3] = l_cell_wire[189];							inform_L[183][3] = l_cell_wire[190];							inform_L[191][3] = l_cell_wire[191];							inform_L[192][3] = l_cell_wire[192];							inform_L[200][3] = l_cell_wire[193];							inform_L[193][3] = l_cell_wire[194];							inform_L[201][3] = l_cell_wire[195];							inform_L[194][3] = l_cell_wire[196];							inform_L[202][3] = l_cell_wire[197];							inform_L[195][3] = l_cell_wire[198];							inform_L[203][3] = l_cell_wire[199];							inform_L[196][3] = l_cell_wire[200];							inform_L[204][3] = l_cell_wire[201];							inform_L[197][3] = l_cell_wire[202];							inform_L[205][3] = l_cell_wire[203];							inform_L[198][3] = l_cell_wire[204];							inform_L[206][3] = l_cell_wire[205];							inform_L[199][3] = l_cell_wire[206];							inform_L[207][3] = l_cell_wire[207];							inform_L[208][3] = l_cell_wire[208];							inform_L[216][3] = l_cell_wire[209];							inform_L[209][3] = l_cell_wire[210];							inform_L[217][3] = l_cell_wire[211];							inform_L[210][3] = l_cell_wire[212];							inform_L[218][3] = l_cell_wire[213];							inform_L[211][3] = l_cell_wire[214];							inform_L[219][3] = l_cell_wire[215];							inform_L[212][3] = l_cell_wire[216];							inform_L[220][3] = l_cell_wire[217];							inform_L[213][3] = l_cell_wire[218];							inform_L[221][3] = l_cell_wire[219];							inform_L[214][3] = l_cell_wire[220];							inform_L[222][3] = l_cell_wire[221];							inform_L[215][3] = l_cell_wire[222];							inform_L[223][3] = l_cell_wire[223];							inform_L[224][3] = l_cell_wire[224];							inform_L[232][3] = l_cell_wire[225];							inform_L[225][3] = l_cell_wire[226];							inform_L[233][3] = l_cell_wire[227];							inform_L[226][3] = l_cell_wire[228];							inform_L[234][3] = l_cell_wire[229];							inform_L[227][3] = l_cell_wire[230];							inform_L[235][3] = l_cell_wire[231];							inform_L[228][3] = l_cell_wire[232];							inform_L[236][3] = l_cell_wire[233];							inform_L[229][3] = l_cell_wire[234];							inform_L[237][3] = l_cell_wire[235];							inform_L[230][3] = l_cell_wire[236];							inform_L[238][3] = l_cell_wire[237];							inform_L[231][3] = l_cell_wire[238];							inform_L[239][3] = l_cell_wire[239];							inform_L[240][3] = l_cell_wire[240];							inform_L[248][3] = l_cell_wire[241];							inform_L[241][3] = l_cell_wire[242];							inform_L[249][3] = l_cell_wire[243];							inform_L[242][3] = l_cell_wire[244];							inform_L[250][3] = l_cell_wire[245];							inform_L[243][3] = l_cell_wire[246];							inform_L[251][3] = l_cell_wire[247];							inform_L[244][3] = l_cell_wire[248];							inform_L[252][3] = l_cell_wire[249];							inform_L[245][3] = l_cell_wire[250];							inform_L[253][3] = l_cell_wire[251];							inform_L[246][3] = l_cell_wire[252];							inform_L[254][3] = l_cell_wire[253];							inform_L[247][3] = l_cell_wire[254];							inform_L[255][3] = l_cell_wire[255];							inform_L[256][3] = l_cell_wire[256];							inform_L[264][3] = l_cell_wire[257];							inform_L[257][3] = l_cell_wire[258];							inform_L[265][3] = l_cell_wire[259];							inform_L[258][3] = l_cell_wire[260];							inform_L[266][3] = l_cell_wire[261];							inform_L[259][3] = l_cell_wire[262];							inform_L[267][3] = l_cell_wire[263];							inform_L[260][3] = l_cell_wire[264];							inform_L[268][3] = l_cell_wire[265];							inform_L[261][3] = l_cell_wire[266];							inform_L[269][3] = l_cell_wire[267];							inform_L[262][3] = l_cell_wire[268];							inform_L[270][3] = l_cell_wire[269];							inform_L[263][3] = l_cell_wire[270];							inform_L[271][3] = l_cell_wire[271];							inform_L[272][3] = l_cell_wire[272];							inform_L[280][3] = l_cell_wire[273];							inform_L[273][3] = l_cell_wire[274];							inform_L[281][3] = l_cell_wire[275];							inform_L[274][3] = l_cell_wire[276];							inform_L[282][3] = l_cell_wire[277];							inform_L[275][3] = l_cell_wire[278];							inform_L[283][3] = l_cell_wire[279];							inform_L[276][3] = l_cell_wire[280];							inform_L[284][3] = l_cell_wire[281];							inform_L[277][3] = l_cell_wire[282];							inform_L[285][3] = l_cell_wire[283];							inform_L[278][3] = l_cell_wire[284];							inform_L[286][3] = l_cell_wire[285];							inform_L[279][3] = l_cell_wire[286];							inform_L[287][3] = l_cell_wire[287];							inform_L[288][3] = l_cell_wire[288];							inform_L[296][3] = l_cell_wire[289];							inform_L[289][3] = l_cell_wire[290];							inform_L[297][3] = l_cell_wire[291];							inform_L[290][3] = l_cell_wire[292];							inform_L[298][3] = l_cell_wire[293];							inform_L[291][3] = l_cell_wire[294];							inform_L[299][3] = l_cell_wire[295];							inform_L[292][3] = l_cell_wire[296];							inform_L[300][3] = l_cell_wire[297];							inform_L[293][3] = l_cell_wire[298];							inform_L[301][3] = l_cell_wire[299];							inform_L[294][3] = l_cell_wire[300];							inform_L[302][3] = l_cell_wire[301];							inform_L[295][3] = l_cell_wire[302];							inform_L[303][3] = l_cell_wire[303];							inform_L[304][3] = l_cell_wire[304];							inform_L[312][3] = l_cell_wire[305];							inform_L[305][3] = l_cell_wire[306];							inform_L[313][3] = l_cell_wire[307];							inform_L[306][3] = l_cell_wire[308];							inform_L[314][3] = l_cell_wire[309];							inform_L[307][3] = l_cell_wire[310];							inform_L[315][3] = l_cell_wire[311];							inform_L[308][3] = l_cell_wire[312];							inform_L[316][3] = l_cell_wire[313];							inform_L[309][3] = l_cell_wire[314];							inform_L[317][3] = l_cell_wire[315];							inform_L[310][3] = l_cell_wire[316];							inform_L[318][3] = l_cell_wire[317];							inform_L[311][3] = l_cell_wire[318];							inform_L[319][3] = l_cell_wire[319];							inform_L[320][3] = l_cell_wire[320];							inform_L[328][3] = l_cell_wire[321];							inform_L[321][3] = l_cell_wire[322];							inform_L[329][3] = l_cell_wire[323];							inform_L[322][3] = l_cell_wire[324];							inform_L[330][3] = l_cell_wire[325];							inform_L[323][3] = l_cell_wire[326];							inform_L[331][3] = l_cell_wire[327];							inform_L[324][3] = l_cell_wire[328];							inform_L[332][3] = l_cell_wire[329];							inform_L[325][3] = l_cell_wire[330];							inform_L[333][3] = l_cell_wire[331];							inform_L[326][3] = l_cell_wire[332];							inform_L[334][3] = l_cell_wire[333];							inform_L[327][3] = l_cell_wire[334];							inform_L[335][3] = l_cell_wire[335];							inform_L[336][3] = l_cell_wire[336];							inform_L[344][3] = l_cell_wire[337];							inform_L[337][3] = l_cell_wire[338];							inform_L[345][3] = l_cell_wire[339];							inform_L[338][3] = l_cell_wire[340];							inform_L[346][3] = l_cell_wire[341];							inform_L[339][3] = l_cell_wire[342];							inform_L[347][3] = l_cell_wire[343];							inform_L[340][3] = l_cell_wire[344];							inform_L[348][3] = l_cell_wire[345];							inform_L[341][3] = l_cell_wire[346];							inform_L[349][3] = l_cell_wire[347];							inform_L[342][3] = l_cell_wire[348];							inform_L[350][3] = l_cell_wire[349];							inform_L[343][3] = l_cell_wire[350];							inform_L[351][3] = l_cell_wire[351];							inform_L[352][3] = l_cell_wire[352];							inform_L[360][3] = l_cell_wire[353];							inform_L[353][3] = l_cell_wire[354];							inform_L[361][3] = l_cell_wire[355];							inform_L[354][3] = l_cell_wire[356];							inform_L[362][3] = l_cell_wire[357];							inform_L[355][3] = l_cell_wire[358];							inform_L[363][3] = l_cell_wire[359];							inform_L[356][3] = l_cell_wire[360];							inform_L[364][3] = l_cell_wire[361];							inform_L[357][3] = l_cell_wire[362];							inform_L[365][3] = l_cell_wire[363];							inform_L[358][3] = l_cell_wire[364];							inform_L[366][3] = l_cell_wire[365];							inform_L[359][3] = l_cell_wire[366];							inform_L[367][3] = l_cell_wire[367];							inform_L[368][3] = l_cell_wire[368];							inform_L[376][3] = l_cell_wire[369];							inform_L[369][3] = l_cell_wire[370];							inform_L[377][3] = l_cell_wire[371];							inform_L[370][3] = l_cell_wire[372];							inform_L[378][3] = l_cell_wire[373];							inform_L[371][3] = l_cell_wire[374];							inform_L[379][3] = l_cell_wire[375];							inform_L[372][3] = l_cell_wire[376];							inform_L[380][3] = l_cell_wire[377];							inform_L[373][3] = l_cell_wire[378];							inform_L[381][3] = l_cell_wire[379];							inform_L[374][3] = l_cell_wire[380];							inform_L[382][3] = l_cell_wire[381];							inform_L[375][3] = l_cell_wire[382];							inform_L[383][3] = l_cell_wire[383];							inform_L[384][3] = l_cell_wire[384];							inform_L[392][3] = l_cell_wire[385];							inform_L[385][3] = l_cell_wire[386];							inform_L[393][3] = l_cell_wire[387];							inform_L[386][3] = l_cell_wire[388];							inform_L[394][3] = l_cell_wire[389];							inform_L[387][3] = l_cell_wire[390];							inform_L[395][3] = l_cell_wire[391];							inform_L[388][3] = l_cell_wire[392];							inform_L[396][3] = l_cell_wire[393];							inform_L[389][3] = l_cell_wire[394];							inform_L[397][3] = l_cell_wire[395];							inform_L[390][3] = l_cell_wire[396];							inform_L[398][3] = l_cell_wire[397];							inform_L[391][3] = l_cell_wire[398];							inform_L[399][3] = l_cell_wire[399];							inform_L[400][3] = l_cell_wire[400];							inform_L[408][3] = l_cell_wire[401];							inform_L[401][3] = l_cell_wire[402];							inform_L[409][3] = l_cell_wire[403];							inform_L[402][3] = l_cell_wire[404];							inform_L[410][3] = l_cell_wire[405];							inform_L[403][3] = l_cell_wire[406];							inform_L[411][3] = l_cell_wire[407];							inform_L[404][3] = l_cell_wire[408];							inform_L[412][3] = l_cell_wire[409];							inform_L[405][3] = l_cell_wire[410];							inform_L[413][3] = l_cell_wire[411];							inform_L[406][3] = l_cell_wire[412];							inform_L[414][3] = l_cell_wire[413];							inform_L[407][3] = l_cell_wire[414];							inform_L[415][3] = l_cell_wire[415];							inform_L[416][3] = l_cell_wire[416];							inform_L[424][3] = l_cell_wire[417];							inform_L[417][3] = l_cell_wire[418];							inform_L[425][3] = l_cell_wire[419];							inform_L[418][3] = l_cell_wire[420];							inform_L[426][3] = l_cell_wire[421];							inform_L[419][3] = l_cell_wire[422];							inform_L[427][3] = l_cell_wire[423];							inform_L[420][3] = l_cell_wire[424];							inform_L[428][3] = l_cell_wire[425];							inform_L[421][3] = l_cell_wire[426];							inform_L[429][3] = l_cell_wire[427];							inform_L[422][3] = l_cell_wire[428];							inform_L[430][3] = l_cell_wire[429];							inform_L[423][3] = l_cell_wire[430];							inform_L[431][3] = l_cell_wire[431];							inform_L[432][3] = l_cell_wire[432];							inform_L[440][3] = l_cell_wire[433];							inform_L[433][3] = l_cell_wire[434];							inform_L[441][3] = l_cell_wire[435];							inform_L[434][3] = l_cell_wire[436];							inform_L[442][3] = l_cell_wire[437];							inform_L[435][3] = l_cell_wire[438];							inform_L[443][3] = l_cell_wire[439];							inform_L[436][3] = l_cell_wire[440];							inform_L[444][3] = l_cell_wire[441];							inform_L[437][3] = l_cell_wire[442];							inform_L[445][3] = l_cell_wire[443];							inform_L[438][3] = l_cell_wire[444];							inform_L[446][3] = l_cell_wire[445];							inform_L[439][3] = l_cell_wire[446];							inform_L[447][3] = l_cell_wire[447];							inform_L[448][3] = l_cell_wire[448];							inform_L[456][3] = l_cell_wire[449];							inform_L[449][3] = l_cell_wire[450];							inform_L[457][3] = l_cell_wire[451];							inform_L[450][3] = l_cell_wire[452];							inform_L[458][3] = l_cell_wire[453];							inform_L[451][3] = l_cell_wire[454];							inform_L[459][3] = l_cell_wire[455];							inform_L[452][3] = l_cell_wire[456];							inform_L[460][3] = l_cell_wire[457];							inform_L[453][3] = l_cell_wire[458];							inform_L[461][3] = l_cell_wire[459];							inform_L[454][3] = l_cell_wire[460];							inform_L[462][3] = l_cell_wire[461];							inform_L[455][3] = l_cell_wire[462];							inform_L[463][3] = l_cell_wire[463];							inform_L[464][3] = l_cell_wire[464];							inform_L[472][3] = l_cell_wire[465];							inform_L[465][3] = l_cell_wire[466];							inform_L[473][3] = l_cell_wire[467];							inform_L[466][3] = l_cell_wire[468];							inform_L[474][3] = l_cell_wire[469];							inform_L[467][3] = l_cell_wire[470];							inform_L[475][3] = l_cell_wire[471];							inform_L[468][3] = l_cell_wire[472];							inform_L[476][3] = l_cell_wire[473];							inform_L[469][3] = l_cell_wire[474];							inform_L[477][3] = l_cell_wire[475];							inform_L[470][3] = l_cell_wire[476];							inform_L[478][3] = l_cell_wire[477];							inform_L[471][3] = l_cell_wire[478];							inform_L[479][3] = l_cell_wire[479];							inform_L[480][3] = l_cell_wire[480];							inform_L[488][3] = l_cell_wire[481];							inform_L[481][3] = l_cell_wire[482];							inform_L[489][3] = l_cell_wire[483];							inform_L[482][3] = l_cell_wire[484];							inform_L[490][3] = l_cell_wire[485];							inform_L[483][3] = l_cell_wire[486];							inform_L[491][3] = l_cell_wire[487];							inform_L[484][3] = l_cell_wire[488];							inform_L[492][3] = l_cell_wire[489];							inform_L[485][3] = l_cell_wire[490];							inform_L[493][3] = l_cell_wire[491];							inform_L[486][3] = l_cell_wire[492];							inform_L[494][3] = l_cell_wire[493];							inform_L[487][3] = l_cell_wire[494];							inform_L[495][3] = l_cell_wire[495];							inform_L[496][3] = l_cell_wire[496];							inform_L[504][3] = l_cell_wire[497];							inform_L[497][3] = l_cell_wire[498];							inform_L[505][3] = l_cell_wire[499];							inform_L[498][3] = l_cell_wire[500];							inform_L[506][3] = l_cell_wire[501];							inform_L[499][3] = l_cell_wire[502];							inform_L[507][3] = l_cell_wire[503];							inform_L[500][3] = l_cell_wire[504];							inform_L[508][3] = l_cell_wire[505];							inform_L[501][3] = l_cell_wire[506];							inform_L[509][3] = l_cell_wire[507];							inform_L[502][3] = l_cell_wire[508];							inform_L[510][3] = l_cell_wire[509];							inform_L[503][3] = l_cell_wire[510];							inform_L[511][3] = l_cell_wire[511];							inform_L[512][3] = l_cell_wire[512];							inform_L[520][3] = l_cell_wire[513];							inform_L[513][3] = l_cell_wire[514];							inform_L[521][3] = l_cell_wire[515];							inform_L[514][3] = l_cell_wire[516];							inform_L[522][3] = l_cell_wire[517];							inform_L[515][3] = l_cell_wire[518];							inform_L[523][3] = l_cell_wire[519];							inform_L[516][3] = l_cell_wire[520];							inform_L[524][3] = l_cell_wire[521];							inform_L[517][3] = l_cell_wire[522];							inform_L[525][3] = l_cell_wire[523];							inform_L[518][3] = l_cell_wire[524];							inform_L[526][3] = l_cell_wire[525];							inform_L[519][3] = l_cell_wire[526];							inform_L[527][3] = l_cell_wire[527];							inform_L[528][3] = l_cell_wire[528];							inform_L[536][3] = l_cell_wire[529];							inform_L[529][3] = l_cell_wire[530];							inform_L[537][3] = l_cell_wire[531];							inform_L[530][3] = l_cell_wire[532];							inform_L[538][3] = l_cell_wire[533];							inform_L[531][3] = l_cell_wire[534];							inform_L[539][3] = l_cell_wire[535];							inform_L[532][3] = l_cell_wire[536];							inform_L[540][3] = l_cell_wire[537];							inform_L[533][3] = l_cell_wire[538];							inform_L[541][3] = l_cell_wire[539];							inform_L[534][3] = l_cell_wire[540];							inform_L[542][3] = l_cell_wire[541];							inform_L[535][3] = l_cell_wire[542];							inform_L[543][3] = l_cell_wire[543];							inform_L[544][3] = l_cell_wire[544];							inform_L[552][3] = l_cell_wire[545];							inform_L[545][3] = l_cell_wire[546];							inform_L[553][3] = l_cell_wire[547];							inform_L[546][3] = l_cell_wire[548];							inform_L[554][3] = l_cell_wire[549];							inform_L[547][3] = l_cell_wire[550];							inform_L[555][3] = l_cell_wire[551];							inform_L[548][3] = l_cell_wire[552];							inform_L[556][3] = l_cell_wire[553];							inform_L[549][3] = l_cell_wire[554];							inform_L[557][3] = l_cell_wire[555];							inform_L[550][3] = l_cell_wire[556];							inform_L[558][3] = l_cell_wire[557];							inform_L[551][3] = l_cell_wire[558];							inform_L[559][3] = l_cell_wire[559];							inform_L[560][3] = l_cell_wire[560];							inform_L[568][3] = l_cell_wire[561];							inform_L[561][3] = l_cell_wire[562];							inform_L[569][3] = l_cell_wire[563];							inform_L[562][3] = l_cell_wire[564];							inform_L[570][3] = l_cell_wire[565];							inform_L[563][3] = l_cell_wire[566];							inform_L[571][3] = l_cell_wire[567];							inform_L[564][3] = l_cell_wire[568];							inform_L[572][3] = l_cell_wire[569];							inform_L[565][3] = l_cell_wire[570];							inform_L[573][3] = l_cell_wire[571];							inform_L[566][3] = l_cell_wire[572];							inform_L[574][3] = l_cell_wire[573];							inform_L[567][3] = l_cell_wire[574];							inform_L[575][3] = l_cell_wire[575];							inform_L[576][3] = l_cell_wire[576];							inform_L[584][3] = l_cell_wire[577];							inform_L[577][3] = l_cell_wire[578];							inform_L[585][3] = l_cell_wire[579];							inform_L[578][3] = l_cell_wire[580];							inform_L[586][3] = l_cell_wire[581];							inform_L[579][3] = l_cell_wire[582];							inform_L[587][3] = l_cell_wire[583];							inform_L[580][3] = l_cell_wire[584];							inform_L[588][3] = l_cell_wire[585];							inform_L[581][3] = l_cell_wire[586];							inform_L[589][3] = l_cell_wire[587];							inform_L[582][3] = l_cell_wire[588];							inform_L[590][3] = l_cell_wire[589];							inform_L[583][3] = l_cell_wire[590];							inform_L[591][3] = l_cell_wire[591];							inform_L[592][3] = l_cell_wire[592];							inform_L[600][3] = l_cell_wire[593];							inform_L[593][3] = l_cell_wire[594];							inform_L[601][3] = l_cell_wire[595];							inform_L[594][3] = l_cell_wire[596];							inform_L[602][3] = l_cell_wire[597];							inform_L[595][3] = l_cell_wire[598];							inform_L[603][3] = l_cell_wire[599];							inform_L[596][3] = l_cell_wire[600];							inform_L[604][3] = l_cell_wire[601];							inform_L[597][3] = l_cell_wire[602];							inform_L[605][3] = l_cell_wire[603];							inform_L[598][3] = l_cell_wire[604];							inform_L[606][3] = l_cell_wire[605];							inform_L[599][3] = l_cell_wire[606];							inform_L[607][3] = l_cell_wire[607];							inform_L[608][3] = l_cell_wire[608];							inform_L[616][3] = l_cell_wire[609];							inform_L[609][3] = l_cell_wire[610];							inform_L[617][3] = l_cell_wire[611];							inform_L[610][3] = l_cell_wire[612];							inform_L[618][3] = l_cell_wire[613];							inform_L[611][3] = l_cell_wire[614];							inform_L[619][3] = l_cell_wire[615];							inform_L[612][3] = l_cell_wire[616];							inform_L[620][3] = l_cell_wire[617];							inform_L[613][3] = l_cell_wire[618];							inform_L[621][3] = l_cell_wire[619];							inform_L[614][3] = l_cell_wire[620];							inform_L[622][3] = l_cell_wire[621];							inform_L[615][3] = l_cell_wire[622];							inform_L[623][3] = l_cell_wire[623];							inform_L[624][3] = l_cell_wire[624];							inform_L[632][3] = l_cell_wire[625];							inform_L[625][3] = l_cell_wire[626];							inform_L[633][3] = l_cell_wire[627];							inform_L[626][3] = l_cell_wire[628];							inform_L[634][3] = l_cell_wire[629];							inform_L[627][3] = l_cell_wire[630];							inform_L[635][3] = l_cell_wire[631];							inform_L[628][3] = l_cell_wire[632];							inform_L[636][3] = l_cell_wire[633];							inform_L[629][3] = l_cell_wire[634];							inform_L[637][3] = l_cell_wire[635];							inform_L[630][3] = l_cell_wire[636];							inform_L[638][3] = l_cell_wire[637];							inform_L[631][3] = l_cell_wire[638];							inform_L[639][3] = l_cell_wire[639];							inform_L[640][3] = l_cell_wire[640];							inform_L[648][3] = l_cell_wire[641];							inform_L[641][3] = l_cell_wire[642];							inform_L[649][3] = l_cell_wire[643];							inform_L[642][3] = l_cell_wire[644];							inform_L[650][3] = l_cell_wire[645];							inform_L[643][3] = l_cell_wire[646];							inform_L[651][3] = l_cell_wire[647];							inform_L[644][3] = l_cell_wire[648];							inform_L[652][3] = l_cell_wire[649];							inform_L[645][3] = l_cell_wire[650];							inform_L[653][3] = l_cell_wire[651];							inform_L[646][3] = l_cell_wire[652];							inform_L[654][3] = l_cell_wire[653];							inform_L[647][3] = l_cell_wire[654];							inform_L[655][3] = l_cell_wire[655];							inform_L[656][3] = l_cell_wire[656];							inform_L[664][3] = l_cell_wire[657];							inform_L[657][3] = l_cell_wire[658];							inform_L[665][3] = l_cell_wire[659];							inform_L[658][3] = l_cell_wire[660];							inform_L[666][3] = l_cell_wire[661];							inform_L[659][3] = l_cell_wire[662];							inform_L[667][3] = l_cell_wire[663];							inform_L[660][3] = l_cell_wire[664];							inform_L[668][3] = l_cell_wire[665];							inform_L[661][3] = l_cell_wire[666];							inform_L[669][3] = l_cell_wire[667];							inform_L[662][3] = l_cell_wire[668];							inform_L[670][3] = l_cell_wire[669];							inform_L[663][3] = l_cell_wire[670];							inform_L[671][3] = l_cell_wire[671];							inform_L[672][3] = l_cell_wire[672];							inform_L[680][3] = l_cell_wire[673];							inform_L[673][3] = l_cell_wire[674];							inform_L[681][3] = l_cell_wire[675];							inform_L[674][3] = l_cell_wire[676];							inform_L[682][3] = l_cell_wire[677];							inform_L[675][3] = l_cell_wire[678];							inform_L[683][3] = l_cell_wire[679];							inform_L[676][3] = l_cell_wire[680];							inform_L[684][3] = l_cell_wire[681];							inform_L[677][3] = l_cell_wire[682];							inform_L[685][3] = l_cell_wire[683];							inform_L[678][3] = l_cell_wire[684];							inform_L[686][3] = l_cell_wire[685];							inform_L[679][3] = l_cell_wire[686];							inform_L[687][3] = l_cell_wire[687];							inform_L[688][3] = l_cell_wire[688];							inform_L[696][3] = l_cell_wire[689];							inform_L[689][3] = l_cell_wire[690];							inform_L[697][3] = l_cell_wire[691];							inform_L[690][3] = l_cell_wire[692];							inform_L[698][3] = l_cell_wire[693];							inform_L[691][3] = l_cell_wire[694];							inform_L[699][3] = l_cell_wire[695];							inform_L[692][3] = l_cell_wire[696];							inform_L[700][3] = l_cell_wire[697];							inform_L[693][3] = l_cell_wire[698];							inform_L[701][3] = l_cell_wire[699];							inform_L[694][3] = l_cell_wire[700];							inform_L[702][3] = l_cell_wire[701];							inform_L[695][3] = l_cell_wire[702];							inform_L[703][3] = l_cell_wire[703];							inform_L[704][3] = l_cell_wire[704];							inform_L[712][3] = l_cell_wire[705];							inform_L[705][3] = l_cell_wire[706];							inform_L[713][3] = l_cell_wire[707];							inform_L[706][3] = l_cell_wire[708];							inform_L[714][3] = l_cell_wire[709];							inform_L[707][3] = l_cell_wire[710];							inform_L[715][3] = l_cell_wire[711];							inform_L[708][3] = l_cell_wire[712];							inform_L[716][3] = l_cell_wire[713];							inform_L[709][3] = l_cell_wire[714];							inform_L[717][3] = l_cell_wire[715];							inform_L[710][3] = l_cell_wire[716];							inform_L[718][3] = l_cell_wire[717];							inform_L[711][3] = l_cell_wire[718];							inform_L[719][3] = l_cell_wire[719];							inform_L[720][3] = l_cell_wire[720];							inform_L[728][3] = l_cell_wire[721];							inform_L[721][3] = l_cell_wire[722];							inform_L[729][3] = l_cell_wire[723];							inform_L[722][3] = l_cell_wire[724];							inform_L[730][3] = l_cell_wire[725];							inform_L[723][3] = l_cell_wire[726];							inform_L[731][3] = l_cell_wire[727];							inform_L[724][3] = l_cell_wire[728];							inform_L[732][3] = l_cell_wire[729];							inform_L[725][3] = l_cell_wire[730];							inform_L[733][3] = l_cell_wire[731];							inform_L[726][3] = l_cell_wire[732];							inform_L[734][3] = l_cell_wire[733];							inform_L[727][3] = l_cell_wire[734];							inform_L[735][3] = l_cell_wire[735];							inform_L[736][3] = l_cell_wire[736];							inform_L[744][3] = l_cell_wire[737];							inform_L[737][3] = l_cell_wire[738];							inform_L[745][3] = l_cell_wire[739];							inform_L[738][3] = l_cell_wire[740];							inform_L[746][3] = l_cell_wire[741];							inform_L[739][3] = l_cell_wire[742];							inform_L[747][3] = l_cell_wire[743];							inform_L[740][3] = l_cell_wire[744];							inform_L[748][3] = l_cell_wire[745];							inform_L[741][3] = l_cell_wire[746];							inform_L[749][3] = l_cell_wire[747];							inform_L[742][3] = l_cell_wire[748];							inform_L[750][3] = l_cell_wire[749];							inform_L[743][3] = l_cell_wire[750];							inform_L[751][3] = l_cell_wire[751];							inform_L[752][3] = l_cell_wire[752];							inform_L[760][3] = l_cell_wire[753];							inform_L[753][3] = l_cell_wire[754];							inform_L[761][3] = l_cell_wire[755];							inform_L[754][3] = l_cell_wire[756];							inform_L[762][3] = l_cell_wire[757];							inform_L[755][3] = l_cell_wire[758];							inform_L[763][3] = l_cell_wire[759];							inform_L[756][3] = l_cell_wire[760];							inform_L[764][3] = l_cell_wire[761];							inform_L[757][3] = l_cell_wire[762];							inform_L[765][3] = l_cell_wire[763];							inform_L[758][3] = l_cell_wire[764];							inform_L[766][3] = l_cell_wire[765];							inform_L[759][3] = l_cell_wire[766];							inform_L[767][3] = l_cell_wire[767];							inform_L[768][3] = l_cell_wire[768];							inform_L[776][3] = l_cell_wire[769];							inform_L[769][3] = l_cell_wire[770];							inform_L[777][3] = l_cell_wire[771];							inform_L[770][3] = l_cell_wire[772];							inform_L[778][3] = l_cell_wire[773];							inform_L[771][3] = l_cell_wire[774];							inform_L[779][3] = l_cell_wire[775];							inform_L[772][3] = l_cell_wire[776];							inform_L[780][3] = l_cell_wire[777];							inform_L[773][3] = l_cell_wire[778];							inform_L[781][3] = l_cell_wire[779];							inform_L[774][3] = l_cell_wire[780];							inform_L[782][3] = l_cell_wire[781];							inform_L[775][3] = l_cell_wire[782];							inform_L[783][3] = l_cell_wire[783];							inform_L[784][3] = l_cell_wire[784];							inform_L[792][3] = l_cell_wire[785];							inform_L[785][3] = l_cell_wire[786];							inform_L[793][3] = l_cell_wire[787];							inform_L[786][3] = l_cell_wire[788];							inform_L[794][3] = l_cell_wire[789];							inform_L[787][3] = l_cell_wire[790];							inform_L[795][3] = l_cell_wire[791];							inform_L[788][3] = l_cell_wire[792];							inform_L[796][3] = l_cell_wire[793];							inform_L[789][3] = l_cell_wire[794];							inform_L[797][3] = l_cell_wire[795];							inform_L[790][3] = l_cell_wire[796];							inform_L[798][3] = l_cell_wire[797];							inform_L[791][3] = l_cell_wire[798];							inform_L[799][3] = l_cell_wire[799];							inform_L[800][3] = l_cell_wire[800];							inform_L[808][3] = l_cell_wire[801];							inform_L[801][3] = l_cell_wire[802];							inform_L[809][3] = l_cell_wire[803];							inform_L[802][3] = l_cell_wire[804];							inform_L[810][3] = l_cell_wire[805];							inform_L[803][3] = l_cell_wire[806];							inform_L[811][3] = l_cell_wire[807];							inform_L[804][3] = l_cell_wire[808];							inform_L[812][3] = l_cell_wire[809];							inform_L[805][3] = l_cell_wire[810];							inform_L[813][3] = l_cell_wire[811];							inform_L[806][3] = l_cell_wire[812];							inform_L[814][3] = l_cell_wire[813];							inform_L[807][3] = l_cell_wire[814];							inform_L[815][3] = l_cell_wire[815];							inform_L[816][3] = l_cell_wire[816];							inform_L[824][3] = l_cell_wire[817];							inform_L[817][3] = l_cell_wire[818];							inform_L[825][3] = l_cell_wire[819];							inform_L[818][3] = l_cell_wire[820];							inform_L[826][3] = l_cell_wire[821];							inform_L[819][3] = l_cell_wire[822];							inform_L[827][3] = l_cell_wire[823];							inform_L[820][3] = l_cell_wire[824];							inform_L[828][3] = l_cell_wire[825];							inform_L[821][3] = l_cell_wire[826];							inform_L[829][3] = l_cell_wire[827];							inform_L[822][3] = l_cell_wire[828];							inform_L[830][3] = l_cell_wire[829];							inform_L[823][3] = l_cell_wire[830];							inform_L[831][3] = l_cell_wire[831];							inform_L[832][3] = l_cell_wire[832];							inform_L[840][3] = l_cell_wire[833];							inform_L[833][3] = l_cell_wire[834];							inform_L[841][3] = l_cell_wire[835];							inform_L[834][3] = l_cell_wire[836];							inform_L[842][3] = l_cell_wire[837];							inform_L[835][3] = l_cell_wire[838];							inform_L[843][3] = l_cell_wire[839];							inform_L[836][3] = l_cell_wire[840];							inform_L[844][3] = l_cell_wire[841];							inform_L[837][3] = l_cell_wire[842];							inform_L[845][3] = l_cell_wire[843];							inform_L[838][3] = l_cell_wire[844];							inform_L[846][3] = l_cell_wire[845];							inform_L[839][3] = l_cell_wire[846];							inform_L[847][3] = l_cell_wire[847];							inform_L[848][3] = l_cell_wire[848];							inform_L[856][3] = l_cell_wire[849];							inform_L[849][3] = l_cell_wire[850];							inform_L[857][3] = l_cell_wire[851];							inform_L[850][3] = l_cell_wire[852];							inform_L[858][3] = l_cell_wire[853];							inform_L[851][3] = l_cell_wire[854];							inform_L[859][3] = l_cell_wire[855];							inform_L[852][3] = l_cell_wire[856];							inform_L[860][3] = l_cell_wire[857];							inform_L[853][3] = l_cell_wire[858];							inform_L[861][3] = l_cell_wire[859];							inform_L[854][3] = l_cell_wire[860];							inform_L[862][3] = l_cell_wire[861];							inform_L[855][3] = l_cell_wire[862];							inform_L[863][3] = l_cell_wire[863];							inform_L[864][3] = l_cell_wire[864];							inform_L[872][3] = l_cell_wire[865];							inform_L[865][3] = l_cell_wire[866];							inform_L[873][3] = l_cell_wire[867];							inform_L[866][3] = l_cell_wire[868];							inform_L[874][3] = l_cell_wire[869];							inform_L[867][3] = l_cell_wire[870];							inform_L[875][3] = l_cell_wire[871];							inform_L[868][3] = l_cell_wire[872];							inform_L[876][3] = l_cell_wire[873];							inform_L[869][3] = l_cell_wire[874];							inform_L[877][3] = l_cell_wire[875];							inform_L[870][3] = l_cell_wire[876];							inform_L[878][3] = l_cell_wire[877];							inform_L[871][3] = l_cell_wire[878];							inform_L[879][3] = l_cell_wire[879];							inform_L[880][3] = l_cell_wire[880];							inform_L[888][3] = l_cell_wire[881];							inform_L[881][3] = l_cell_wire[882];							inform_L[889][3] = l_cell_wire[883];							inform_L[882][3] = l_cell_wire[884];							inform_L[890][3] = l_cell_wire[885];							inform_L[883][3] = l_cell_wire[886];							inform_L[891][3] = l_cell_wire[887];							inform_L[884][3] = l_cell_wire[888];							inform_L[892][3] = l_cell_wire[889];							inform_L[885][3] = l_cell_wire[890];							inform_L[893][3] = l_cell_wire[891];							inform_L[886][3] = l_cell_wire[892];							inform_L[894][3] = l_cell_wire[893];							inform_L[887][3] = l_cell_wire[894];							inform_L[895][3] = l_cell_wire[895];							inform_L[896][3] = l_cell_wire[896];							inform_L[904][3] = l_cell_wire[897];							inform_L[897][3] = l_cell_wire[898];							inform_L[905][3] = l_cell_wire[899];							inform_L[898][3] = l_cell_wire[900];							inform_L[906][3] = l_cell_wire[901];							inform_L[899][3] = l_cell_wire[902];							inform_L[907][3] = l_cell_wire[903];							inform_L[900][3] = l_cell_wire[904];							inform_L[908][3] = l_cell_wire[905];							inform_L[901][3] = l_cell_wire[906];							inform_L[909][3] = l_cell_wire[907];							inform_L[902][3] = l_cell_wire[908];							inform_L[910][3] = l_cell_wire[909];							inform_L[903][3] = l_cell_wire[910];							inform_L[911][3] = l_cell_wire[911];							inform_L[912][3] = l_cell_wire[912];							inform_L[920][3] = l_cell_wire[913];							inform_L[913][3] = l_cell_wire[914];							inform_L[921][3] = l_cell_wire[915];							inform_L[914][3] = l_cell_wire[916];							inform_L[922][3] = l_cell_wire[917];							inform_L[915][3] = l_cell_wire[918];							inform_L[923][3] = l_cell_wire[919];							inform_L[916][3] = l_cell_wire[920];							inform_L[924][3] = l_cell_wire[921];							inform_L[917][3] = l_cell_wire[922];							inform_L[925][3] = l_cell_wire[923];							inform_L[918][3] = l_cell_wire[924];							inform_L[926][3] = l_cell_wire[925];							inform_L[919][3] = l_cell_wire[926];							inform_L[927][3] = l_cell_wire[927];							inform_L[928][3] = l_cell_wire[928];							inform_L[936][3] = l_cell_wire[929];							inform_L[929][3] = l_cell_wire[930];							inform_L[937][3] = l_cell_wire[931];							inform_L[930][3] = l_cell_wire[932];							inform_L[938][3] = l_cell_wire[933];							inform_L[931][3] = l_cell_wire[934];							inform_L[939][3] = l_cell_wire[935];							inform_L[932][3] = l_cell_wire[936];							inform_L[940][3] = l_cell_wire[937];							inform_L[933][3] = l_cell_wire[938];							inform_L[941][3] = l_cell_wire[939];							inform_L[934][3] = l_cell_wire[940];							inform_L[942][3] = l_cell_wire[941];							inform_L[935][3] = l_cell_wire[942];							inform_L[943][3] = l_cell_wire[943];							inform_L[944][3] = l_cell_wire[944];							inform_L[952][3] = l_cell_wire[945];							inform_L[945][3] = l_cell_wire[946];							inform_L[953][3] = l_cell_wire[947];							inform_L[946][3] = l_cell_wire[948];							inform_L[954][3] = l_cell_wire[949];							inform_L[947][3] = l_cell_wire[950];							inform_L[955][3] = l_cell_wire[951];							inform_L[948][3] = l_cell_wire[952];							inform_L[956][3] = l_cell_wire[953];							inform_L[949][3] = l_cell_wire[954];							inform_L[957][3] = l_cell_wire[955];							inform_L[950][3] = l_cell_wire[956];							inform_L[958][3] = l_cell_wire[957];							inform_L[951][3] = l_cell_wire[958];							inform_L[959][3] = l_cell_wire[959];							inform_L[960][3] = l_cell_wire[960];							inform_L[968][3] = l_cell_wire[961];							inform_L[961][3] = l_cell_wire[962];							inform_L[969][3] = l_cell_wire[963];							inform_L[962][3] = l_cell_wire[964];							inform_L[970][3] = l_cell_wire[965];							inform_L[963][3] = l_cell_wire[966];							inform_L[971][3] = l_cell_wire[967];							inform_L[964][3] = l_cell_wire[968];							inform_L[972][3] = l_cell_wire[969];							inform_L[965][3] = l_cell_wire[970];							inform_L[973][3] = l_cell_wire[971];							inform_L[966][3] = l_cell_wire[972];							inform_L[974][3] = l_cell_wire[973];							inform_L[967][3] = l_cell_wire[974];							inform_L[975][3] = l_cell_wire[975];							inform_L[976][3] = l_cell_wire[976];							inform_L[984][3] = l_cell_wire[977];							inform_L[977][3] = l_cell_wire[978];							inform_L[985][3] = l_cell_wire[979];							inform_L[978][3] = l_cell_wire[980];							inform_L[986][3] = l_cell_wire[981];							inform_L[979][3] = l_cell_wire[982];							inform_L[987][3] = l_cell_wire[983];							inform_L[980][3] = l_cell_wire[984];							inform_L[988][3] = l_cell_wire[985];							inform_L[981][3] = l_cell_wire[986];							inform_L[989][3] = l_cell_wire[987];							inform_L[982][3] = l_cell_wire[988];							inform_L[990][3] = l_cell_wire[989];							inform_L[983][3] = l_cell_wire[990];							inform_L[991][3] = l_cell_wire[991];							inform_L[992][3] = l_cell_wire[992];							inform_L[1000][3] = l_cell_wire[993];							inform_L[993][3] = l_cell_wire[994];							inform_L[1001][3] = l_cell_wire[995];							inform_L[994][3] = l_cell_wire[996];							inform_L[1002][3] = l_cell_wire[997];							inform_L[995][3] = l_cell_wire[998];							inform_L[1003][3] = l_cell_wire[999];							inform_L[996][3] = l_cell_wire[1000];							inform_L[1004][3] = l_cell_wire[1001];							inform_L[997][3] = l_cell_wire[1002];							inform_L[1005][3] = l_cell_wire[1003];							inform_L[998][3] = l_cell_wire[1004];							inform_L[1006][3] = l_cell_wire[1005];							inform_L[999][3] = l_cell_wire[1006];							inform_L[1007][3] = l_cell_wire[1007];							inform_L[1008][3] = l_cell_wire[1008];							inform_L[1016][3] = l_cell_wire[1009];							inform_L[1009][3] = l_cell_wire[1010];							inform_L[1017][3] = l_cell_wire[1011];							inform_L[1010][3] = l_cell_wire[1012];							inform_L[1018][3] = l_cell_wire[1013];							inform_L[1011][3] = l_cell_wire[1014];							inform_L[1019][3] = l_cell_wire[1015];							inform_L[1012][3] = l_cell_wire[1016];							inform_L[1020][3] = l_cell_wire[1017];							inform_L[1013][3] = l_cell_wire[1018];							inform_L[1021][3] = l_cell_wire[1019];							inform_L[1014][3] = l_cell_wire[1020];							inform_L[1022][3] = l_cell_wire[1021];							inform_L[1015][3] = l_cell_wire[1022];							inform_L[1023][3] = l_cell_wire[1023];						end
						5:						begin							inform_R[0][5] = r_cell_wire[0];							inform_R[16][5] = r_cell_wire[1];							inform_R[1][5] = r_cell_wire[2];							inform_R[17][5] = r_cell_wire[3];							inform_R[2][5] = r_cell_wire[4];							inform_R[18][5] = r_cell_wire[5];							inform_R[3][5] = r_cell_wire[6];							inform_R[19][5] = r_cell_wire[7];							inform_R[4][5] = r_cell_wire[8];							inform_R[20][5] = r_cell_wire[9];							inform_R[5][5] = r_cell_wire[10];							inform_R[21][5] = r_cell_wire[11];							inform_R[6][5] = r_cell_wire[12];							inform_R[22][5] = r_cell_wire[13];							inform_R[7][5] = r_cell_wire[14];							inform_R[23][5] = r_cell_wire[15];							inform_R[8][5] = r_cell_wire[16];							inform_R[24][5] = r_cell_wire[17];							inform_R[9][5] = r_cell_wire[18];							inform_R[25][5] = r_cell_wire[19];							inform_R[10][5] = r_cell_wire[20];							inform_R[26][5] = r_cell_wire[21];							inform_R[11][5] = r_cell_wire[22];							inform_R[27][5] = r_cell_wire[23];							inform_R[12][5] = r_cell_wire[24];							inform_R[28][5] = r_cell_wire[25];							inform_R[13][5] = r_cell_wire[26];							inform_R[29][5] = r_cell_wire[27];							inform_R[14][5] = r_cell_wire[28];							inform_R[30][5] = r_cell_wire[29];							inform_R[15][5] = r_cell_wire[30];							inform_R[31][5] = r_cell_wire[31];							inform_R[32][5] = r_cell_wire[32];							inform_R[48][5] = r_cell_wire[33];							inform_R[33][5] = r_cell_wire[34];							inform_R[49][5] = r_cell_wire[35];							inform_R[34][5] = r_cell_wire[36];							inform_R[50][5] = r_cell_wire[37];							inform_R[35][5] = r_cell_wire[38];							inform_R[51][5] = r_cell_wire[39];							inform_R[36][5] = r_cell_wire[40];							inform_R[52][5] = r_cell_wire[41];							inform_R[37][5] = r_cell_wire[42];							inform_R[53][5] = r_cell_wire[43];							inform_R[38][5] = r_cell_wire[44];							inform_R[54][5] = r_cell_wire[45];							inform_R[39][5] = r_cell_wire[46];							inform_R[55][5] = r_cell_wire[47];							inform_R[40][5] = r_cell_wire[48];							inform_R[56][5] = r_cell_wire[49];							inform_R[41][5] = r_cell_wire[50];							inform_R[57][5] = r_cell_wire[51];							inform_R[42][5] = r_cell_wire[52];							inform_R[58][5] = r_cell_wire[53];							inform_R[43][5] = r_cell_wire[54];							inform_R[59][5] = r_cell_wire[55];							inform_R[44][5] = r_cell_wire[56];							inform_R[60][5] = r_cell_wire[57];							inform_R[45][5] = r_cell_wire[58];							inform_R[61][5] = r_cell_wire[59];							inform_R[46][5] = r_cell_wire[60];							inform_R[62][5] = r_cell_wire[61];							inform_R[47][5] = r_cell_wire[62];							inform_R[63][5] = r_cell_wire[63];							inform_R[64][5] = r_cell_wire[64];							inform_R[80][5] = r_cell_wire[65];							inform_R[65][5] = r_cell_wire[66];							inform_R[81][5] = r_cell_wire[67];							inform_R[66][5] = r_cell_wire[68];							inform_R[82][5] = r_cell_wire[69];							inform_R[67][5] = r_cell_wire[70];							inform_R[83][5] = r_cell_wire[71];							inform_R[68][5] = r_cell_wire[72];							inform_R[84][5] = r_cell_wire[73];							inform_R[69][5] = r_cell_wire[74];							inform_R[85][5] = r_cell_wire[75];							inform_R[70][5] = r_cell_wire[76];							inform_R[86][5] = r_cell_wire[77];							inform_R[71][5] = r_cell_wire[78];							inform_R[87][5] = r_cell_wire[79];							inform_R[72][5] = r_cell_wire[80];							inform_R[88][5] = r_cell_wire[81];							inform_R[73][5] = r_cell_wire[82];							inform_R[89][5] = r_cell_wire[83];							inform_R[74][5] = r_cell_wire[84];							inform_R[90][5] = r_cell_wire[85];							inform_R[75][5] = r_cell_wire[86];							inform_R[91][5] = r_cell_wire[87];							inform_R[76][5] = r_cell_wire[88];							inform_R[92][5] = r_cell_wire[89];							inform_R[77][5] = r_cell_wire[90];							inform_R[93][5] = r_cell_wire[91];							inform_R[78][5] = r_cell_wire[92];							inform_R[94][5] = r_cell_wire[93];							inform_R[79][5] = r_cell_wire[94];							inform_R[95][5] = r_cell_wire[95];							inform_R[96][5] = r_cell_wire[96];							inform_R[112][5] = r_cell_wire[97];							inform_R[97][5] = r_cell_wire[98];							inform_R[113][5] = r_cell_wire[99];							inform_R[98][5] = r_cell_wire[100];							inform_R[114][5] = r_cell_wire[101];							inform_R[99][5] = r_cell_wire[102];							inform_R[115][5] = r_cell_wire[103];							inform_R[100][5] = r_cell_wire[104];							inform_R[116][5] = r_cell_wire[105];							inform_R[101][5] = r_cell_wire[106];							inform_R[117][5] = r_cell_wire[107];							inform_R[102][5] = r_cell_wire[108];							inform_R[118][5] = r_cell_wire[109];							inform_R[103][5] = r_cell_wire[110];							inform_R[119][5] = r_cell_wire[111];							inform_R[104][5] = r_cell_wire[112];							inform_R[120][5] = r_cell_wire[113];							inform_R[105][5] = r_cell_wire[114];							inform_R[121][5] = r_cell_wire[115];							inform_R[106][5] = r_cell_wire[116];							inform_R[122][5] = r_cell_wire[117];							inform_R[107][5] = r_cell_wire[118];							inform_R[123][5] = r_cell_wire[119];							inform_R[108][5] = r_cell_wire[120];							inform_R[124][5] = r_cell_wire[121];							inform_R[109][5] = r_cell_wire[122];							inform_R[125][5] = r_cell_wire[123];							inform_R[110][5] = r_cell_wire[124];							inform_R[126][5] = r_cell_wire[125];							inform_R[111][5] = r_cell_wire[126];							inform_R[127][5] = r_cell_wire[127];							inform_R[128][5] = r_cell_wire[128];							inform_R[144][5] = r_cell_wire[129];							inform_R[129][5] = r_cell_wire[130];							inform_R[145][5] = r_cell_wire[131];							inform_R[130][5] = r_cell_wire[132];							inform_R[146][5] = r_cell_wire[133];							inform_R[131][5] = r_cell_wire[134];							inform_R[147][5] = r_cell_wire[135];							inform_R[132][5] = r_cell_wire[136];							inform_R[148][5] = r_cell_wire[137];							inform_R[133][5] = r_cell_wire[138];							inform_R[149][5] = r_cell_wire[139];							inform_R[134][5] = r_cell_wire[140];							inform_R[150][5] = r_cell_wire[141];							inform_R[135][5] = r_cell_wire[142];							inform_R[151][5] = r_cell_wire[143];							inform_R[136][5] = r_cell_wire[144];							inform_R[152][5] = r_cell_wire[145];							inform_R[137][5] = r_cell_wire[146];							inform_R[153][5] = r_cell_wire[147];							inform_R[138][5] = r_cell_wire[148];							inform_R[154][5] = r_cell_wire[149];							inform_R[139][5] = r_cell_wire[150];							inform_R[155][5] = r_cell_wire[151];							inform_R[140][5] = r_cell_wire[152];							inform_R[156][5] = r_cell_wire[153];							inform_R[141][5] = r_cell_wire[154];							inform_R[157][5] = r_cell_wire[155];							inform_R[142][5] = r_cell_wire[156];							inform_R[158][5] = r_cell_wire[157];							inform_R[143][5] = r_cell_wire[158];							inform_R[159][5] = r_cell_wire[159];							inform_R[160][5] = r_cell_wire[160];							inform_R[176][5] = r_cell_wire[161];							inform_R[161][5] = r_cell_wire[162];							inform_R[177][5] = r_cell_wire[163];							inform_R[162][5] = r_cell_wire[164];							inform_R[178][5] = r_cell_wire[165];							inform_R[163][5] = r_cell_wire[166];							inform_R[179][5] = r_cell_wire[167];							inform_R[164][5] = r_cell_wire[168];							inform_R[180][5] = r_cell_wire[169];							inform_R[165][5] = r_cell_wire[170];							inform_R[181][5] = r_cell_wire[171];							inform_R[166][5] = r_cell_wire[172];							inform_R[182][5] = r_cell_wire[173];							inform_R[167][5] = r_cell_wire[174];							inform_R[183][5] = r_cell_wire[175];							inform_R[168][5] = r_cell_wire[176];							inform_R[184][5] = r_cell_wire[177];							inform_R[169][5] = r_cell_wire[178];							inform_R[185][5] = r_cell_wire[179];							inform_R[170][5] = r_cell_wire[180];							inform_R[186][5] = r_cell_wire[181];							inform_R[171][5] = r_cell_wire[182];							inform_R[187][5] = r_cell_wire[183];							inform_R[172][5] = r_cell_wire[184];							inform_R[188][5] = r_cell_wire[185];							inform_R[173][5] = r_cell_wire[186];							inform_R[189][5] = r_cell_wire[187];							inform_R[174][5] = r_cell_wire[188];							inform_R[190][5] = r_cell_wire[189];							inform_R[175][5] = r_cell_wire[190];							inform_R[191][5] = r_cell_wire[191];							inform_R[192][5] = r_cell_wire[192];							inform_R[208][5] = r_cell_wire[193];							inform_R[193][5] = r_cell_wire[194];							inform_R[209][5] = r_cell_wire[195];							inform_R[194][5] = r_cell_wire[196];							inform_R[210][5] = r_cell_wire[197];							inform_R[195][5] = r_cell_wire[198];							inform_R[211][5] = r_cell_wire[199];							inform_R[196][5] = r_cell_wire[200];							inform_R[212][5] = r_cell_wire[201];							inform_R[197][5] = r_cell_wire[202];							inform_R[213][5] = r_cell_wire[203];							inform_R[198][5] = r_cell_wire[204];							inform_R[214][5] = r_cell_wire[205];							inform_R[199][5] = r_cell_wire[206];							inform_R[215][5] = r_cell_wire[207];							inform_R[200][5] = r_cell_wire[208];							inform_R[216][5] = r_cell_wire[209];							inform_R[201][5] = r_cell_wire[210];							inform_R[217][5] = r_cell_wire[211];							inform_R[202][5] = r_cell_wire[212];							inform_R[218][5] = r_cell_wire[213];							inform_R[203][5] = r_cell_wire[214];							inform_R[219][5] = r_cell_wire[215];							inform_R[204][5] = r_cell_wire[216];							inform_R[220][5] = r_cell_wire[217];							inform_R[205][5] = r_cell_wire[218];							inform_R[221][5] = r_cell_wire[219];							inform_R[206][5] = r_cell_wire[220];							inform_R[222][5] = r_cell_wire[221];							inform_R[207][5] = r_cell_wire[222];							inform_R[223][5] = r_cell_wire[223];							inform_R[224][5] = r_cell_wire[224];							inform_R[240][5] = r_cell_wire[225];							inform_R[225][5] = r_cell_wire[226];							inform_R[241][5] = r_cell_wire[227];							inform_R[226][5] = r_cell_wire[228];							inform_R[242][5] = r_cell_wire[229];							inform_R[227][5] = r_cell_wire[230];							inform_R[243][5] = r_cell_wire[231];							inform_R[228][5] = r_cell_wire[232];							inform_R[244][5] = r_cell_wire[233];							inform_R[229][5] = r_cell_wire[234];							inform_R[245][5] = r_cell_wire[235];							inform_R[230][5] = r_cell_wire[236];							inform_R[246][5] = r_cell_wire[237];							inform_R[231][5] = r_cell_wire[238];							inform_R[247][5] = r_cell_wire[239];							inform_R[232][5] = r_cell_wire[240];							inform_R[248][5] = r_cell_wire[241];							inform_R[233][5] = r_cell_wire[242];							inform_R[249][5] = r_cell_wire[243];							inform_R[234][5] = r_cell_wire[244];							inform_R[250][5] = r_cell_wire[245];							inform_R[235][5] = r_cell_wire[246];							inform_R[251][5] = r_cell_wire[247];							inform_R[236][5] = r_cell_wire[248];							inform_R[252][5] = r_cell_wire[249];							inform_R[237][5] = r_cell_wire[250];							inform_R[253][5] = r_cell_wire[251];							inform_R[238][5] = r_cell_wire[252];							inform_R[254][5] = r_cell_wire[253];							inform_R[239][5] = r_cell_wire[254];							inform_R[255][5] = r_cell_wire[255];							inform_R[256][5] = r_cell_wire[256];							inform_R[272][5] = r_cell_wire[257];							inform_R[257][5] = r_cell_wire[258];							inform_R[273][5] = r_cell_wire[259];							inform_R[258][5] = r_cell_wire[260];							inform_R[274][5] = r_cell_wire[261];							inform_R[259][5] = r_cell_wire[262];							inform_R[275][5] = r_cell_wire[263];							inform_R[260][5] = r_cell_wire[264];							inform_R[276][5] = r_cell_wire[265];							inform_R[261][5] = r_cell_wire[266];							inform_R[277][5] = r_cell_wire[267];							inform_R[262][5] = r_cell_wire[268];							inform_R[278][5] = r_cell_wire[269];							inform_R[263][5] = r_cell_wire[270];							inform_R[279][5] = r_cell_wire[271];							inform_R[264][5] = r_cell_wire[272];							inform_R[280][5] = r_cell_wire[273];							inform_R[265][5] = r_cell_wire[274];							inform_R[281][5] = r_cell_wire[275];							inform_R[266][5] = r_cell_wire[276];							inform_R[282][5] = r_cell_wire[277];							inform_R[267][5] = r_cell_wire[278];							inform_R[283][5] = r_cell_wire[279];							inform_R[268][5] = r_cell_wire[280];							inform_R[284][5] = r_cell_wire[281];							inform_R[269][5] = r_cell_wire[282];							inform_R[285][5] = r_cell_wire[283];							inform_R[270][5] = r_cell_wire[284];							inform_R[286][5] = r_cell_wire[285];							inform_R[271][5] = r_cell_wire[286];							inform_R[287][5] = r_cell_wire[287];							inform_R[288][5] = r_cell_wire[288];							inform_R[304][5] = r_cell_wire[289];							inform_R[289][5] = r_cell_wire[290];							inform_R[305][5] = r_cell_wire[291];							inform_R[290][5] = r_cell_wire[292];							inform_R[306][5] = r_cell_wire[293];							inform_R[291][5] = r_cell_wire[294];							inform_R[307][5] = r_cell_wire[295];							inform_R[292][5] = r_cell_wire[296];							inform_R[308][5] = r_cell_wire[297];							inform_R[293][5] = r_cell_wire[298];							inform_R[309][5] = r_cell_wire[299];							inform_R[294][5] = r_cell_wire[300];							inform_R[310][5] = r_cell_wire[301];							inform_R[295][5] = r_cell_wire[302];							inform_R[311][5] = r_cell_wire[303];							inform_R[296][5] = r_cell_wire[304];							inform_R[312][5] = r_cell_wire[305];							inform_R[297][5] = r_cell_wire[306];							inform_R[313][5] = r_cell_wire[307];							inform_R[298][5] = r_cell_wire[308];							inform_R[314][5] = r_cell_wire[309];							inform_R[299][5] = r_cell_wire[310];							inform_R[315][5] = r_cell_wire[311];							inform_R[300][5] = r_cell_wire[312];							inform_R[316][5] = r_cell_wire[313];							inform_R[301][5] = r_cell_wire[314];							inform_R[317][5] = r_cell_wire[315];							inform_R[302][5] = r_cell_wire[316];							inform_R[318][5] = r_cell_wire[317];							inform_R[303][5] = r_cell_wire[318];							inform_R[319][5] = r_cell_wire[319];							inform_R[320][5] = r_cell_wire[320];							inform_R[336][5] = r_cell_wire[321];							inform_R[321][5] = r_cell_wire[322];							inform_R[337][5] = r_cell_wire[323];							inform_R[322][5] = r_cell_wire[324];							inform_R[338][5] = r_cell_wire[325];							inform_R[323][5] = r_cell_wire[326];							inform_R[339][5] = r_cell_wire[327];							inform_R[324][5] = r_cell_wire[328];							inform_R[340][5] = r_cell_wire[329];							inform_R[325][5] = r_cell_wire[330];							inform_R[341][5] = r_cell_wire[331];							inform_R[326][5] = r_cell_wire[332];							inform_R[342][5] = r_cell_wire[333];							inform_R[327][5] = r_cell_wire[334];							inform_R[343][5] = r_cell_wire[335];							inform_R[328][5] = r_cell_wire[336];							inform_R[344][5] = r_cell_wire[337];							inform_R[329][5] = r_cell_wire[338];							inform_R[345][5] = r_cell_wire[339];							inform_R[330][5] = r_cell_wire[340];							inform_R[346][5] = r_cell_wire[341];							inform_R[331][5] = r_cell_wire[342];							inform_R[347][5] = r_cell_wire[343];							inform_R[332][5] = r_cell_wire[344];							inform_R[348][5] = r_cell_wire[345];							inform_R[333][5] = r_cell_wire[346];							inform_R[349][5] = r_cell_wire[347];							inform_R[334][5] = r_cell_wire[348];							inform_R[350][5] = r_cell_wire[349];							inform_R[335][5] = r_cell_wire[350];							inform_R[351][5] = r_cell_wire[351];							inform_R[352][5] = r_cell_wire[352];							inform_R[368][5] = r_cell_wire[353];							inform_R[353][5] = r_cell_wire[354];							inform_R[369][5] = r_cell_wire[355];							inform_R[354][5] = r_cell_wire[356];							inform_R[370][5] = r_cell_wire[357];							inform_R[355][5] = r_cell_wire[358];							inform_R[371][5] = r_cell_wire[359];							inform_R[356][5] = r_cell_wire[360];							inform_R[372][5] = r_cell_wire[361];							inform_R[357][5] = r_cell_wire[362];							inform_R[373][5] = r_cell_wire[363];							inform_R[358][5] = r_cell_wire[364];							inform_R[374][5] = r_cell_wire[365];							inform_R[359][5] = r_cell_wire[366];							inform_R[375][5] = r_cell_wire[367];							inform_R[360][5] = r_cell_wire[368];							inform_R[376][5] = r_cell_wire[369];							inform_R[361][5] = r_cell_wire[370];							inform_R[377][5] = r_cell_wire[371];							inform_R[362][5] = r_cell_wire[372];							inform_R[378][5] = r_cell_wire[373];							inform_R[363][5] = r_cell_wire[374];							inform_R[379][5] = r_cell_wire[375];							inform_R[364][5] = r_cell_wire[376];							inform_R[380][5] = r_cell_wire[377];							inform_R[365][5] = r_cell_wire[378];							inform_R[381][5] = r_cell_wire[379];							inform_R[366][5] = r_cell_wire[380];							inform_R[382][5] = r_cell_wire[381];							inform_R[367][5] = r_cell_wire[382];							inform_R[383][5] = r_cell_wire[383];							inform_R[384][5] = r_cell_wire[384];							inform_R[400][5] = r_cell_wire[385];							inform_R[385][5] = r_cell_wire[386];							inform_R[401][5] = r_cell_wire[387];							inform_R[386][5] = r_cell_wire[388];							inform_R[402][5] = r_cell_wire[389];							inform_R[387][5] = r_cell_wire[390];							inform_R[403][5] = r_cell_wire[391];							inform_R[388][5] = r_cell_wire[392];							inform_R[404][5] = r_cell_wire[393];							inform_R[389][5] = r_cell_wire[394];							inform_R[405][5] = r_cell_wire[395];							inform_R[390][5] = r_cell_wire[396];							inform_R[406][5] = r_cell_wire[397];							inform_R[391][5] = r_cell_wire[398];							inform_R[407][5] = r_cell_wire[399];							inform_R[392][5] = r_cell_wire[400];							inform_R[408][5] = r_cell_wire[401];							inform_R[393][5] = r_cell_wire[402];							inform_R[409][5] = r_cell_wire[403];							inform_R[394][5] = r_cell_wire[404];							inform_R[410][5] = r_cell_wire[405];							inform_R[395][5] = r_cell_wire[406];							inform_R[411][5] = r_cell_wire[407];							inform_R[396][5] = r_cell_wire[408];							inform_R[412][5] = r_cell_wire[409];							inform_R[397][5] = r_cell_wire[410];							inform_R[413][5] = r_cell_wire[411];							inform_R[398][5] = r_cell_wire[412];							inform_R[414][5] = r_cell_wire[413];							inform_R[399][5] = r_cell_wire[414];							inform_R[415][5] = r_cell_wire[415];							inform_R[416][5] = r_cell_wire[416];							inform_R[432][5] = r_cell_wire[417];							inform_R[417][5] = r_cell_wire[418];							inform_R[433][5] = r_cell_wire[419];							inform_R[418][5] = r_cell_wire[420];							inform_R[434][5] = r_cell_wire[421];							inform_R[419][5] = r_cell_wire[422];							inform_R[435][5] = r_cell_wire[423];							inform_R[420][5] = r_cell_wire[424];							inform_R[436][5] = r_cell_wire[425];							inform_R[421][5] = r_cell_wire[426];							inform_R[437][5] = r_cell_wire[427];							inform_R[422][5] = r_cell_wire[428];							inform_R[438][5] = r_cell_wire[429];							inform_R[423][5] = r_cell_wire[430];							inform_R[439][5] = r_cell_wire[431];							inform_R[424][5] = r_cell_wire[432];							inform_R[440][5] = r_cell_wire[433];							inform_R[425][5] = r_cell_wire[434];							inform_R[441][5] = r_cell_wire[435];							inform_R[426][5] = r_cell_wire[436];							inform_R[442][5] = r_cell_wire[437];							inform_R[427][5] = r_cell_wire[438];							inform_R[443][5] = r_cell_wire[439];							inform_R[428][5] = r_cell_wire[440];							inform_R[444][5] = r_cell_wire[441];							inform_R[429][5] = r_cell_wire[442];							inform_R[445][5] = r_cell_wire[443];							inform_R[430][5] = r_cell_wire[444];							inform_R[446][5] = r_cell_wire[445];							inform_R[431][5] = r_cell_wire[446];							inform_R[447][5] = r_cell_wire[447];							inform_R[448][5] = r_cell_wire[448];							inform_R[464][5] = r_cell_wire[449];							inform_R[449][5] = r_cell_wire[450];							inform_R[465][5] = r_cell_wire[451];							inform_R[450][5] = r_cell_wire[452];							inform_R[466][5] = r_cell_wire[453];							inform_R[451][5] = r_cell_wire[454];							inform_R[467][5] = r_cell_wire[455];							inform_R[452][5] = r_cell_wire[456];							inform_R[468][5] = r_cell_wire[457];							inform_R[453][5] = r_cell_wire[458];							inform_R[469][5] = r_cell_wire[459];							inform_R[454][5] = r_cell_wire[460];							inform_R[470][5] = r_cell_wire[461];							inform_R[455][5] = r_cell_wire[462];							inform_R[471][5] = r_cell_wire[463];							inform_R[456][5] = r_cell_wire[464];							inform_R[472][5] = r_cell_wire[465];							inform_R[457][5] = r_cell_wire[466];							inform_R[473][5] = r_cell_wire[467];							inform_R[458][5] = r_cell_wire[468];							inform_R[474][5] = r_cell_wire[469];							inform_R[459][5] = r_cell_wire[470];							inform_R[475][5] = r_cell_wire[471];							inform_R[460][5] = r_cell_wire[472];							inform_R[476][5] = r_cell_wire[473];							inform_R[461][5] = r_cell_wire[474];							inform_R[477][5] = r_cell_wire[475];							inform_R[462][5] = r_cell_wire[476];							inform_R[478][5] = r_cell_wire[477];							inform_R[463][5] = r_cell_wire[478];							inform_R[479][5] = r_cell_wire[479];							inform_R[480][5] = r_cell_wire[480];							inform_R[496][5] = r_cell_wire[481];							inform_R[481][5] = r_cell_wire[482];							inform_R[497][5] = r_cell_wire[483];							inform_R[482][5] = r_cell_wire[484];							inform_R[498][5] = r_cell_wire[485];							inform_R[483][5] = r_cell_wire[486];							inform_R[499][5] = r_cell_wire[487];							inform_R[484][5] = r_cell_wire[488];							inform_R[500][5] = r_cell_wire[489];							inform_R[485][5] = r_cell_wire[490];							inform_R[501][5] = r_cell_wire[491];							inform_R[486][5] = r_cell_wire[492];							inform_R[502][5] = r_cell_wire[493];							inform_R[487][5] = r_cell_wire[494];							inform_R[503][5] = r_cell_wire[495];							inform_R[488][5] = r_cell_wire[496];							inform_R[504][5] = r_cell_wire[497];							inform_R[489][5] = r_cell_wire[498];							inform_R[505][5] = r_cell_wire[499];							inform_R[490][5] = r_cell_wire[500];							inform_R[506][5] = r_cell_wire[501];							inform_R[491][5] = r_cell_wire[502];							inform_R[507][5] = r_cell_wire[503];							inform_R[492][5] = r_cell_wire[504];							inform_R[508][5] = r_cell_wire[505];							inform_R[493][5] = r_cell_wire[506];							inform_R[509][5] = r_cell_wire[507];							inform_R[494][5] = r_cell_wire[508];							inform_R[510][5] = r_cell_wire[509];							inform_R[495][5] = r_cell_wire[510];							inform_R[511][5] = r_cell_wire[511];							inform_R[512][5] = r_cell_wire[512];							inform_R[528][5] = r_cell_wire[513];							inform_R[513][5] = r_cell_wire[514];							inform_R[529][5] = r_cell_wire[515];							inform_R[514][5] = r_cell_wire[516];							inform_R[530][5] = r_cell_wire[517];							inform_R[515][5] = r_cell_wire[518];							inform_R[531][5] = r_cell_wire[519];							inform_R[516][5] = r_cell_wire[520];							inform_R[532][5] = r_cell_wire[521];							inform_R[517][5] = r_cell_wire[522];							inform_R[533][5] = r_cell_wire[523];							inform_R[518][5] = r_cell_wire[524];							inform_R[534][5] = r_cell_wire[525];							inform_R[519][5] = r_cell_wire[526];							inform_R[535][5] = r_cell_wire[527];							inform_R[520][5] = r_cell_wire[528];							inform_R[536][5] = r_cell_wire[529];							inform_R[521][5] = r_cell_wire[530];							inform_R[537][5] = r_cell_wire[531];							inform_R[522][5] = r_cell_wire[532];							inform_R[538][5] = r_cell_wire[533];							inform_R[523][5] = r_cell_wire[534];							inform_R[539][5] = r_cell_wire[535];							inform_R[524][5] = r_cell_wire[536];							inform_R[540][5] = r_cell_wire[537];							inform_R[525][5] = r_cell_wire[538];							inform_R[541][5] = r_cell_wire[539];							inform_R[526][5] = r_cell_wire[540];							inform_R[542][5] = r_cell_wire[541];							inform_R[527][5] = r_cell_wire[542];							inform_R[543][5] = r_cell_wire[543];							inform_R[544][5] = r_cell_wire[544];							inform_R[560][5] = r_cell_wire[545];							inform_R[545][5] = r_cell_wire[546];							inform_R[561][5] = r_cell_wire[547];							inform_R[546][5] = r_cell_wire[548];							inform_R[562][5] = r_cell_wire[549];							inform_R[547][5] = r_cell_wire[550];							inform_R[563][5] = r_cell_wire[551];							inform_R[548][5] = r_cell_wire[552];							inform_R[564][5] = r_cell_wire[553];							inform_R[549][5] = r_cell_wire[554];							inform_R[565][5] = r_cell_wire[555];							inform_R[550][5] = r_cell_wire[556];							inform_R[566][5] = r_cell_wire[557];							inform_R[551][5] = r_cell_wire[558];							inform_R[567][5] = r_cell_wire[559];							inform_R[552][5] = r_cell_wire[560];							inform_R[568][5] = r_cell_wire[561];							inform_R[553][5] = r_cell_wire[562];							inform_R[569][5] = r_cell_wire[563];							inform_R[554][5] = r_cell_wire[564];							inform_R[570][5] = r_cell_wire[565];							inform_R[555][5] = r_cell_wire[566];							inform_R[571][5] = r_cell_wire[567];							inform_R[556][5] = r_cell_wire[568];							inform_R[572][5] = r_cell_wire[569];							inform_R[557][5] = r_cell_wire[570];							inform_R[573][5] = r_cell_wire[571];							inform_R[558][5] = r_cell_wire[572];							inform_R[574][5] = r_cell_wire[573];							inform_R[559][5] = r_cell_wire[574];							inform_R[575][5] = r_cell_wire[575];							inform_R[576][5] = r_cell_wire[576];							inform_R[592][5] = r_cell_wire[577];							inform_R[577][5] = r_cell_wire[578];							inform_R[593][5] = r_cell_wire[579];							inform_R[578][5] = r_cell_wire[580];							inform_R[594][5] = r_cell_wire[581];							inform_R[579][5] = r_cell_wire[582];							inform_R[595][5] = r_cell_wire[583];							inform_R[580][5] = r_cell_wire[584];							inform_R[596][5] = r_cell_wire[585];							inform_R[581][5] = r_cell_wire[586];							inform_R[597][5] = r_cell_wire[587];							inform_R[582][5] = r_cell_wire[588];							inform_R[598][5] = r_cell_wire[589];							inform_R[583][5] = r_cell_wire[590];							inform_R[599][5] = r_cell_wire[591];							inform_R[584][5] = r_cell_wire[592];							inform_R[600][5] = r_cell_wire[593];							inform_R[585][5] = r_cell_wire[594];							inform_R[601][5] = r_cell_wire[595];							inform_R[586][5] = r_cell_wire[596];							inform_R[602][5] = r_cell_wire[597];							inform_R[587][5] = r_cell_wire[598];							inform_R[603][5] = r_cell_wire[599];							inform_R[588][5] = r_cell_wire[600];							inform_R[604][5] = r_cell_wire[601];							inform_R[589][5] = r_cell_wire[602];							inform_R[605][5] = r_cell_wire[603];							inform_R[590][5] = r_cell_wire[604];							inform_R[606][5] = r_cell_wire[605];							inform_R[591][5] = r_cell_wire[606];							inform_R[607][5] = r_cell_wire[607];							inform_R[608][5] = r_cell_wire[608];							inform_R[624][5] = r_cell_wire[609];							inform_R[609][5] = r_cell_wire[610];							inform_R[625][5] = r_cell_wire[611];							inform_R[610][5] = r_cell_wire[612];							inform_R[626][5] = r_cell_wire[613];							inform_R[611][5] = r_cell_wire[614];							inform_R[627][5] = r_cell_wire[615];							inform_R[612][5] = r_cell_wire[616];							inform_R[628][5] = r_cell_wire[617];							inform_R[613][5] = r_cell_wire[618];							inform_R[629][5] = r_cell_wire[619];							inform_R[614][5] = r_cell_wire[620];							inform_R[630][5] = r_cell_wire[621];							inform_R[615][5] = r_cell_wire[622];							inform_R[631][5] = r_cell_wire[623];							inform_R[616][5] = r_cell_wire[624];							inform_R[632][5] = r_cell_wire[625];							inform_R[617][5] = r_cell_wire[626];							inform_R[633][5] = r_cell_wire[627];							inform_R[618][5] = r_cell_wire[628];							inform_R[634][5] = r_cell_wire[629];							inform_R[619][5] = r_cell_wire[630];							inform_R[635][5] = r_cell_wire[631];							inform_R[620][5] = r_cell_wire[632];							inform_R[636][5] = r_cell_wire[633];							inform_R[621][5] = r_cell_wire[634];							inform_R[637][5] = r_cell_wire[635];							inform_R[622][5] = r_cell_wire[636];							inform_R[638][5] = r_cell_wire[637];							inform_R[623][5] = r_cell_wire[638];							inform_R[639][5] = r_cell_wire[639];							inform_R[640][5] = r_cell_wire[640];							inform_R[656][5] = r_cell_wire[641];							inform_R[641][5] = r_cell_wire[642];							inform_R[657][5] = r_cell_wire[643];							inform_R[642][5] = r_cell_wire[644];							inform_R[658][5] = r_cell_wire[645];							inform_R[643][5] = r_cell_wire[646];							inform_R[659][5] = r_cell_wire[647];							inform_R[644][5] = r_cell_wire[648];							inform_R[660][5] = r_cell_wire[649];							inform_R[645][5] = r_cell_wire[650];							inform_R[661][5] = r_cell_wire[651];							inform_R[646][5] = r_cell_wire[652];							inform_R[662][5] = r_cell_wire[653];							inform_R[647][5] = r_cell_wire[654];							inform_R[663][5] = r_cell_wire[655];							inform_R[648][5] = r_cell_wire[656];							inform_R[664][5] = r_cell_wire[657];							inform_R[649][5] = r_cell_wire[658];							inform_R[665][5] = r_cell_wire[659];							inform_R[650][5] = r_cell_wire[660];							inform_R[666][5] = r_cell_wire[661];							inform_R[651][5] = r_cell_wire[662];							inform_R[667][5] = r_cell_wire[663];							inform_R[652][5] = r_cell_wire[664];							inform_R[668][5] = r_cell_wire[665];							inform_R[653][5] = r_cell_wire[666];							inform_R[669][5] = r_cell_wire[667];							inform_R[654][5] = r_cell_wire[668];							inform_R[670][5] = r_cell_wire[669];							inform_R[655][5] = r_cell_wire[670];							inform_R[671][5] = r_cell_wire[671];							inform_R[672][5] = r_cell_wire[672];							inform_R[688][5] = r_cell_wire[673];							inform_R[673][5] = r_cell_wire[674];							inform_R[689][5] = r_cell_wire[675];							inform_R[674][5] = r_cell_wire[676];							inform_R[690][5] = r_cell_wire[677];							inform_R[675][5] = r_cell_wire[678];							inform_R[691][5] = r_cell_wire[679];							inform_R[676][5] = r_cell_wire[680];							inform_R[692][5] = r_cell_wire[681];							inform_R[677][5] = r_cell_wire[682];							inform_R[693][5] = r_cell_wire[683];							inform_R[678][5] = r_cell_wire[684];							inform_R[694][5] = r_cell_wire[685];							inform_R[679][5] = r_cell_wire[686];							inform_R[695][5] = r_cell_wire[687];							inform_R[680][5] = r_cell_wire[688];							inform_R[696][5] = r_cell_wire[689];							inform_R[681][5] = r_cell_wire[690];							inform_R[697][5] = r_cell_wire[691];							inform_R[682][5] = r_cell_wire[692];							inform_R[698][5] = r_cell_wire[693];							inform_R[683][5] = r_cell_wire[694];							inform_R[699][5] = r_cell_wire[695];							inform_R[684][5] = r_cell_wire[696];							inform_R[700][5] = r_cell_wire[697];							inform_R[685][5] = r_cell_wire[698];							inform_R[701][5] = r_cell_wire[699];							inform_R[686][5] = r_cell_wire[700];							inform_R[702][5] = r_cell_wire[701];							inform_R[687][5] = r_cell_wire[702];							inform_R[703][5] = r_cell_wire[703];							inform_R[704][5] = r_cell_wire[704];							inform_R[720][5] = r_cell_wire[705];							inform_R[705][5] = r_cell_wire[706];							inform_R[721][5] = r_cell_wire[707];							inform_R[706][5] = r_cell_wire[708];							inform_R[722][5] = r_cell_wire[709];							inform_R[707][5] = r_cell_wire[710];							inform_R[723][5] = r_cell_wire[711];							inform_R[708][5] = r_cell_wire[712];							inform_R[724][5] = r_cell_wire[713];							inform_R[709][5] = r_cell_wire[714];							inform_R[725][5] = r_cell_wire[715];							inform_R[710][5] = r_cell_wire[716];							inform_R[726][5] = r_cell_wire[717];							inform_R[711][5] = r_cell_wire[718];							inform_R[727][5] = r_cell_wire[719];							inform_R[712][5] = r_cell_wire[720];							inform_R[728][5] = r_cell_wire[721];							inform_R[713][5] = r_cell_wire[722];							inform_R[729][5] = r_cell_wire[723];							inform_R[714][5] = r_cell_wire[724];							inform_R[730][5] = r_cell_wire[725];							inform_R[715][5] = r_cell_wire[726];							inform_R[731][5] = r_cell_wire[727];							inform_R[716][5] = r_cell_wire[728];							inform_R[732][5] = r_cell_wire[729];							inform_R[717][5] = r_cell_wire[730];							inform_R[733][5] = r_cell_wire[731];							inform_R[718][5] = r_cell_wire[732];							inform_R[734][5] = r_cell_wire[733];							inform_R[719][5] = r_cell_wire[734];							inform_R[735][5] = r_cell_wire[735];							inform_R[736][5] = r_cell_wire[736];							inform_R[752][5] = r_cell_wire[737];							inform_R[737][5] = r_cell_wire[738];							inform_R[753][5] = r_cell_wire[739];							inform_R[738][5] = r_cell_wire[740];							inform_R[754][5] = r_cell_wire[741];							inform_R[739][5] = r_cell_wire[742];							inform_R[755][5] = r_cell_wire[743];							inform_R[740][5] = r_cell_wire[744];							inform_R[756][5] = r_cell_wire[745];							inform_R[741][5] = r_cell_wire[746];							inform_R[757][5] = r_cell_wire[747];							inform_R[742][5] = r_cell_wire[748];							inform_R[758][5] = r_cell_wire[749];							inform_R[743][5] = r_cell_wire[750];							inform_R[759][5] = r_cell_wire[751];							inform_R[744][5] = r_cell_wire[752];							inform_R[760][5] = r_cell_wire[753];							inform_R[745][5] = r_cell_wire[754];							inform_R[761][5] = r_cell_wire[755];							inform_R[746][5] = r_cell_wire[756];							inform_R[762][5] = r_cell_wire[757];							inform_R[747][5] = r_cell_wire[758];							inform_R[763][5] = r_cell_wire[759];							inform_R[748][5] = r_cell_wire[760];							inform_R[764][5] = r_cell_wire[761];							inform_R[749][5] = r_cell_wire[762];							inform_R[765][5] = r_cell_wire[763];							inform_R[750][5] = r_cell_wire[764];							inform_R[766][5] = r_cell_wire[765];							inform_R[751][5] = r_cell_wire[766];							inform_R[767][5] = r_cell_wire[767];							inform_R[768][5] = r_cell_wire[768];							inform_R[784][5] = r_cell_wire[769];							inform_R[769][5] = r_cell_wire[770];							inform_R[785][5] = r_cell_wire[771];							inform_R[770][5] = r_cell_wire[772];							inform_R[786][5] = r_cell_wire[773];							inform_R[771][5] = r_cell_wire[774];							inform_R[787][5] = r_cell_wire[775];							inform_R[772][5] = r_cell_wire[776];							inform_R[788][5] = r_cell_wire[777];							inform_R[773][5] = r_cell_wire[778];							inform_R[789][5] = r_cell_wire[779];							inform_R[774][5] = r_cell_wire[780];							inform_R[790][5] = r_cell_wire[781];							inform_R[775][5] = r_cell_wire[782];							inform_R[791][5] = r_cell_wire[783];							inform_R[776][5] = r_cell_wire[784];							inform_R[792][5] = r_cell_wire[785];							inform_R[777][5] = r_cell_wire[786];							inform_R[793][5] = r_cell_wire[787];							inform_R[778][5] = r_cell_wire[788];							inform_R[794][5] = r_cell_wire[789];							inform_R[779][5] = r_cell_wire[790];							inform_R[795][5] = r_cell_wire[791];							inform_R[780][5] = r_cell_wire[792];							inform_R[796][5] = r_cell_wire[793];							inform_R[781][5] = r_cell_wire[794];							inform_R[797][5] = r_cell_wire[795];							inform_R[782][5] = r_cell_wire[796];							inform_R[798][5] = r_cell_wire[797];							inform_R[783][5] = r_cell_wire[798];							inform_R[799][5] = r_cell_wire[799];							inform_R[800][5] = r_cell_wire[800];							inform_R[816][5] = r_cell_wire[801];							inform_R[801][5] = r_cell_wire[802];							inform_R[817][5] = r_cell_wire[803];							inform_R[802][5] = r_cell_wire[804];							inform_R[818][5] = r_cell_wire[805];							inform_R[803][5] = r_cell_wire[806];							inform_R[819][5] = r_cell_wire[807];							inform_R[804][5] = r_cell_wire[808];							inform_R[820][5] = r_cell_wire[809];							inform_R[805][5] = r_cell_wire[810];							inform_R[821][5] = r_cell_wire[811];							inform_R[806][5] = r_cell_wire[812];							inform_R[822][5] = r_cell_wire[813];							inform_R[807][5] = r_cell_wire[814];							inform_R[823][5] = r_cell_wire[815];							inform_R[808][5] = r_cell_wire[816];							inform_R[824][5] = r_cell_wire[817];							inform_R[809][5] = r_cell_wire[818];							inform_R[825][5] = r_cell_wire[819];							inform_R[810][5] = r_cell_wire[820];							inform_R[826][5] = r_cell_wire[821];							inform_R[811][5] = r_cell_wire[822];							inform_R[827][5] = r_cell_wire[823];							inform_R[812][5] = r_cell_wire[824];							inform_R[828][5] = r_cell_wire[825];							inform_R[813][5] = r_cell_wire[826];							inform_R[829][5] = r_cell_wire[827];							inform_R[814][5] = r_cell_wire[828];							inform_R[830][5] = r_cell_wire[829];							inform_R[815][5] = r_cell_wire[830];							inform_R[831][5] = r_cell_wire[831];							inform_R[832][5] = r_cell_wire[832];							inform_R[848][5] = r_cell_wire[833];							inform_R[833][5] = r_cell_wire[834];							inform_R[849][5] = r_cell_wire[835];							inform_R[834][5] = r_cell_wire[836];							inform_R[850][5] = r_cell_wire[837];							inform_R[835][5] = r_cell_wire[838];							inform_R[851][5] = r_cell_wire[839];							inform_R[836][5] = r_cell_wire[840];							inform_R[852][5] = r_cell_wire[841];							inform_R[837][5] = r_cell_wire[842];							inform_R[853][5] = r_cell_wire[843];							inform_R[838][5] = r_cell_wire[844];							inform_R[854][5] = r_cell_wire[845];							inform_R[839][5] = r_cell_wire[846];							inform_R[855][5] = r_cell_wire[847];							inform_R[840][5] = r_cell_wire[848];							inform_R[856][5] = r_cell_wire[849];							inform_R[841][5] = r_cell_wire[850];							inform_R[857][5] = r_cell_wire[851];							inform_R[842][5] = r_cell_wire[852];							inform_R[858][5] = r_cell_wire[853];							inform_R[843][5] = r_cell_wire[854];							inform_R[859][5] = r_cell_wire[855];							inform_R[844][5] = r_cell_wire[856];							inform_R[860][5] = r_cell_wire[857];							inform_R[845][5] = r_cell_wire[858];							inform_R[861][5] = r_cell_wire[859];							inform_R[846][5] = r_cell_wire[860];							inform_R[862][5] = r_cell_wire[861];							inform_R[847][5] = r_cell_wire[862];							inform_R[863][5] = r_cell_wire[863];							inform_R[864][5] = r_cell_wire[864];							inform_R[880][5] = r_cell_wire[865];							inform_R[865][5] = r_cell_wire[866];							inform_R[881][5] = r_cell_wire[867];							inform_R[866][5] = r_cell_wire[868];							inform_R[882][5] = r_cell_wire[869];							inform_R[867][5] = r_cell_wire[870];							inform_R[883][5] = r_cell_wire[871];							inform_R[868][5] = r_cell_wire[872];							inform_R[884][5] = r_cell_wire[873];							inform_R[869][5] = r_cell_wire[874];							inform_R[885][5] = r_cell_wire[875];							inform_R[870][5] = r_cell_wire[876];							inform_R[886][5] = r_cell_wire[877];							inform_R[871][5] = r_cell_wire[878];							inform_R[887][5] = r_cell_wire[879];							inform_R[872][5] = r_cell_wire[880];							inform_R[888][5] = r_cell_wire[881];							inform_R[873][5] = r_cell_wire[882];							inform_R[889][5] = r_cell_wire[883];							inform_R[874][5] = r_cell_wire[884];							inform_R[890][5] = r_cell_wire[885];							inform_R[875][5] = r_cell_wire[886];							inform_R[891][5] = r_cell_wire[887];							inform_R[876][5] = r_cell_wire[888];							inform_R[892][5] = r_cell_wire[889];							inform_R[877][5] = r_cell_wire[890];							inform_R[893][5] = r_cell_wire[891];							inform_R[878][5] = r_cell_wire[892];							inform_R[894][5] = r_cell_wire[893];							inform_R[879][5] = r_cell_wire[894];							inform_R[895][5] = r_cell_wire[895];							inform_R[896][5] = r_cell_wire[896];							inform_R[912][5] = r_cell_wire[897];							inform_R[897][5] = r_cell_wire[898];							inform_R[913][5] = r_cell_wire[899];							inform_R[898][5] = r_cell_wire[900];							inform_R[914][5] = r_cell_wire[901];							inform_R[899][5] = r_cell_wire[902];							inform_R[915][5] = r_cell_wire[903];							inform_R[900][5] = r_cell_wire[904];							inform_R[916][5] = r_cell_wire[905];							inform_R[901][5] = r_cell_wire[906];							inform_R[917][5] = r_cell_wire[907];							inform_R[902][5] = r_cell_wire[908];							inform_R[918][5] = r_cell_wire[909];							inform_R[903][5] = r_cell_wire[910];							inform_R[919][5] = r_cell_wire[911];							inform_R[904][5] = r_cell_wire[912];							inform_R[920][5] = r_cell_wire[913];							inform_R[905][5] = r_cell_wire[914];							inform_R[921][5] = r_cell_wire[915];							inform_R[906][5] = r_cell_wire[916];							inform_R[922][5] = r_cell_wire[917];							inform_R[907][5] = r_cell_wire[918];							inform_R[923][5] = r_cell_wire[919];							inform_R[908][5] = r_cell_wire[920];							inform_R[924][5] = r_cell_wire[921];							inform_R[909][5] = r_cell_wire[922];							inform_R[925][5] = r_cell_wire[923];							inform_R[910][5] = r_cell_wire[924];							inform_R[926][5] = r_cell_wire[925];							inform_R[911][5] = r_cell_wire[926];							inform_R[927][5] = r_cell_wire[927];							inform_R[928][5] = r_cell_wire[928];							inform_R[944][5] = r_cell_wire[929];							inform_R[929][5] = r_cell_wire[930];							inform_R[945][5] = r_cell_wire[931];							inform_R[930][5] = r_cell_wire[932];							inform_R[946][5] = r_cell_wire[933];							inform_R[931][5] = r_cell_wire[934];							inform_R[947][5] = r_cell_wire[935];							inform_R[932][5] = r_cell_wire[936];							inform_R[948][5] = r_cell_wire[937];							inform_R[933][5] = r_cell_wire[938];							inform_R[949][5] = r_cell_wire[939];							inform_R[934][5] = r_cell_wire[940];							inform_R[950][5] = r_cell_wire[941];							inform_R[935][5] = r_cell_wire[942];							inform_R[951][5] = r_cell_wire[943];							inform_R[936][5] = r_cell_wire[944];							inform_R[952][5] = r_cell_wire[945];							inform_R[937][5] = r_cell_wire[946];							inform_R[953][5] = r_cell_wire[947];							inform_R[938][5] = r_cell_wire[948];							inform_R[954][5] = r_cell_wire[949];							inform_R[939][5] = r_cell_wire[950];							inform_R[955][5] = r_cell_wire[951];							inform_R[940][5] = r_cell_wire[952];							inform_R[956][5] = r_cell_wire[953];							inform_R[941][5] = r_cell_wire[954];							inform_R[957][5] = r_cell_wire[955];							inform_R[942][5] = r_cell_wire[956];							inform_R[958][5] = r_cell_wire[957];							inform_R[943][5] = r_cell_wire[958];							inform_R[959][5] = r_cell_wire[959];							inform_R[960][5] = r_cell_wire[960];							inform_R[976][5] = r_cell_wire[961];							inform_R[961][5] = r_cell_wire[962];							inform_R[977][5] = r_cell_wire[963];							inform_R[962][5] = r_cell_wire[964];							inform_R[978][5] = r_cell_wire[965];							inform_R[963][5] = r_cell_wire[966];							inform_R[979][5] = r_cell_wire[967];							inform_R[964][5] = r_cell_wire[968];							inform_R[980][5] = r_cell_wire[969];							inform_R[965][5] = r_cell_wire[970];							inform_R[981][5] = r_cell_wire[971];							inform_R[966][5] = r_cell_wire[972];							inform_R[982][5] = r_cell_wire[973];							inform_R[967][5] = r_cell_wire[974];							inform_R[983][5] = r_cell_wire[975];							inform_R[968][5] = r_cell_wire[976];							inform_R[984][5] = r_cell_wire[977];							inform_R[969][5] = r_cell_wire[978];							inform_R[985][5] = r_cell_wire[979];							inform_R[970][5] = r_cell_wire[980];							inform_R[986][5] = r_cell_wire[981];							inform_R[971][5] = r_cell_wire[982];							inform_R[987][5] = r_cell_wire[983];							inform_R[972][5] = r_cell_wire[984];							inform_R[988][5] = r_cell_wire[985];							inform_R[973][5] = r_cell_wire[986];							inform_R[989][5] = r_cell_wire[987];							inform_R[974][5] = r_cell_wire[988];							inform_R[990][5] = r_cell_wire[989];							inform_R[975][5] = r_cell_wire[990];							inform_R[991][5] = r_cell_wire[991];							inform_R[992][5] = r_cell_wire[992];							inform_R[1008][5] = r_cell_wire[993];							inform_R[993][5] = r_cell_wire[994];							inform_R[1009][5] = r_cell_wire[995];							inform_R[994][5] = r_cell_wire[996];							inform_R[1010][5] = r_cell_wire[997];							inform_R[995][5] = r_cell_wire[998];							inform_R[1011][5] = r_cell_wire[999];							inform_R[996][5] = r_cell_wire[1000];							inform_R[1012][5] = r_cell_wire[1001];							inform_R[997][5] = r_cell_wire[1002];							inform_R[1013][5] = r_cell_wire[1003];							inform_R[998][5] = r_cell_wire[1004];							inform_R[1014][5] = r_cell_wire[1005];							inform_R[999][5] = r_cell_wire[1006];							inform_R[1015][5] = r_cell_wire[1007];							inform_R[1000][5] = r_cell_wire[1008];							inform_R[1016][5] = r_cell_wire[1009];							inform_R[1001][5] = r_cell_wire[1010];							inform_R[1017][5] = r_cell_wire[1011];							inform_R[1002][5] = r_cell_wire[1012];							inform_R[1018][5] = r_cell_wire[1013];							inform_R[1003][5] = r_cell_wire[1014];							inform_R[1019][5] = r_cell_wire[1015];							inform_R[1004][5] = r_cell_wire[1016];							inform_R[1020][5] = r_cell_wire[1017];							inform_R[1005][5] = r_cell_wire[1018];							inform_R[1021][5] = r_cell_wire[1019];							inform_R[1006][5] = r_cell_wire[1020];							inform_R[1022][5] = r_cell_wire[1021];							inform_R[1007][5] = r_cell_wire[1022];							inform_R[1023][5] = r_cell_wire[1023];							inform_L[0][4] = l_cell_wire[0];							inform_L[16][4] = l_cell_wire[1];							inform_L[1][4] = l_cell_wire[2];							inform_L[17][4] = l_cell_wire[3];							inform_L[2][4] = l_cell_wire[4];							inform_L[18][4] = l_cell_wire[5];							inform_L[3][4] = l_cell_wire[6];							inform_L[19][4] = l_cell_wire[7];							inform_L[4][4] = l_cell_wire[8];							inform_L[20][4] = l_cell_wire[9];							inform_L[5][4] = l_cell_wire[10];							inform_L[21][4] = l_cell_wire[11];							inform_L[6][4] = l_cell_wire[12];							inform_L[22][4] = l_cell_wire[13];							inform_L[7][4] = l_cell_wire[14];							inform_L[23][4] = l_cell_wire[15];							inform_L[8][4] = l_cell_wire[16];							inform_L[24][4] = l_cell_wire[17];							inform_L[9][4] = l_cell_wire[18];							inform_L[25][4] = l_cell_wire[19];							inform_L[10][4] = l_cell_wire[20];							inform_L[26][4] = l_cell_wire[21];							inform_L[11][4] = l_cell_wire[22];							inform_L[27][4] = l_cell_wire[23];							inform_L[12][4] = l_cell_wire[24];							inform_L[28][4] = l_cell_wire[25];							inform_L[13][4] = l_cell_wire[26];							inform_L[29][4] = l_cell_wire[27];							inform_L[14][4] = l_cell_wire[28];							inform_L[30][4] = l_cell_wire[29];							inform_L[15][4] = l_cell_wire[30];							inform_L[31][4] = l_cell_wire[31];							inform_L[32][4] = l_cell_wire[32];							inform_L[48][4] = l_cell_wire[33];							inform_L[33][4] = l_cell_wire[34];							inform_L[49][4] = l_cell_wire[35];							inform_L[34][4] = l_cell_wire[36];							inform_L[50][4] = l_cell_wire[37];							inform_L[35][4] = l_cell_wire[38];							inform_L[51][4] = l_cell_wire[39];							inform_L[36][4] = l_cell_wire[40];							inform_L[52][4] = l_cell_wire[41];							inform_L[37][4] = l_cell_wire[42];							inform_L[53][4] = l_cell_wire[43];							inform_L[38][4] = l_cell_wire[44];							inform_L[54][4] = l_cell_wire[45];							inform_L[39][4] = l_cell_wire[46];							inform_L[55][4] = l_cell_wire[47];							inform_L[40][4] = l_cell_wire[48];							inform_L[56][4] = l_cell_wire[49];							inform_L[41][4] = l_cell_wire[50];							inform_L[57][4] = l_cell_wire[51];							inform_L[42][4] = l_cell_wire[52];							inform_L[58][4] = l_cell_wire[53];							inform_L[43][4] = l_cell_wire[54];							inform_L[59][4] = l_cell_wire[55];							inform_L[44][4] = l_cell_wire[56];							inform_L[60][4] = l_cell_wire[57];							inform_L[45][4] = l_cell_wire[58];							inform_L[61][4] = l_cell_wire[59];							inform_L[46][4] = l_cell_wire[60];							inform_L[62][4] = l_cell_wire[61];							inform_L[47][4] = l_cell_wire[62];							inform_L[63][4] = l_cell_wire[63];							inform_L[64][4] = l_cell_wire[64];							inform_L[80][4] = l_cell_wire[65];							inform_L[65][4] = l_cell_wire[66];							inform_L[81][4] = l_cell_wire[67];							inform_L[66][4] = l_cell_wire[68];							inform_L[82][4] = l_cell_wire[69];							inform_L[67][4] = l_cell_wire[70];							inform_L[83][4] = l_cell_wire[71];							inform_L[68][4] = l_cell_wire[72];							inform_L[84][4] = l_cell_wire[73];							inform_L[69][4] = l_cell_wire[74];							inform_L[85][4] = l_cell_wire[75];							inform_L[70][4] = l_cell_wire[76];							inform_L[86][4] = l_cell_wire[77];							inform_L[71][4] = l_cell_wire[78];							inform_L[87][4] = l_cell_wire[79];							inform_L[72][4] = l_cell_wire[80];							inform_L[88][4] = l_cell_wire[81];							inform_L[73][4] = l_cell_wire[82];							inform_L[89][4] = l_cell_wire[83];							inform_L[74][4] = l_cell_wire[84];							inform_L[90][4] = l_cell_wire[85];							inform_L[75][4] = l_cell_wire[86];							inform_L[91][4] = l_cell_wire[87];							inform_L[76][4] = l_cell_wire[88];							inform_L[92][4] = l_cell_wire[89];							inform_L[77][4] = l_cell_wire[90];							inform_L[93][4] = l_cell_wire[91];							inform_L[78][4] = l_cell_wire[92];							inform_L[94][4] = l_cell_wire[93];							inform_L[79][4] = l_cell_wire[94];							inform_L[95][4] = l_cell_wire[95];							inform_L[96][4] = l_cell_wire[96];							inform_L[112][4] = l_cell_wire[97];							inform_L[97][4] = l_cell_wire[98];							inform_L[113][4] = l_cell_wire[99];							inform_L[98][4] = l_cell_wire[100];							inform_L[114][4] = l_cell_wire[101];							inform_L[99][4] = l_cell_wire[102];							inform_L[115][4] = l_cell_wire[103];							inform_L[100][4] = l_cell_wire[104];							inform_L[116][4] = l_cell_wire[105];							inform_L[101][4] = l_cell_wire[106];							inform_L[117][4] = l_cell_wire[107];							inform_L[102][4] = l_cell_wire[108];							inform_L[118][4] = l_cell_wire[109];							inform_L[103][4] = l_cell_wire[110];							inform_L[119][4] = l_cell_wire[111];							inform_L[104][4] = l_cell_wire[112];							inform_L[120][4] = l_cell_wire[113];							inform_L[105][4] = l_cell_wire[114];							inform_L[121][4] = l_cell_wire[115];							inform_L[106][4] = l_cell_wire[116];							inform_L[122][4] = l_cell_wire[117];							inform_L[107][4] = l_cell_wire[118];							inform_L[123][4] = l_cell_wire[119];							inform_L[108][4] = l_cell_wire[120];							inform_L[124][4] = l_cell_wire[121];							inform_L[109][4] = l_cell_wire[122];							inform_L[125][4] = l_cell_wire[123];							inform_L[110][4] = l_cell_wire[124];							inform_L[126][4] = l_cell_wire[125];							inform_L[111][4] = l_cell_wire[126];							inform_L[127][4] = l_cell_wire[127];							inform_L[128][4] = l_cell_wire[128];							inform_L[144][4] = l_cell_wire[129];							inform_L[129][4] = l_cell_wire[130];							inform_L[145][4] = l_cell_wire[131];							inform_L[130][4] = l_cell_wire[132];							inform_L[146][4] = l_cell_wire[133];							inform_L[131][4] = l_cell_wire[134];							inform_L[147][4] = l_cell_wire[135];							inform_L[132][4] = l_cell_wire[136];							inform_L[148][4] = l_cell_wire[137];							inform_L[133][4] = l_cell_wire[138];							inform_L[149][4] = l_cell_wire[139];							inform_L[134][4] = l_cell_wire[140];							inform_L[150][4] = l_cell_wire[141];							inform_L[135][4] = l_cell_wire[142];							inform_L[151][4] = l_cell_wire[143];							inform_L[136][4] = l_cell_wire[144];							inform_L[152][4] = l_cell_wire[145];							inform_L[137][4] = l_cell_wire[146];							inform_L[153][4] = l_cell_wire[147];							inform_L[138][4] = l_cell_wire[148];							inform_L[154][4] = l_cell_wire[149];							inform_L[139][4] = l_cell_wire[150];							inform_L[155][4] = l_cell_wire[151];							inform_L[140][4] = l_cell_wire[152];							inform_L[156][4] = l_cell_wire[153];							inform_L[141][4] = l_cell_wire[154];							inform_L[157][4] = l_cell_wire[155];							inform_L[142][4] = l_cell_wire[156];							inform_L[158][4] = l_cell_wire[157];							inform_L[143][4] = l_cell_wire[158];							inform_L[159][4] = l_cell_wire[159];							inform_L[160][4] = l_cell_wire[160];							inform_L[176][4] = l_cell_wire[161];							inform_L[161][4] = l_cell_wire[162];							inform_L[177][4] = l_cell_wire[163];							inform_L[162][4] = l_cell_wire[164];							inform_L[178][4] = l_cell_wire[165];							inform_L[163][4] = l_cell_wire[166];							inform_L[179][4] = l_cell_wire[167];							inform_L[164][4] = l_cell_wire[168];							inform_L[180][4] = l_cell_wire[169];							inform_L[165][4] = l_cell_wire[170];							inform_L[181][4] = l_cell_wire[171];							inform_L[166][4] = l_cell_wire[172];							inform_L[182][4] = l_cell_wire[173];							inform_L[167][4] = l_cell_wire[174];							inform_L[183][4] = l_cell_wire[175];							inform_L[168][4] = l_cell_wire[176];							inform_L[184][4] = l_cell_wire[177];							inform_L[169][4] = l_cell_wire[178];							inform_L[185][4] = l_cell_wire[179];							inform_L[170][4] = l_cell_wire[180];							inform_L[186][4] = l_cell_wire[181];							inform_L[171][4] = l_cell_wire[182];							inform_L[187][4] = l_cell_wire[183];							inform_L[172][4] = l_cell_wire[184];							inform_L[188][4] = l_cell_wire[185];							inform_L[173][4] = l_cell_wire[186];							inform_L[189][4] = l_cell_wire[187];							inform_L[174][4] = l_cell_wire[188];							inform_L[190][4] = l_cell_wire[189];							inform_L[175][4] = l_cell_wire[190];							inform_L[191][4] = l_cell_wire[191];							inform_L[192][4] = l_cell_wire[192];							inform_L[208][4] = l_cell_wire[193];							inform_L[193][4] = l_cell_wire[194];							inform_L[209][4] = l_cell_wire[195];							inform_L[194][4] = l_cell_wire[196];							inform_L[210][4] = l_cell_wire[197];							inform_L[195][4] = l_cell_wire[198];							inform_L[211][4] = l_cell_wire[199];							inform_L[196][4] = l_cell_wire[200];							inform_L[212][4] = l_cell_wire[201];							inform_L[197][4] = l_cell_wire[202];							inform_L[213][4] = l_cell_wire[203];							inform_L[198][4] = l_cell_wire[204];							inform_L[214][4] = l_cell_wire[205];							inform_L[199][4] = l_cell_wire[206];							inform_L[215][4] = l_cell_wire[207];							inform_L[200][4] = l_cell_wire[208];							inform_L[216][4] = l_cell_wire[209];							inform_L[201][4] = l_cell_wire[210];							inform_L[217][4] = l_cell_wire[211];							inform_L[202][4] = l_cell_wire[212];							inform_L[218][4] = l_cell_wire[213];							inform_L[203][4] = l_cell_wire[214];							inform_L[219][4] = l_cell_wire[215];							inform_L[204][4] = l_cell_wire[216];							inform_L[220][4] = l_cell_wire[217];							inform_L[205][4] = l_cell_wire[218];							inform_L[221][4] = l_cell_wire[219];							inform_L[206][4] = l_cell_wire[220];							inform_L[222][4] = l_cell_wire[221];							inform_L[207][4] = l_cell_wire[222];							inform_L[223][4] = l_cell_wire[223];							inform_L[224][4] = l_cell_wire[224];							inform_L[240][4] = l_cell_wire[225];							inform_L[225][4] = l_cell_wire[226];							inform_L[241][4] = l_cell_wire[227];							inform_L[226][4] = l_cell_wire[228];							inform_L[242][4] = l_cell_wire[229];							inform_L[227][4] = l_cell_wire[230];							inform_L[243][4] = l_cell_wire[231];							inform_L[228][4] = l_cell_wire[232];							inform_L[244][4] = l_cell_wire[233];							inform_L[229][4] = l_cell_wire[234];							inform_L[245][4] = l_cell_wire[235];							inform_L[230][4] = l_cell_wire[236];							inform_L[246][4] = l_cell_wire[237];							inform_L[231][4] = l_cell_wire[238];							inform_L[247][4] = l_cell_wire[239];							inform_L[232][4] = l_cell_wire[240];							inform_L[248][4] = l_cell_wire[241];							inform_L[233][4] = l_cell_wire[242];							inform_L[249][4] = l_cell_wire[243];							inform_L[234][4] = l_cell_wire[244];							inform_L[250][4] = l_cell_wire[245];							inform_L[235][4] = l_cell_wire[246];							inform_L[251][4] = l_cell_wire[247];							inform_L[236][4] = l_cell_wire[248];							inform_L[252][4] = l_cell_wire[249];							inform_L[237][4] = l_cell_wire[250];							inform_L[253][4] = l_cell_wire[251];							inform_L[238][4] = l_cell_wire[252];							inform_L[254][4] = l_cell_wire[253];							inform_L[239][4] = l_cell_wire[254];							inform_L[255][4] = l_cell_wire[255];							inform_L[256][4] = l_cell_wire[256];							inform_L[272][4] = l_cell_wire[257];							inform_L[257][4] = l_cell_wire[258];							inform_L[273][4] = l_cell_wire[259];							inform_L[258][4] = l_cell_wire[260];							inform_L[274][4] = l_cell_wire[261];							inform_L[259][4] = l_cell_wire[262];							inform_L[275][4] = l_cell_wire[263];							inform_L[260][4] = l_cell_wire[264];							inform_L[276][4] = l_cell_wire[265];							inform_L[261][4] = l_cell_wire[266];							inform_L[277][4] = l_cell_wire[267];							inform_L[262][4] = l_cell_wire[268];							inform_L[278][4] = l_cell_wire[269];							inform_L[263][4] = l_cell_wire[270];							inform_L[279][4] = l_cell_wire[271];							inform_L[264][4] = l_cell_wire[272];							inform_L[280][4] = l_cell_wire[273];							inform_L[265][4] = l_cell_wire[274];							inform_L[281][4] = l_cell_wire[275];							inform_L[266][4] = l_cell_wire[276];							inform_L[282][4] = l_cell_wire[277];							inform_L[267][4] = l_cell_wire[278];							inform_L[283][4] = l_cell_wire[279];							inform_L[268][4] = l_cell_wire[280];							inform_L[284][4] = l_cell_wire[281];							inform_L[269][4] = l_cell_wire[282];							inform_L[285][4] = l_cell_wire[283];							inform_L[270][4] = l_cell_wire[284];							inform_L[286][4] = l_cell_wire[285];							inform_L[271][4] = l_cell_wire[286];							inform_L[287][4] = l_cell_wire[287];							inform_L[288][4] = l_cell_wire[288];							inform_L[304][4] = l_cell_wire[289];							inform_L[289][4] = l_cell_wire[290];							inform_L[305][4] = l_cell_wire[291];							inform_L[290][4] = l_cell_wire[292];							inform_L[306][4] = l_cell_wire[293];							inform_L[291][4] = l_cell_wire[294];							inform_L[307][4] = l_cell_wire[295];							inform_L[292][4] = l_cell_wire[296];							inform_L[308][4] = l_cell_wire[297];							inform_L[293][4] = l_cell_wire[298];							inform_L[309][4] = l_cell_wire[299];							inform_L[294][4] = l_cell_wire[300];							inform_L[310][4] = l_cell_wire[301];							inform_L[295][4] = l_cell_wire[302];							inform_L[311][4] = l_cell_wire[303];							inform_L[296][4] = l_cell_wire[304];							inform_L[312][4] = l_cell_wire[305];							inform_L[297][4] = l_cell_wire[306];							inform_L[313][4] = l_cell_wire[307];							inform_L[298][4] = l_cell_wire[308];							inform_L[314][4] = l_cell_wire[309];							inform_L[299][4] = l_cell_wire[310];							inform_L[315][4] = l_cell_wire[311];							inform_L[300][4] = l_cell_wire[312];							inform_L[316][4] = l_cell_wire[313];							inform_L[301][4] = l_cell_wire[314];							inform_L[317][4] = l_cell_wire[315];							inform_L[302][4] = l_cell_wire[316];							inform_L[318][4] = l_cell_wire[317];							inform_L[303][4] = l_cell_wire[318];							inform_L[319][4] = l_cell_wire[319];							inform_L[320][4] = l_cell_wire[320];							inform_L[336][4] = l_cell_wire[321];							inform_L[321][4] = l_cell_wire[322];							inform_L[337][4] = l_cell_wire[323];							inform_L[322][4] = l_cell_wire[324];							inform_L[338][4] = l_cell_wire[325];							inform_L[323][4] = l_cell_wire[326];							inform_L[339][4] = l_cell_wire[327];							inform_L[324][4] = l_cell_wire[328];							inform_L[340][4] = l_cell_wire[329];							inform_L[325][4] = l_cell_wire[330];							inform_L[341][4] = l_cell_wire[331];							inform_L[326][4] = l_cell_wire[332];							inform_L[342][4] = l_cell_wire[333];							inform_L[327][4] = l_cell_wire[334];							inform_L[343][4] = l_cell_wire[335];							inform_L[328][4] = l_cell_wire[336];							inform_L[344][4] = l_cell_wire[337];							inform_L[329][4] = l_cell_wire[338];							inform_L[345][4] = l_cell_wire[339];							inform_L[330][4] = l_cell_wire[340];							inform_L[346][4] = l_cell_wire[341];							inform_L[331][4] = l_cell_wire[342];							inform_L[347][4] = l_cell_wire[343];							inform_L[332][4] = l_cell_wire[344];							inform_L[348][4] = l_cell_wire[345];							inform_L[333][4] = l_cell_wire[346];							inform_L[349][4] = l_cell_wire[347];							inform_L[334][4] = l_cell_wire[348];							inform_L[350][4] = l_cell_wire[349];							inform_L[335][4] = l_cell_wire[350];							inform_L[351][4] = l_cell_wire[351];							inform_L[352][4] = l_cell_wire[352];							inform_L[368][4] = l_cell_wire[353];							inform_L[353][4] = l_cell_wire[354];							inform_L[369][4] = l_cell_wire[355];							inform_L[354][4] = l_cell_wire[356];							inform_L[370][4] = l_cell_wire[357];							inform_L[355][4] = l_cell_wire[358];							inform_L[371][4] = l_cell_wire[359];							inform_L[356][4] = l_cell_wire[360];							inform_L[372][4] = l_cell_wire[361];							inform_L[357][4] = l_cell_wire[362];							inform_L[373][4] = l_cell_wire[363];							inform_L[358][4] = l_cell_wire[364];							inform_L[374][4] = l_cell_wire[365];							inform_L[359][4] = l_cell_wire[366];							inform_L[375][4] = l_cell_wire[367];							inform_L[360][4] = l_cell_wire[368];							inform_L[376][4] = l_cell_wire[369];							inform_L[361][4] = l_cell_wire[370];							inform_L[377][4] = l_cell_wire[371];							inform_L[362][4] = l_cell_wire[372];							inform_L[378][4] = l_cell_wire[373];							inform_L[363][4] = l_cell_wire[374];							inform_L[379][4] = l_cell_wire[375];							inform_L[364][4] = l_cell_wire[376];							inform_L[380][4] = l_cell_wire[377];							inform_L[365][4] = l_cell_wire[378];							inform_L[381][4] = l_cell_wire[379];							inform_L[366][4] = l_cell_wire[380];							inform_L[382][4] = l_cell_wire[381];							inform_L[367][4] = l_cell_wire[382];							inform_L[383][4] = l_cell_wire[383];							inform_L[384][4] = l_cell_wire[384];							inform_L[400][4] = l_cell_wire[385];							inform_L[385][4] = l_cell_wire[386];							inform_L[401][4] = l_cell_wire[387];							inform_L[386][4] = l_cell_wire[388];							inform_L[402][4] = l_cell_wire[389];							inform_L[387][4] = l_cell_wire[390];							inform_L[403][4] = l_cell_wire[391];							inform_L[388][4] = l_cell_wire[392];							inform_L[404][4] = l_cell_wire[393];							inform_L[389][4] = l_cell_wire[394];							inform_L[405][4] = l_cell_wire[395];							inform_L[390][4] = l_cell_wire[396];							inform_L[406][4] = l_cell_wire[397];							inform_L[391][4] = l_cell_wire[398];							inform_L[407][4] = l_cell_wire[399];							inform_L[392][4] = l_cell_wire[400];							inform_L[408][4] = l_cell_wire[401];							inform_L[393][4] = l_cell_wire[402];							inform_L[409][4] = l_cell_wire[403];							inform_L[394][4] = l_cell_wire[404];							inform_L[410][4] = l_cell_wire[405];							inform_L[395][4] = l_cell_wire[406];							inform_L[411][4] = l_cell_wire[407];							inform_L[396][4] = l_cell_wire[408];							inform_L[412][4] = l_cell_wire[409];							inform_L[397][4] = l_cell_wire[410];							inform_L[413][4] = l_cell_wire[411];							inform_L[398][4] = l_cell_wire[412];							inform_L[414][4] = l_cell_wire[413];							inform_L[399][4] = l_cell_wire[414];							inform_L[415][4] = l_cell_wire[415];							inform_L[416][4] = l_cell_wire[416];							inform_L[432][4] = l_cell_wire[417];							inform_L[417][4] = l_cell_wire[418];							inform_L[433][4] = l_cell_wire[419];							inform_L[418][4] = l_cell_wire[420];							inform_L[434][4] = l_cell_wire[421];							inform_L[419][4] = l_cell_wire[422];							inform_L[435][4] = l_cell_wire[423];							inform_L[420][4] = l_cell_wire[424];							inform_L[436][4] = l_cell_wire[425];							inform_L[421][4] = l_cell_wire[426];							inform_L[437][4] = l_cell_wire[427];							inform_L[422][4] = l_cell_wire[428];							inform_L[438][4] = l_cell_wire[429];							inform_L[423][4] = l_cell_wire[430];							inform_L[439][4] = l_cell_wire[431];							inform_L[424][4] = l_cell_wire[432];							inform_L[440][4] = l_cell_wire[433];							inform_L[425][4] = l_cell_wire[434];							inform_L[441][4] = l_cell_wire[435];							inform_L[426][4] = l_cell_wire[436];							inform_L[442][4] = l_cell_wire[437];							inform_L[427][4] = l_cell_wire[438];							inform_L[443][4] = l_cell_wire[439];							inform_L[428][4] = l_cell_wire[440];							inform_L[444][4] = l_cell_wire[441];							inform_L[429][4] = l_cell_wire[442];							inform_L[445][4] = l_cell_wire[443];							inform_L[430][4] = l_cell_wire[444];							inform_L[446][4] = l_cell_wire[445];							inform_L[431][4] = l_cell_wire[446];							inform_L[447][4] = l_cell_wire[447];							inform_L[448][4] = l_cell_wire[448];							inform_L[464][4] = l_cell_wire[449];							inform_L[449][4] = l_cell_wire[450];							inform_L[465][4] = l_cell_wire[451];							inform_L[450][4] = l_cell_wire[452];							inform_L[466][4] = l_cell_wire[453];							inform_L[451][4] = l_cell_wire[454];							inform_L[467][4] = l_cell_wire[455];							inform_L[452][4] = l_cell_wire[456];							inform_L[468][4] = l_cell_wire[457];							inform_L[453][4] = l_cell_wire[458];							inform_L[469][4] = l_cell_wire[459];							inform_L[454][4] = l_cell_wire[460];							inform_L[470][4] = l_cell_wire[461];							inform_L[455][4] = l_cell_wire[462];							inform_L[471][4] = l_cell_wire[463];							inform_L[456][4] = l_cell_wire[464];							inform_L[472][4] = l_cell_wire[465];							inform_L[457][4] = l_cell_wire[466];							inform_L[473][4] = l_cell_wire[467];							inform_L[458][4] = l_cell_wire[468];							inform_L[474][4] = l_cell_wire[469];							inform_L[459][4] = l_cell_wire[470];							inform_L[475][4] = l_cell_wire[471];							inform_L[460][4] = l_cell_wire[472];							inform_L[476][4] = l_cell_wire[473];							inform_L[461][4] = l_cell_wire[474];							inform_L[477][4] = l_cell_wire[475];							inform_L[462][4] = l_cell_wire[476];							inform_L[478][4] = l_cell_wire[477];							inform_L[463][4] = l_cell_wire[478];							inform_L[479][4] = l_cell_wire[479];							inform_L[480][4] = l_cell_wire[480];							inform_L[496][4] = l_cell_wire[481];							inform_L[481][4] = l_cell_wire[482];							inform_L[497][4] = l_cell_wire[483];							inform_L[482][4] = l_cell_wire[484];							inform_L[498][4] = l_cell_wire[485];							inform_L[483][4] = l_cell_wire[486];							inform_L[499][4] = l_cell_wire[487];							inform_L[484][4] = l_cell_wire[488];							inform_L[500][4] = l_cell_wire[489];							inform_L[485][4] = l_cell_wire[490];							inform_L[501][4] = l_cell_wire[491];							inform_L[486][4] = l_cell_wire[492];							inform_L[502][4] = l_cell_wire[493];							inform_L[487][4] = l_cell_wire[494];							inform_L[503][4] = l_cell_wire[495];							inform_L[488][4] = l_cell_wire[496];							inform_L[504][4] = l_cell_wire[497];							inform_L[489][4] = l_cell_wire[498];							inform_L[505][4] = l_cell_wire[499];							inform_L[490][4] = l_cell_wire[500];							inform_L[506][4] = l_cell_wire[501];							inform_L[491][4] = l_cell_wire[502];							inform_L[507][4] = l_cell_wire[503];							inform_L[492][4] = l_cell_wire[504];							inform_L[508][4] = l_cell_wire[505];							inform_L[493][4] = l_cell_wire[506];							inform_L[509][4] = l_cell_wire[507];							inform_L[494][4] = l_cell_wire[508];							inform_L[510][4] = l_cell_wire[509];							inform_L[495][4] = l_cell_wire[510];							inform_L[511][4] = l_cell_wire[511];							inform_L[512][4] = l_cell_wire[512];							inform_L[528][4] = l_cell_wire[513];							inform_L[513][4] = l_cell_wire[514];							inform_L[529][4] = l_cell_wire[515];							inform_L[514][4] = l_cell_wire[516];							inform_L[530][4] = l_cell_wire[517];							inform_L[515][4] = l_cell_wire[518];							inform_L[531][4] = l_cell_wire[519];							inform_L[516][4] = l_cell_wire[520];							inform_L[532][4] = l_cell_wire[521];							inform_L[517][4] = l_cell_wire[522];							inform_L[533][4] = l_cell_wire[523];							inform_L[518][4] = l_cell_wire[524];							inform_L[534][4] = l_cell_wire[525];							inform_L[519][4] = l_cell_wire[526];							inform_L[535][4] = l_cell_wire[527];							inform_L[520][4] = l_cell_wire[528];							inform_L[536][4] = l_cell_wire[529];							inform_L[521][4] = l_cell_wire[530];							inform_L[537][4] = l_cell_wire[531];							inform_L[522][4] = l_cell_wire[532];							inform_L[538][4] = l_cell_wire[533];							inform_L[523][4] = l_cell_wire[534];							inform_L[539][4] = l_cell_wire[535];							inform_L[524][4] = l_cell_wire[536];							inform_L[540][4] = l_cell_wire[537];							inform_L[525][4] = l_cell_wire[538];							inform_L[541][4] = l_cell_wire[539];							inform_L[526][4] = l_cell_wire[540];							inform_L[542][4] = l_cell_wire[541];							inform_L[527][4] = l_cell_wire[542];							inform_L[543][4] = l_cell_wire[543];							inform_L[544][4] = l_cell_wire[544];							inform_L[560][4] = l_cell_wire[545];							inform_L[545][4] = l_cell_wire[546];							inform_L[561][4] = l_cell_wire[547];							inform_L[546][4] = l_cell_wire[548];							inform_L[562][4] = l_cell_wire[549];							inform_L[547][4] = l_cell_wire[550];							inform_L[563][4] = l_cell_wire[551];							inform_L[548][4] = l_cell_wire[552];							inform_L[564][4] = l_cell_wire[553];							inform_L[549][4] = l_cell_wire[554];							inform_L[565][4] = l_cell_wire[555];							inform_L[550][4] = l_cell_wire[556];							inform_L[566][4] = l_cell_wire[557];							inform_L[551][4] = l_cell_wire[558];							inform_L[567][4] = l_cell_wire[559];							inform_L[552][4] = l_cell_wire[560];							inform_L[568][4] = l_cell_wire[561];							inform_L[553][4] = l_cell_wire[562];							inform_L[569][4] = l_cell_wire[563];							inform_L[554][4] = l_cell_wire[564];							inform_L[570][4] = l_cell_wire[565];							inform_L[555][4] = l_cell_wire[566];							inform_L[571][4] = l_cell_wire[567];							inform_L[556][4] = l_cell_wire[568];							inform_L[572][4] = l_cell_wire[569];							inform_L[557][4] = l_cell_wire[570];							inform_L[573][4] = l_cell_wire[571];							inform_L[558][4] = l_cell_wire[572];							inform_L[574][4] = l_cell_wire[573];							inform_L[559][4] = l_cell_wire[574];							inform_L[575][4] = l_cell_wire[575];							inform_L[576][4] = l_cell_wire[576];							inform_L[592][4] = l_cell_wire[577];							inform_L[577][4] = l_cell_wire[578];							inform_L[593][4] = l_cell_wire[579];							inform_L[578][4] = l_cell_wire[580];							inform_L[594][4] = l_cell_wire[581];							inform_L[579][4] = l_cell_wire[582];							inform_L[595][4] = l_cell_wire[583];							inform_L[580][4] = l_cell_wire[584];							inform_L[596][4] = l_cell_wire[585];							inform_L[581][4] = l_cell_wire[586];							inform_L[597][4] = l_cell_wire[587];							inform_L[582][4] = l_cell_wire[588];							inform_L[598][4] = l_cell_wire[589];							inform_L[583][4] = l_cell_wire[590];							inform_L[599][4] = l_cell_wire[591];							inform_L[584][4] = l_cell_wire[592];							inform_L[600][4] = l_cell_wire[593];							inform_L[585][4] = l_cell_wire[594];							inform_L[601][4] = l_cell_wire[595];							inform_L[586][4] = l_cell_wire[596];							inform_L[602][4] = l_cell_wire[597];							inform_L[587][4] = l_cell_wire[598];							inform_L[603][4] = l_cell_wire[599];							inform_L[588][4] = l_cell_wire[600];							inform_L[604][4] = l_cell_wire[601];							inform_L[589][4] = l_cell_wire[602];							inform_L[605][4] = l_cell_wire[603];							inform_L[590][4] = l_cell_wire[604];							inform_L[606][4] = l_cell_wire[605];							inform_L[591][4] = l_cell_wire[606];							inform_L[607][4] = l_cell_wire[607];							inform_L[608][4] = l_cell_wire[608];							inform_L[624][4] = l_cell_wire[609];							inform_L[609][4] = l_cell_wire[610];							inform_L[625][4] = l_cell_wire[611];							inform_L[610][4] = l_cell_wire[612];							inform_L[626][4] = l_cell_wire[613];							inform_L[611][4] = l_cell_wire[614];							inform_L[627][4] = l_cell_wire[615];							inform_L[612][4] = l_cell_wire[616];							inform_L[628][4] = l_cell_wire[617];							inform_L[613][4] = l_cell_wire[618];							inform_L[629][4] = l_cell_wire[619];							inform_L[614][4] = l_cell_wire[620];							inform_L[630][4] = l_cell_wire[621];							inform_L[615][4] = l_cell_wire[622];							inform_L[631][4] = l_cell_wire[623];							inform_L[616][4] = l_cell_wire[624];							inform_L[632][4] = l_cell_wire[625];							inform_L[617][4] = l_cell_wire[626];							inform_L[633][4] = l_cell_wire[627];							inform_L[618][4] = l_cell_wire[628];							inform_L[634][4] = l_cell_wire[629];							inform_L[619][4] = l_cell_wire[630];							inform_L[635][4] = l_cell_wire[631];							inform_L[620][4] = l_cell_wire[632];							inform_L[636][4] = l_cell_wire[633];							inform_L[621][4] = l_cell_wire[634];							inform_L[637][4] = l_cell_wire[635];							inform_L[622][4] = l_cell_wire[636];							inform_L[638][4] = l_cell_wire[637];							inform_L[623][4] = l_cell_wire[638];							inform_L[639][4] = l_cell_wire[639];							inform_L[640][4] = l_cell_wire[640];							inform_L[656][4] = l_cell_wire[641];							inform_L[641][4] = l_cell_wire[642];							inform_L[657][4] = l_cell_wire[643];							inform_L[642][4] = l_cell_wire[644];							inform_L[658][4] = l_cell_wire[645];							inform_L[643][4] = l_cell_wire[646];							inform_L[659][4] = l_cell_wire[647];							inform_L[644][4] = l_cell_wire[648];							inform_L[660][4] = l_cell_wire[649];							inform_L[645][4] = l_cell_wire[650];							inform_L[661][4] = l_cell_wire[651];							inform_L[646][4] = l_cell_wire[652];							inform_L[662][4] = l_cell_wire[653];							inform_L[647][4] = l_cell_wire[654];							inform_L[663][4] = l_cell_wire[655];							inform_L[648][4] = l_cell_wire[656];							inform_L[664][4] = l_cell_wire[657];							inform_L[649][4] = l_cell_wire[658];							inform_L[665][4] = l_cell_wire[659];							inform_L[650][4] = l_cell_wire[660];							inform_L[666][4] = l_cell_wire[661];							inform_L[651][4] = l_cell_wire[662];							inform_L[667][4] = l_cell_wire[663];							inform_L[652][4] = l_cell_wire[664];							inform_L[668][4] = l_cell_wire[665];							inform_L[653][4] = l_cell_wire[666];							inform_L[669][4] = l_cell_wire[667];							inform_L[654][4] = l_cell_wire[668];							inform_L[670][4] = l_cell_wire[669];							inform_L[655][4] = l_cell_wire[670];							inform_L[671][4] = l_cell_wire[671];							inform_L[672][4] = l_cell_wire[672];							inform_L[688][4] = l_cell_wire[673];							inform_L[673][4] = l_cell_wire[674];							inform_L[689][4] = l_cell_wire[675];							inform_L[674][4] = l_cell_wire[676];							inform_L[690][4] = l_cell_wire[677];							inform_L[675][4] = l_cell_wire[678];							inform_L[691][4] = l_cell_wire[679];							inform_L[676][4] = l_cell_wire[680];							inform_L[692][4] = l_cell_wire[681];							inform_L[677][4] = l_cell_wire[682];							inform_L[693][4] = l_cell_wire[683];							inform_L[678][4] = l_cell_wire[684];							inform_L[694][4] = l_cell_wire[685];							inform_L[679][4] = l_cell_wire[686];							inform_L[695][4] = l_cell_wire[687];							inform_L[680][4] = l_cell_wire[688];							inform_L[696][4] = l_cell_wire[689];							inform_L[681][4] = l_cell_wire[690];							inform_L[697][4] = l_cell_wire[691];							inform_L[682][4] = l_cell_wire[692];							inform_L[698][4] = l_cell_wire[693];							inform_L[683][4] = l_cell_wire[694];							inform_L[699][4] = l_cell_wire[695];							inform_L[684][4] = l_cell_wire[696];							inform_L[700][4] = l_cell_wire[697];							inform_L[685][4] = l_cell_wire[698];							inform_L[701][4] = l_cell_wire[699];							inform_L[686][4] = l_cell_wire[700];							inform_L[702][4] = l_cell_wire[701];							inform_L[687][4] = l_cell_wire[702];							inform_L[703][4] = l_cell_wire[703];							inform_L[704][4] = l_cell_wire[704];							inform_L[720][4] = l_cell_wire[705];							inform_L[705][4] = l_cell_wire[706];							inform_L[721][4] = l_cell_wire[707];							inform_L[706][4] = l_cell_wire[708];							inform_L[722][4] = l_cell_wire[709];							inform_L[707][4] = l_cell_wire[710];							inform_L[723][4] = l_cell_wire[711];							inform_L[708][4] = l_cell_wire[712];							inform_L[724][4] = l_cell_wire[713];							inform_L[709][4] = l_cell_wire[714];							inform_L[725][4] = l_cell_wire[715];							inform_L[710][4] = l_cell_wire[716];							inform_L[726][4] = l_cell_wire[717];							inform_L[711][4] = l_cell_wire[718];							inform_L[727][4] = l_cell_wire[719];							inform_L[712][4] = l_cell_wire[720];							inform_L[728][4] = l_cell_wire[721];							inform_L[713][4] = l_cell_wire[722];							inform_L[729][4] = l_cell_wire[723];							inform_L[714][4] = l_cell_wire[724];							inform_L[730][4] = l_cell_wire[725];							inform_L[715][4] = l_cell_wire[726];							inform_L[731][4] = l_cell_wire[727];							inform_L[716][4] = l_cell_wire[728];							inform_L[732][4] = l_cell_wire[729];							inform_L[717][4] = l_cell_wire[730];							inform_L[733][4] = l_cell_wire[731];							inform_L[718][4] = l_cell_wire[732];							inform_L[734][4] = l_cell_wire[733];							inform_L[719][4] = l_cell_wire[734];							inform_L[735][4] = l_cell_wire[735];							inform_L[736][4] = l_cell_wire[736];							inform_L[752][4] = l_cell_wire[737];							inform_L[737][4] = l_cell_wire[738];							inform_L[753][4] = l_cell_wire[739];							inform_L[738][4] = l_cell_wire[740];							inform_L[754][4] = l_cell_wire[741];							inform_L[739][4] = l_cell_wire[742];							inform_L[755][4] = l_cell_wire[743];							inform_L[740][4] = l_cell_wire[744];							inform_L[756][4] = l_cell_wire[745];							inform_L[741][4] = l_cell_wire[746];							inform_L[757][4] = l_cell_wire[747];							inform_L[742][4] = l_cell_wire[748];							inform_L[758][4] = l_cell_wire[749];							inform_L[743][4] = l_cell_wire[750];							inform_L[759][4] = l_cell_wire[751];							inform_L[744][4] = l_cell_wire[752];							inform_L[760][4] = l_cell_wire[753];							inform_L[745][4] = l_cell_wire[754];							inform_L[761][4] = l_cell_wire[755];							inform_L[746][4] = l_cell_wire[756];							inform_L[762][4] = l_cell_wire[757];							inform_L[747][4] = l_cell_wire[758];							inform_L[763][4] = l_cell_wire[759];							inform_L[748][4] = l_cell_wire[760];							inform_L[764][4] = l_cell_wire[761];							inform_L[749][4] = l_cell_wire[762];							inform_L[765][4] = l_cell_wire[763];							inform_L[750][4] = l_cell_wire[764];							inform_L[766][4] = l_cell_wire[765];							inform_L[751][4] = l_cell_wire[766];							inform_L[767][4] = l_cell_wire[767];							inform_L[768][4] = l_cell_wire[768];							inform_L[784][4] = l_cell_wire[769];							inform_L[769][4] = l_cell_wire[770];							inform_L[785][4] = l_cell_wire[771];							inform_L[770][4] = l_cell_wire[772];							inform_L[786][4] = l_cell_wire[773];							inform_L[771][4] = l_cell_wire[774];							inform_L[787][4] = l_cell_wire[775];							inform_L[772][4] = l_cell_wire[776];							inform_L[788][4] = l_cell_wire[777];							inform_L[773][4] = l_cell_wire[778];							inform_L[789][4] = l_cell_wire[779];							inform_L[774][4] = l_cell_wire[780];							inform_L[790][4] = l_cell_wire[781];							inform_L[775][4] = l_cell_wire[782];							inform_L[791][4] = l_cell_wire[783];							inform_L[776][4] = l_cell_wire[784];							inform_L[792][4] = l_cell_wire[785];							inform_L[777][4] = l_cell_wire[786];							inform_L[793][4] = l_cell_wire[787];							inform_L[778][4] = l_cell_wire[788];							inform_L[794][4] = l_cell_wire[789];							inform_L[779][4] = l_cell_wire[790];							inform_L[795][4] = l_cell_wire[791];							inform_L[780][4] = l_cell_wire[792];							inform_L[796][4] = l_cell_wire[793];							inform_L[781][4] = l_cell_wire[794];							inform_L[797][4] = l_cell_wire[795];							inform_L[782][4] = l_cell_wire[796];							inform_L[798][4] = l_cell_wire[797];							inform_L[783][4] = l_cell_wire[798];							inform_L[799][4] = l_cell_wire[799];							inform_L[800][4] = l_cell_wire[800];							inform_L[816][4] = l_cell_wire[801];							inform_L[801][4] = l_cell_wire[802];							inform_L[817][4] = l_cell_wire[803];							inform_L[802][4] = l_cell_wire[804];							inform_L[818][4] = l_cell_wire[805];							inform_L[803][4] = l_cell_wire[806];							inform_L[819][4] = l_cell_wire[807];							inform_L[804][4] = l_cell_wire[808];							inform_L[820][4] = l_cell_wire[809];							inform_L[805][4] = l_cell_wire[810];							inform_L[821][4] = l_cell_wire[811];							inform_L[806][4] = l_cell_wire[812];							inform_L[822][4] = l_cell_wire[813];							inform_L[807][4] = l_cell_wire[814];							inform_L[823][4] = l_cell_wire[815];							inform_L[808][4] = l_cell_wire[816];							inform_L[824][4] = l_cell_wire[817];							inform_L[809][4] = l_cell_wire[818];							inform_L[825][4] = l_cell_wire[819];							inform_L[810][4] = l_cell_wire[820];							inform_L[826][4] = l_cell_wire[821];							inform_L[811][4] = l_cell_wire[822];							inform_L[827][4] = l_cell_wire[823];							inform_L[812][4] = l_cell_wire[824];							inform_L[828][4] = l_cell_wire[825];							inform_L[813][4] = l_cell_wire[826];							inform_L[829][4] = l_cell_wire[827];							inform_L[814][4] = l_cell_wire[828];							inform_L[830][4] = l_cell_wire[829];							inform_L[815][4] = l_cell_wire[830];							inform_L[831][4] = l_cell_wire[831];							inform_L[832][4] = l_cell_wire[832];							inform_L[848][4] = l_cell_wire[833];							inform_L[833][4] = l_cell_wire[834];							inform_L[849][4] = l_cell_wire[835];							inform_L[834][4] = l_cell_wire[836];							inform_L[850][4] = l_cell_wire[837];							inform_L[835][4] = l_cell_wire[838];							inform_L[851][4] = l_cell_wire[839];							inform_L[836][4] = l_cell_wire[840];							inform_L[852][4] = l_cell_wire[841];							inform_L[837][4] = l_cell_wire[842];							inform_L[853][4] = l_cell_wire[843];							inform_L[838][4] = l_cell_wire[844];							inform_L[854][4] = l_cell_wire[845];							inform_L[839][4] = l_cell_wire[846];							inform_L[855][4] = l_cell_wire[847];							inform_L[840][4] = l_cell_wire[848];							inform_L[856][4] = l_cell_wire[849];							inform_L[841][4] = l_cell_wire[850];							inform_L[857][4] = l_cell_wire[851];							inform_L[842][4] = l_cell_wire[852];							inform_L[858][4] = l_cell_wire[853];							inform_L[843][4] = l_cell_wire[854];							inform_L[859][4] = l_cell_wire[855];							inform_L[844][4] = l_cell_wire[856];							inform_L[860][4] = l_cell_wire[857];							inform_L[845][4] = l_cell_wire[858];							inform_L[861][4] = l_cell_wire[859];							inform_L[846][4] = l_cell_wire[860];							inform_L[862][4] = l_cell_wire[861];							inform_L[847][4] = l_cell_wire[862];							inform_L[863][4] = l_cell_wire[863];							inform_L[864][4] = l_cell_wire[864];							inform_L[880][4] = l_cell_wire[865];							inform_L[865][4] = l_cell_wire[866];							inform_L[881][4] = l_cell_wire[867];							inform_L[866][4] = l_cell_wire[868];							inform_L[882][4] = l_cell_wire[869];							inform_L[867][4] = l_cell_wire[870];							inform_L[883][4] = l_cell_wire[871];							inform_L[868][4] = l_cell_wire[872];							inform_L[884][4] = l_cell_wire[873];							inform_L[869][4] = l_cell_wire[874];							inform_L[885][4] = l_cell_wire[875];							inform_L[870][4] = l_cell_wire[876];							inform_L[886][4] = l_cell_wire[877];							inform_L[871][4] = l_cell_wire[878];							inform_L[887][4] = l_cell_wire[879];							inform_L[872][4] = l_cell_wire[880];							inform_L[888][4] = l_cell_wire[881];							inform_L[873][4] = l_cell_wire[882];							inform_L[889][4] = l_cell_wire[883];							inform_L[874][4] = l_cell_wire[884];							inform_L[890][4] = l_cell_wire[885];							inform_L[875][4] = l_cell_wire[886];							inform_L[891][4] = l_cell_wire[887];							inform_L[876][4] = l_cell_wire[888];							inform_L[892][4] = l_cell_wire[889];							inform_L[877][4] = l_cell_wire[890];							inform_L[893][4] = l_cell_wire[891];							inform_L[878][4] = l_cell_wire[892];							inform_L[894][4] = l_cell_wire[893];							inform_L[879][4] = l_cell_wire[894];							inform_L[895][4] = l_cell_wire[895];							inform_L[896][4] = l_cell_wire[896];							inform_L[912][4] = l_cell_wire[897];							inform_L[897][4] = l_cell_wire[898];							inform_L[913][4] = l_cell_wire[899];							inform_L[898][4] = l_cell_wire[900];							inform_L[914][4] = l_cell_wire[901];							inform_L[899][4] = l_cell_wire[902];							inform_L[915][4] = l_cell_wire[903];							inform_L[900][4] = l_cell_wire[904];							inform_L[916][4] = l_cell_wire[905];							inform_L[901][4] = l_cell_wire[906];							inform_L[917][4] = l_cell_wire[907];							inform_L[902][4] = l_cell_wire[908];							inform_L[918][4] = l_cell_wire[909];							inform_L[903][4] = l_cell_wire[910];							inform_L[919][4] = l_cell_wire[911];							inform_L[904][4] = l_cell_wire[912];							inform_L[920][4] = l_cell_wire[913];							inform_L[905][4] = l_cell_wire[914];							inform_L[921][4] = l_cell_wire[915];							inform_L[906][4] = l_cell_wire[916];							inform_L[922][4] = l_cell_wire[917];							inform_L[907][4] = l_cell_wire[918];							inform_L[923][4] = l_cell_wire[919];							inform_L[908][4] = l_cell_wire[920];							inform_L[924][4] = l_cell_wire[921];							inform_L[909][4] = l_cell_wire[922];							inform_L[925][4] = l_cell_wire[923];							inform_L[910][4] = l_cell_wire[924];							inform_L[926][4] = l_cell_wire[925];							inform_L[911][4] = l_cell_wire[926];							inform_L[927][4] = l_cell_wire[927];							inform_L[928][4] = l_cell_wire[928];							inform_L[944][4] = l_cell_wire[929];							inform_L[929][4] = l_cell_wire[930];							inform_L[945][4] = l_cell_wire[931];							inform_L[930][4] = l_cell_wire[932];							inform_L[946][4] = l_cell_wire[933];							inform_L[931][4] = l_cell_wire[934];							inform_L[947][4] = l_cell_wire[935];							inform_L[932][4] = l_cell_wire[936];							inform_L[948][4] = l_cell_wire[937];							inform_L[933][4] = l_cell_wire[938];							inform_L[949][4] = l_cell_wire[939];							inform_L[934][4] = l_cell_wire[940];							inform_L[950][4] = l_cell_wire[941];							inform_L[935][4] = l_cell_wire[942];							inform_L[951][4] = l_cell_wire[943];							inform_L[936][4] = l_cell_wire[944];							inform_L[952][4] = l_cell_wire[945];							inform_L[937][4] = l_cell_wire[946];							inform_L[953][4] = l_cell_wire[947];							inform_L[938][4] = l_cell_wire[948];							inform_L[954][4] = l_cell_wire[949];							inform_L[939][4] = l_cell_wire[950];							inform_L[955][4] = l_cell_wire[951];							inform_L[940][4] = l_cell_wire[952];							inform_L[956][4] = l_cell_wire[953];							inform_L[941][4] = l_cell_wire[954];							inform_L[957][4] = l_cell_wire[955];							inform_L[942][4] = l_cell_wire[956];							inform_L[958][4] = l_cell_wire[957];							inform_L[943][4] = l_cell_wire[958];							inform_L[959][4] = l_cell_wire[959];							inform_L[960][4] = l_cell_wire[960];							inform_L[976][4] = l_cell_wire[961];							inform_L[961][4] = l_cell_wire[962];							inform_L[977][4] = l_cell_wire[963];							inform_L[962][4] = l_cell_wire[964];							inform_L[978][4] = l_cell_wire[965];							inform_L[963][4] = l_cell_wire[966];							inform_L[979][4] = l_cell_wire[967];							inform_L[964][4] = l_cell_wire[968];							inform_L[980][4] = l_cell_wire[969];							inform_L[965][4] = l_cell_wire[970];							inform_L[981][4] = l_cell_wire[971];							inform_L[966][4] = l_cell_wire[972];							inform_L[982][4] = l_cell_wire[973];							inform_L[967][4] = l_cell_wire[974];							inform_L[983][4] = l_cell_wire[975];							inform_L[968][4] = l_cell_wire[976];							inform_L[984][4] = l_cell_wire[977];							inform_L[969][4] = l_cell_wire[978];							inform_L[985][4] = l_cell_wire[979];							inform_L[970][4] = l_cell_wire[980];							inform_L[986][4] = l_cell_wire[981];							inform_L[971][4] = l_cell_wire[982];							inform_L[987][4] = l_cell_wire[983];							inform_L[972][4] = l_cell_wire[984];							inform_L[988][4] = l_cell_wire[985];							inform_L[973][4] = l_cell_wire[986];							inform_L[989][4] = l_cell_wire[987];							inform_L[974][4] = l_cell_wire[988];							inform_L[990][4] = l_cell_wire[989];							inform_L[975][4] = l_cell_wire[990];							inform_L[991][4] = l_cell_wire[991];							inform_L[992][4] = l_cell_wire[992];							inform_L[1008][4] = l_cell_wire[993];							inform_L[993][4] = l_cell_wire[994];							inform_L[1009][4] = l_cell_wire[995];							inform_L[994][4] = l_cell_wire[996];							inform_L[1010][4] = l_cell_wire[997];							inform_L[995][4] = l_cell_wire[998];							inform_L[1011][4] = l_cell_wire[999];							inform_L[996][4] = l_cell_wire[1000];							inform_L[1012][4] = l_cell_wire[1001];							inform_L[997][4] = l_cell_wire[1002];							inform_L[1013][4] = l_cell_wire[1003];							inform_L[998][4] = l_cell_wire[1004];							inform_L[1014][4] = l_cell_wire[1005];							inform_L[999][4] = l_cell_wire[1006];							inform_L[1015][4] = l_cell_wire[1007];							inform_L[1000][4] = l_cell_wire[1008];							inform_L[1016][4] = l_cell_wire[1009];							inform_L[1001][4] = l_cell_wire[1010];							inform_L[1017][4] = l_cell_wire[1011];							inform_L[1002][4] = l_cell_wire[1012];							inform_L[1018][4] = l_cell_wire[1013];							inform_L[1003][4] = l_cell_wire[1014];							inform_L[1019][4] = l_cell_wire[1015];							inform_L[1004][4] = l_cell_wire[1016];							inform_L[1020][4] = l_cell_wire[1017];							inform_L[1005][4] = l_cell_wire[1018];							inform_L[1021][4] = l_cell_wire[1019];							inform_L[1006][4] = l_cell_wire[1020];							inform_L[1022][4] = l_cell_wire[1021];							inform_L[1007][4] = l_cell_wire[1022];							inform_L[1023][4] = l_cell_wire[1023];						end
						6:						begin							inform_R[0][6] = r_cell_wire[0];							inform_R[32][6] = r_cell_wire[1];							inform_R[1][6] = r_cell_wire[2];							inform_R[33][6] = r_cell_wire[3];							inform_R[2][6] = r_cell_wire[4];							inform_R[34][6] = r_cell_wire[5];							inform_R[3][6] = r_cell_wire[6];							inform_R[35][6] = r_cell_wire[7];							inform_R[4][6] = r_cell_wire[8];							inform_R[36][6] = r_cell_wire[9];							inform_R[5][6] = r_cell_wire[10];							inform_R[37][6] = r_cell_wire[11];							inform_R[6][6] = r_cell_wire[12];							inform_R[38][6] = r_cell_wire[13];							inform_R[7][6] = r_cell_wire[14];							inform_R[39][6] = r_cell_wire[15];							inform_R[8][6] = r_cell_wire[16];							inform_R[40][6] = r_cell_wire[17];							inform_R[9][6] = r_cell_wire[18];							inform_R[41][6] = r_cell_wire[19];							inform_R[10][6] = r_cell_wire[20];							inform_R[42][6] = r_cell_wire[21];							inform_R[11][6] = r_cell_wire[22];							inform_R[43][6] = r_cell_wire[23];							inform_R[12][6] = r_cell_wire[24];							inform_R[44][6] = r_cell_wire[25];							inform_R[13][6] = r_cell_wire[26];							inform_R[45][6] = r_cell_wire[27];							inform_R[14][6] = r_cell_wire[28];							inform_R[46][6] = r_cell_wire[29];							inform_R[15][6] = r_cell_wire[30];							inform_R[47][6] = r_cell_wire[31];							inform_R[16][6] = r_cell_wire[32];							inform_R[48][6] = r_cell_wire[33];							inform_R[17][6] = r_cell_wire[34];							inform_R[49][6] = r_cell_wire[35];							inform_R[18][6] = r_cell_wire[36];							inform_R[50][6] = r_cell_wire[37];							inform_R[19][6] = r_cell_wire[38];							inform_R[51][6] = r_cell_wire[39];							inform_R[20][6] = r_cell_wire[40];							inform_R[52][6] = r_cell_wire[41];							inform_R[21][6] = r_cell_wire[42];							inform_R[53][6] = r_cell_wire[43];							inform_R[22][6] = r_cell_wire[44];							inform_R[54][6] = r_cell_wire[45];							inform_R[23][6] = r_cell_wire[46];							inform_R[55][6] = r_cell_wire[47];							inform_R[24][6] = r_cell_wire[48];							inform_R[56][6] = r_cell_wire[49];							inform_R[25][6] = r_cell_wire[50];							inform_R[57][6] = r_cell_wire[51];							inform_R[26][6] = r_cell_wire[52];							inform_R[58][6] = r_cell_wire[53];							inform_R[27][6] = r_cell_wire[54];							inform_R[59][6] = r_cell_wire[55];							inform_R[28][6] = r_cell_wire[56];							inform_R[60][6] = r_cell_wire[57];							inform_R[29][6] = r_cell_wire[58];							inform_R[61][6] = r_cell_wire[59];							inform_R[30][6] = r_cell_wire[60];							inform_R[62][6] = r_cell_wire[61];							inform_R[31][6] = r_cell_wire[62];							inform_R[63][6] = r_cell_wire[63];							inform_R[64][6] = r_cell_wire[64];							inform_R[96][6] = r_cell_wire[65];							inform_R[65][6] = r_cell_wire[66];							inform_R[97][6] = r_cell_wire[67];							inform_R[66][6] = r_cell_wire[68];							inform_R[98][6] = r_cell_wire[69];							inform_R[67][6] = r_cell_wire[70];							inform_R[99][6] = r_cell_wire[71];							inform_R[68][6] = r_cell_wire[72];							inform_R[100][6] = r_cell_wire[73];							inform_R[69][6] = r_cell_wire[74];							inform_R[101][6] = r_cell_wire[75];							inform_R[70][6] = r_cell_wire[76];							inform_R[102][6] = r_cell_wire[77];							inform_R[71][6] = r_cell_wire[78];							inform_R[103][6] = r_cell_wire[79];							inform_R[72][6] = r_cell_wire[80];							inform_R[104][6] = r_cell_wire[81];							inform_R[73][6] = r_cell_wire[82];							inform_R[105][6] = r_cell_wire[83];							inform_R[74][6] = r_cell_wire[84];							inform_R[106][6] = r_cell_wire[85];							inform_R[75][6] = r_cell_wire[86];							inform_R[107][6] = r_cell_wire[87];							inform_R[76][6] = r_cell_wire[88];							inform_R[108][6] = r_cell_wire[89];							inform_R[77][6] = r_cell_wire[90];							inform_R[109][6] = r_cell_wire[91];							inform_R[78][6] = r_cell_wire[92];							inform_R[110][6] = r_cell_wire[93];							inform_R[79][6] = r_cell_wire[94];							inform_R[111][6] = r_cell_wire[95];							inform_R[80][6] = r_cell_wire[96];							inform_R[112][6] = r_cell_wire[97];							inform_R[81][6] = r_cell_wire[98];							inform_R[113][6] = r_cell_wire[99];							inform_R[82][6] = r_cell_wire[100];							inform_R[114][6] = r_cell_wire[101];							inform_R[83][6] = r_cell_wire[102];							inform_R[115][6] = r_cell_wire[103];							inform_R[84][6] = r_cell_wire[104];							inform_R[116][6] = r_cell_wire[105];							inform_R[85][6] = r_cell_wire[106];							inform_R[117][6] = r_cell_wire[107];							inform_R[86][6] = r_cell_wire[108];							inform_R[118][6] = r_cell_wire[109];							inform_R[87][6] = r_cell_wire[110];							inform_R[119][6] = r_cell_wire[111];							inform_R[88][6] = r_cell_wire[112];							inform_R[120][6] = r_cell_wire[113];							inform_R[89][6] = r_cell_wire[114];							inform_R[121][6] = r_cell_wire[115];							inform_R[90][6] = r_cell_wire[116];							inform_R[122][6] = r_cell_wire[117];							inform_R[91][6] = r_cell_wire[118];							inform_R[123][6] = r_cell_wire[119];							inform_R[92][6] = r_cell_wire[120];							inform_R[124][6] = r_cell_wire[121];							inform_R[93][6] = r_cell_wire[122];							inform_R[125][6] = r_cell_wire[123];							inform_R[94][6] = r_cell_wire[124];							inform_R[126][6] = r_cell_wire[125];							inform_R[95][6] = r_cell_wire[126];							inform_R[127][6] = r_cell_wire[127];							inform_R[128][6] = r_cell_wire[128];							inform_R[160][6] = r_cell_wire[129];							inform_R[129][6] = r_cell_wire[130];							inform_R[161][6] = r_cell_wire[131];							inform_R[130][6] = r_cell_wire[132];							inform_R[162][6] = r_cell_wire[133];							inform_R[131][6] = r_cell_wire[134];							inform_R[163][6] = r_cell_wire[135];							inform_R[132][6] = r_cell_wire[136];							inform_R[164][6] = r_cell_wire[137];							inform_R[133][6] = r_cell_wire[138];							inform_R[165][6] = r_cell_wire[139];							inform_R[134][6] = r_cell_wire[140];							inform_R[166][6] = r_cell_wire[141];							inform_R[135][6] = r_cell_wire[142];							inform_R[167][6] = r_cell_wire[143];							inform_R[136][6] = r_cell_wire[144];							inform_R[168][6] = r_cell_wire[145];							inform_R[137][6] = r_cell_wire[146];							inform_R[169][6] = r_cell_wire[147];							inform_R[138][6] = r_cell_wire[148];							inform_R[170][6] = r_cell_wire[149];							inform_R[139][6] = r_cell_wire[150];							inform_R[171][6] = r_cell_wire[151];							inform_R[140][6] = r_cell_wire[152];							inform_R[172][6] = r_cell_wire[153];							inform_R[141][6] = r_cell_wire[154];							inform_R[173][6] = r_cell_wire[155];							inform_R[142][6] = r_cell_wire[156];							inform_R[174][6] = r_cell_wire[157];							inform_R[143][6] = r_cell_wire[158];							inform_R[175][6] = r_cell_wire[159];							inform_R[144][6] = r_cell_wire[160];							inform_R[176][6] = r_cell_wire[161];							inform_R[145][6] = r_cell_wire[162];							inform_R[177][6] = r_cell_wire[163];							inform_R[146][6] = r_cell_wire[164];							inform_R[178][6] = r_cell_wire[165];							inform_R[147][6] = r_cell_wire[166];							inform_R[179][6] = r_cell_wire[167];							inform_R[148][6] = r_cell_wire[168];							inform_R[180][6] = r_cell_wire[169];							inform_R[149][6] = r_cell_wire[170];							inform_R[181][6] = r_cell_wire[171];							inform_R[150][6] = r_cell_wire[172];							inform_R[182][6] = r_cell_wire[173];							inform_R[151][6] = r_cell_wire[174];							inform_R[183][6] = r_cell_wire[175];							inform_R[152][6] = r_cell_wire[176];							inform_R[184][6] = r_cell_wire[177];							inform_R[153][6] = r_cell_wire[178];							inform_R[185][6] = r_cell_wire[179];							inform_R[154][6] = r_cell_wire[180];							inform_R[186][6] = r_cell_wire[181];							inform_R[155][6] = r_cell_wire[182];							inform_R[187][6] = r_cell_wire[183];							inform_R[156][6] = r_cell_wire[184];							inform_R[188][6] = r_cell_wire[185];							inform_R[157][6] = r_cell_wire[186];							inform_R[189][6] = r_cell_wire[187];							inform_R[158][6] = r_cell_wire[188];							inform_R[190][6] = r_cell_wire[189];							inform_R[159][6] = r_cell_wire[190];							inform_R[191][6] = r_cell_wire[191];							inform_R[192][6] = r_cell_wire[192];							inform_R[224][6] = r_cell_wire[193];							inform_R[193][6] = r_cell_wire[194];							inform_R[225][6] = r_cell_wire[195];							inform_R[194][6] = r_cell_wire[196];							inform_R[226][6] = r_cell_wire[197];							inform_R[195][6] = r_cell_wire[198];							inform_R[227][6] = r_cell_wire[199];							inform_R[196][6] = r_cell_wire[200];							inform_R[228][6] = r_cell_wire[201];							inform_R[197][6] = r_cell_wire[202];							inform_R[229][6] = r_cell_wire[203];							inform_R[198][6] = r_cell_wire[204];							inform_R[230][6] = r_cell_wire[205];							inform_R[199][6] = r_cell_wire[206];							inform_R[231][6] = r_cell_wire[207];							inform_R[200][6] = r_cell_wire[208];							inform_R[232][6] = r_cell_wire[209];							inform_R[201][6] = r_cell_wire[210];							inform_R[233][6] = r_cell_wire[211];							inform_R[202][6] = r_cell_wire[212];							inform_R[234][6] = r_cell_wire[213];							inform_R[203][6] = r_cell_wire[214];							inform_R[235][6] = r_cell_wire[215];							inform_R[204][6] = r_cell_wire[216];							inform_R[236][6] = r_cell_wire[217];							inform_R[205][6] = r_cell_wire[218];							inform_R[237][6] = r_cell_wire[219];							inform_R[206][6] = r_cell_wire[220];							inform_R[238][6] = r_cell_wire[221];							inform_R[207][6] = r_cell_wire[222];							inform_R[239][6] = r_cell_wire[223];							inform_R[208][6] = r_cell_wire[224];							inform_R[240][6] = r_cell_wire[225];							inform_R[209][6] = r_cell_wire[226];							inform_R[241][6] = r_cell_wire[227];							inform_R[210][6] = r_cell_wire[228];							inform_R[242][6] = r_cell_wire[229];							inform_R[211][6] = r_cell_wire[230];							inform_R[243][6] = r_cell_wire[231];							inform_R[212][6] = r_cell_wire[232];							inform_R[244][6] = r_cell_wire[233];							inform_R[213][6] = r_cell_wire[234];							inform_R[245][6] = r_cell_wire[235];							inform_R[214][6] = r_cell_wire[236];							inform_R[246][6] = r_cell_wire[237];							inform_R[215][6] = r_cell_wire[238];							inform_R[247][6] = r_cell_wire[239];							inform_R[216][6] = r_cell_wire[240];							inform_R[248][6] = r_cell_wire[241];							inform_R[217][6] = r_cell_wire[242];							inform_R[249][6] = r_cell_wire[243];							inform_R[218][6] = r_cell_wire[244];							inform_R[250][6] = r_cell_wire[245];							inform_R[219][6] = r_cell_wire[246];							inform_R[251][6] = r_cell_wire[247];							inform_R[220][6] = r_cell_wire[248];							inform_R[252][6] = r_cell_wire[249];							inform_R[221][6] = r_cell_wire[250];							inform_R[253][6] = r_cell_wire[251];							inform_R[222][6] = r_cell_wire[252];							inform_R[254][6] = r_cell_wire[253];							inform_R[223][6] = r_cell_wire[254];							inform_R[255][6] = r_cell_wire[255];							inform_R[256][6] = r_cell_wire[256];							inform_R[288][6] = r_cell_wire[257];							inform_R[257][6] = r_cell_wire[258];							inform_R[289][6] = r_cell_wire[259];							inform_R[258][6] = r_cell_wire[260];							inform_R[290][6] = r_cell_wire[261];							inform_R[259][6] = r_cell_wire[262];							inform_R[291][6] = r_cell_wire[263];							inform_R[260][6] = r_cell_wire[264];							inform_R[292][6] = r_cell_wire[265];							inform_R[261][6] = r_cell_wire[266];							inform_R[293][6] = r_cell_wire[267];							inform_R[262][6] = r_cell_wire[268];							inform_R[294][6] = r_cell_wire[269];							inform_R[263][6] = r_cell_wire[270];							inform_R[295][6] = r_cell_wire[271];							inform_R[264][6] = r_cell_wire[272];							inform_R[296][6] = r_cell_wire[273];							inform_R[265][6] = r_cell_wire[274];							inform_R[297][6] = r_cell_wire[275];							inform_R[266][6] = r_cell_wire[276];							inform_R[298][6] = r_cell_wire[277];							inform_R[267][6] = r_cell_wire[278];							inform_R[299][6] = r_cell_wire[279];							inform_R[268][6] = r_cell_wire[280];							inform_R[300][6] = r_cell_wire[281];							inform_R[269][6] = r_cell_wire[282];							inform_R[301][6] = r_cell_wire[283];							inform_R[270][6] = r_cell_wire[284];							inform_R[302][6] = r_cell_wire[285];							inform_R[271][6] = r_cell_wire[286];							inform_R[303][6] = r_cell_wire[287];							inform_R[272][6] = r_cell_wire[288];							inform_R[304][6] = r_cell_wire[289];							inform_R[273][6] = r_cell_wire[290];							inform_R[305][6] = r_cell_wire[291];							inform_R[274][6] = r_cell_wire[292];							inform_R[306][6] = r_cell_wire[293];							inform_R[275][6] = r_cell_wire[294];							inform_R[307][6] = r_cell_wire[295];							inform_R[276][6] = r_cell_wire[296];							inform_R[308][6] = r_cell_wire[297];							inform_R[277][6] = r_cell_wire[298];							inform_R[309][6] = r_cell_wire[299];							inform_R[278][6] = r_cell_wire[300];							inform_R[310][6] = r_cell_wire[301];							inform_R[279][6] = r_cell_wire[302];							inform_R[311][6] = r_cell_wire[303];							inform_R[280][6] = r_cell_wire[304];							inform_R[312][6] = r_cell_wire[305];							inform_R[281][6] = r_cell_wire[306];							inform_R[313][6] = r_cell_wire[307];							inform_R[282][6] = r_cell_wire[308];							inform_R[314][6] = r_cell_wire[309];							inform_R[283][6] = r_cell_wire[310];							inform_R[315][6] = r_cell_wire[311];							inform_R[284][6] = r_cell_wire[312];							inform_R[316][6] = r_cell_wire[313];							inform_R[285][6] = r_cell_wire[314];							inform_R[317][6] = r_cell_wire[315];							inform_R[286][6] = r_cell_wire[316];							inform_R[318][6] = r_cell_wire[317];							inform_R[287][6] = r_cell_wire[318];							inform_R[319][6] = r_cell_wire[319];							inform_R[320][6] = r_cell_wire[320];							inform_R[352][6] = r_cell_wire[321];							inform_R[321][6] = r_cell_wire[322];							inform_R[353][6] = r_cell_wire[323];							inform_R[322][6] = r_cell_wire[324];							inform_R[354][6] = r_cell_wire[325];							inform_R[323][6] = r_cell_wire[326];							inform_R[355][6] = r_cell_wire[327];							inform_R[324][6] = r_cell_wire[328];							inform_R[356][6] = r_cell_wire[329];							inform_R[325][6] = r_cell_wire[330];							inform_R[357][6] = r_cell_wire[331];							inform_R[326][6] = r_cell_wire[332];							inform_R[358][6] = r_cell_wire[333];							inform_R[327][6] = r_cell_wire[334];							inform_R[359][6] = r_cell_wire[335];							inform_R[328][6] = r_cell_wire[336];							inform_R[360][6] = r_cell_wire[337];							inform_R[329][6] = r_cell_wire[338];							inform_R[361][6] = r_cell_wire[339];							inform_R[330][6] = r_cell_wire[340];							inform_R[362][6] = r_cell_wire[341];							inform_R[331][6] = r_cell_wire[342];							inform_R[363][6] = r_cell_wire[343];							inform_R[332][6] = r_cell_wire[344];							inform_R[364][6] = r_cell_wire[345];							inform_R[333][6] = r_cell_wire[346];							inform_R[365][6] = r_cell_wire[347];							inform_R[334][6] = r_cell_wire[348];							inform_R[366][6] = r_cell_wire[349];							inform_R[335][6] = r_cell_wire[350];							inform_R[367][6] = r_cell_wire[351];							inform_R[336][6] = r_cell_wire[352];							inform_R[368][6] = r_cell_wire[353];							inform_R[337][6] = r_cell_wire[354];							inform_R[369][6] = r_cell_wire[355];							inform_R[338][6] = r_cell_wire[356];							inform_R[370][6] = r_cell_wire[357];							inform_R[339][6] = r_cell_wire[358];							inform_R[371][6] = r_cell_wire[359];							inform_R[340][6] = r_cell_wire[360];							inform_R[372][6] = r_cell_wire[361];							inform_R[341][6] = r_cell_wire[362];							inform_R[373][6] = r_cell_wire[363];							inform_R[342][6] = r_cell_wire[364];							inform_R[374][6] = r_cell_wire[365];							inform_R[343][6] = r_cell_wire[366];							inform_R[375][6] = r_cell_wire[367];							inform_R[344][6] = r_cell_wire[368];							inform_R[376][6] = r_cell_wire[369];							inform_R[345][6] = r_cell_wire[370];							inform_R[377][6] = r_cell_wire[371];							inform_R[346][6] = r_cell_wire[372];							inform_R[378][6] = r_cell_wire[373];							inform_R[347][6] = r_cell_wire[374];							inform_R[379][6] = r_cell_wire[375];							inform_R[348][6] = r_cell_wire[376];							inform_R[380][6] = r_cell_wire[377];							inform_R[349][6] = r_cell_wire[378];							inform_R[381][6] = r_cell_wire[379];							inform_R[350][6] = r_cell_wire[380];							inform_R[382][6] = r_cell_wire[381];							inform_R[351][6] = r_cell_wire[382];							inform_R[383][6] = r_cell_wire[383];							inform_R[384][6] = r_cell_wire[384];							inform_R[416][6] = r_cell_wire[385];							inform_R[385][6] = r_cell_wire[386];							inform_R[417][6] = r_cell_wire[387];							inform_R[386][6] = r_cell_wire[388];							inform_R[418][6] = r_cell_wire[389];							inform_R[387][6] = r_cell_wire[390];							inform_R[419][6] = r_cell_wire[391];							inform_R[388][6] = r_cell_wire[392];							inform_R[420][6] = r_cell_wire[393];							inform_R[389][6] = r_cell_wire[394];							inform_R[421][6] = r_cell_wire[395];							inform_R[390][6] = r_cell_wire[396];							inform_R[422][6] = r_cell_wire[397];							inform_R[391][6] = r_cell_wire[398];							inform_R[423][6] = r_cell_wire[399];							inform_R[392][6] = r_cell_wire[400];							inform_R[424][6] = r_cell_wire[401];							inform_R[393][6] = r_cell_wire[402];							inform_R[425][6] = r_cell_wire[403];							inform_R[394][6] = r_cell_wire[404];							inform_R[426][6] = r_cell_wire[405];							inform_R[395][6] = r_cell_wire[406];							inform_R[427][6] = r_cell_wire[407];							inform_R[396][6] = r_cell_wire[408];							inform_R[428][6] = r_cell_wire[409];							inform_R[397][6] = r_cell_wire[410];							inform_R[429][6] = r_cell_wire[411];							inform_R[398][6] = r_cell_wire[412];							inform_R[430][6] = r_cell_wire[413];							inform_R[399][6] = r_cell_wire[414];							inform_R[431][6] = r_cell_wire[415];							inform_R[400][6] = r_cell_wire[416];							inform_R[432][6] = r_cell_wire[417];							inform_R[401][6] = r_cell_wire[418];							inform_R[433][6] = r_cell_wire[419];							inform_R[402][6] = r_cell_wire[420];							inform_R[434][6] = r_cell_wire[421];							inform_R[403][6] = r_cell_wire[422];							inform_R[435][6] = r_cell_wire[423];							inform_R[404][6] = r_cell_wire[424];							inform_R[436][6] = r_cell_wire[425];							inform_R[405][6] = r_cell_wire[426];							inform_R[437][6] = r_cell_wire[427];							inform_R[406][6] = r_cell_wire[428];							inform_R[438][6] = r_cell_wire[429];							inform_R[407][6] = r_cell_wire[430];							inform_R[439][6] = r_cell_wire[431];							inform_R[408][6] = r_cell_wire[432];							inform_R[440][6] = r_cell_wire[433];							inform_R[409][6] = r_cell_wire[434];							inform_R[441][6] = r_cell_wire[435];							inform_R[410][6] = r_cell_wire[436];							inform_R[442][6] = r_cell_wire[437];							inform_R[411][6] = r_cell_wire[438];							inform_R[443][6] = r_cell_wire[439];							inform_R[412][6] = r_cell_wire[440];							inform_R[444][6] = r_cell_wire[441];							inform_R[413][6] = r_cell_wire[442];							inform_R[445][6] = r_cell_wire[443];							inform_R[414][6] = r_cell_wire[444];							inform_R[446][6] = r_cell_wire[445];							inform_R[415][6] = r_cell_wire[446];							inform_R[447][6] = r_cell_wire[447];							inform_R[448][6] = r_cell_wire[448];							inform_R[480][6] = r_cell_wire[449];							inform_R[449][6] = r_cell_wire[450];							inform_R[481][6] = r_cell_wire[451];							inform_R[450][6] = r_cell_wire[452];							inform_R[482][6] = r_cell_wire[453];							inform_R[451][6] = r_cell_wire[454];							inform_R[483][6] = r_cell_wire[455];							inform_R[452][6] = r_cell_wire[456];							inform_R[484][6] = r_cell_wire[457];							inform_R[453][6] = r_cell_wire[458];							inform_R[485][6] = r_cell_wire[459];							inform_R[454][6] = r_cell_wire[460];							inform_R[486][6] = r_cell_wire[461];							inform_R[455][6] = r_cell_wire[462];							inform_R[487][6] = r_cell_wire[463];							inform_R[456][6] = r_cell_wire[464];							inform_R[488][6] = r_cell_wire[465];							inform_R[457][6] = r_cell_wire[466];							inform_R[489][6] = r_cell_wire[467];							inform_R[458][6] = r_cell_wire[468];							inform_R[490][6] = r_cell_wire[469];							inform_R[459][6] = r_cell_wire[470];							inform_R[491][6] = r_cell_wire[471];							inform_R[460][6] = r_cell_wire[472];							inform_R[492][6] = r_cell_wire[473];							inform_R[461][6] = r_cell_wire[474];							inform_R[493][6] = r_cell_wire[475];							inform_R[462][6] = r_cell_wire[476];							inform_R[494][6] = r_cell_wire[477];							inform_R[463][6] = r_cell_wire[478];							inform_R[495][6] = r_cell_wire[479];							inform_R[464][6] = r_cell_wire[480];							inform_R[496][6] = r_cell_wire[481];							inform_R[465][6] = r_cell_wire[482];							inform_R[497][6] = r_cell_wire[483];							inform_R[466][6] = r_cell_wire[484];							inform_R[498][6] = r_cell_wire[485];							inform_R[467][6] = r_cell_wire[486];							inform_R[499][6] = r_cell_wire[487];							inform_R[468][6] = r_cell_wire[488];							inform_R[500][6] = r_cell_wire[489];							inform_R[469][6] = r_cell_wire[490];							inform_R[501][6] = r_cell_wire[491];							inform_R[470][6] = r_cell_wire[492];							inform_R[502][6] = r_cell_wire[493];							inform_R[471][6] = r_cell_wire[494];							inform_R[503][6] = r_cell_wire[495];							inform_R[472][6] = r_cell_wire[496];							inform_R[504][6] = r_cell_wire[497];							inform_R[473][6] = r_cell_wire[498];							inform_R[505][6] = r_cell_wire[499];							inform_R[474][6] = r_cell_wire[500];							inform_R[506][6] = r_cell_wire[501];							inform_R[475][6] = r_cell_wire[502];							inform_R[507][6] = r_cell_wire[503];							inform_R[476][6] = r_cell_wire[504];							inform_R[508][6] = r_cell_wire[505];							inform_R[477][6] = r_cell_wire[506];							inform_R[509][6] = r_cell_wire[507];							inform_R[478][6] = r_cell_wire[508];							inform_R[510][6] = r_cell_wire[509];							inform_R[479][6] = r_cell_wire[510];							inform_R[511][6] = r_cell_wire[511];							inform_R[512][6] = r_cell_wire[512];							inform_R[544][6] = r_cell_wire[513];							inform_R[513][6] = r_cell_wire[514];							inform_R[545][6] = r_cell_wire[515];							inform_R[514][6] = r_cell_wire[516];							inform_R[546][6] = r_cell_wire[517];							inform_R[515][6] = r_cell_wire[518];							inform_R[547][6] = r_cell_wire[519];							inform_R[516][6] = r_cell_wire[520];							inform_R[548][6] = r_cell_wire[521];							inform_R[517][6] = r_cell_wire[522];							inform_R[549][6] = r_cell_wire[523];							inform_R[518][6] = r_cell_wire[524];							inform_R[550][6] = r_cell_wire[525];							inform_R[519][6] = r_cell_wire[526];							inform_R[551][6] = r_cell_wire[527];							inform_R[520][6] = r_cell_wire[528];							inform_R[552][6] = r_cell_wire[529];							inform_R[521][6] = r_cell_wire[530];							inform_R[553][6] = r_cell_wire[531];							inform_R[522][6] = r_cell_wire[532];							inform_R[554][6] = r_cell_wire[533];							inform_R[523][6] = r_cell_wire[534];							inform_R[555][6] = r_cell_wire[535];							inform_R[524][6] = r_cell_wire[536];							inform_R[556][6] = r_cell_wire[537];							inform_R[525][6] = r_cell_wire[538];							inform_R[557][6] = r_cell_wire[539];							inform_R[526][6] = r_cell_wire[540];							inform_R[558][6] = r_cell_wire[541];							inform_R[527][6] = r_cell_wire[542];							inform_R[559][6] = r_cell_wire[543];							inform_R[528][6] = r_cell_wire[544];							inform_R[560][6] = r_cell_wire[545];							inform_R[529][6] = r_cell_wire[546];							inform_R[561][6] = r_cell_wire[547];							inform_R[530][6] = r_cell_wire[548];							inform_R[562][6] = r_cell_wire[549];							inform_R[531][6] = r_cell_wire[550];							inform_R[563][6] = r_cell_wire[551];							inform_R[532][6] = r_cell_wire[552];							inform_R[564][6] = r_cell_wire[553];							inform_R[533][6] = r_cell_wire[554];							inform_R[565][6] = r_cell_wire[555];							inform_R[534][6] = r_cell_wire[556];							inform_R[566][6] = r_cell_wire[557];							inform_R[535][6] = r_cell_wire[558];							inform_R[567][6] = r_cell_wire[559];							inform_R[536][6] = r_cell_wire[560];							inform_R[568][6] = r_cell_wire[561];							inform_R[537][6] = r_cell_wire[562];							inform_R[569][6] = r_cell_wire[563];							inform_R[538][6] = r_cell_wire[564];							inform_R[570][6] = r_cell_wire[565];							inform_R[539][6] = r_cell_wire[566];							inform_R[571][6] = r_cell_wire[567];							inform_R[540][6] = r_cell_wire[568];							inform_R[572][6] = r_cell_wire[569];							inform_R[541][6] = r_cell_wire[570];							inform_R[573][6] = r_cell_wire[571];							inform_R[542][6] = r_cell_wire[572];							inform_R[574][6] = r_cell_wire[573];							inform_R[543][6] = r_cell_wire[574];							inform_R[575][6] = r_cell_wire[575];							inform_R[576][6] = r_cell_wire[576];							inform_R[608][6] = r_cell_wire[577];							inform_R[577][6] = r_cell_wire[578];							inform_R[609][6] = r_cell_wire[579];							inform_R[578][6] = r_cell_wire[580];							inform_R[610][6] = r_cell_wire[581];							inform_R[579][6] = r_cell_wire[582];							inform_R[611][6] = r_cell_wire[583];							inform_R[580][6] = r_cell_wire[584];							inform_R[612][6] = r_cell_wire[585];							inform_R[581][6] = r_cell_wire[586];							inform_R[613][6] = r_cell_wire[587];							inform_R[582][6] = r_cell_wire[588];							inform_R[614][6] = r_cell_wire[589];							inform_R[583][6] = r_cell_wire[590];							inform_R[615][6] = r_cell_wire[591];							inform_R[584][6] = r_cell_wire[592];							inform_R[616][6] = r_cell_wire[593];							inform_R[585][6] = r_cell_wire[594];							inform_R[617][6] = r_cell_wire[595];							inform_R[586][6] = r_cell_wire[596];							inform_R[618][6] = r_cell_wire[597];							inform_R[587][6] = r_cell_wire[598];							inform_R[619][6] = r_cell_wire[599];							inform_R[588][6] = r_cell_wire[600];							inform_R[620][6] = r_cell_wire[601];							inform_R[589][6] = r_cell_wire[602];							inform_R[621][6] = r_cell_wire[603];							inform_R[590][6] = r_cell_wire[604];							inform_R[622][6] = r_cell_wire[605];							inform_R[591][6] = r_cell_wire[606];							inform_R[623][6] = r_cell_wire[607];							inform_R[592][6] = r_cell_wire[608];							inform_R[624][6] = r_cell_wire[609];							inform_R[593][6] = r_cell_wire[610];							inform_R[625][6] = r_cell_wire[611];							inform_R[594][6] = r_cell_wire[612];							inform_R[626][6] = r_cell_wire[613];							inform_R[595][6] = r_cell_wire[614];							inform_R[627][6] = r_cell_wire[615];							inform_R[596][6] = r_cell_wire[616];							inform_R[628][6] = r_cell_wire[617];							inform_R[597][6] = r_cell_wire[618];							inform_R[629][6] = r_cell_wire[619];							inform_R[598][6] = r_cell_wire[620];							inform_R[630][6] = r_cell_wire[621];							inform_R[599][6] = r_cell_wire[622];							inform_R[631][6] = r_cell_wire[623];							inform_R[600][6] = r_cell_wire[624];							inform_R[632][6] = r_cell_wire[625];							inform_R[601][6] = r_cell_wire[626];							inform_R[633][6] = r_cell_wire[627];							inform_R[602][6] = r_cell_wire[628];							inform_R[634][6] = r_cell_wire[629];							inform_R[603][6] = r_cell_wire[630];							inform_R[635][6] = r_cell_wire[631];							inform_R[604][6] = r_cell_wire[632];							inform_R[636][6] = r_cell_wire[633];							inform_R[605][6] = r_cell_wire[634];							inform_R[637][6] = r_cell_wire[635];							inform_R[606][6] = r_cell_wire[636];							inform_R[638][6] = r_cell_wire[637];							inform_R[607][6] = r_cell_wire[638];							inform_R[639][6] = r_cell_wire[639];							inform_R[640][6] = r_cell_wire[640];							inform_R[672][6] = r_cell_wire[641];							inform_R[641][6] = r_cell_wire[642];							inform_R[673][6] = r_cell_wire[643];							inform_R[642][6] = r_cell_wire[644];							inform_R[674][6] = r_cell_wire[645];							inform_R[643][6] = r_cell_wire[646];							inform_R[675][6] = r_cell_wire[647];							inform_R[644][6] = r_cell_wire[648];							inform_R[676][6] = r_cell_wire[649];							inform_R[645][6] = r_cell_wire[650];							inform_R[677][6] = r_cell_wire[651];							inform_R[646][6] = r_cell_wire[652];							inform_R[678][6] = r_cell_wire[653];							inform_R[647][6] = r_cell_wire[654];							inform_R[679][6] = r_cell_wire[655];							inform_R[648][6] = r_cell_wire[656];							inform_R[680][6] = r_cell_wire[657];							inform_R[649][6] = r_cell_wire[658];							inform_R[681][6] = r_cell_wire[659];							inform_R[650][6] = r_cell_wire[660];							inform_R[682][6] = r_cell_wire[661];							inform_R[651][6] = r_cell_wire[662];							inform_R[683][6] = r_cell_wire[663];							inform_R[652][6] = r_cell_wire[664];							inform_R[684][6] = r_cell_wire[665];							inform_R[653][6] = r_cell_wire[666];							inform_R[685][6] = r_cell_wire[667];							inform_R[654][6] = r_cell_wire[668];							inform_R[686][6] = r_cell_wire[669];							inform_R[655][6] = r_cell_wire[670];							inform_R[687][6] = r_cell_wire[671];							inform_R[656][6] = r_cell_wire[672];							inform_R[688][6] = r_cell_wire[673];							inform_R[657][6] = r_cell_wire[674];							inform_R[689][6] = r_cell_wire[675];							inform_R[658][6] = r_cell_wire[676];							inform_R[690][6] = r_cell_wire[677];							inform_R[659][6] = r_cell_wire[678];							inform_R[691][6] = r_cell_wire[679];							inform_R[660][6] = r_cell_wire[680];							inform_R[692][6] = r_cell_wire[681];							inform_R[661][6] = r_cell_wire[682];							inform_R[693][6] = r_cell_wire[683];							inform_R[662][6] = r_cell_wire[684];							inform_R[694][6] = r_cell_wire[685];							inform_R[663][6] = r_cell_wire[686];							inform_R[695][6] = r_cell_wire[687];							inform_R[664][6] = r_cell_wire[688];							inform_R[696][6] = r_cell_wire[689];							inform_R[665][6] = r_cell_wire[690];							inform_R[697][6] = r_cell_wire[691];							inform_R[666][6] = r_cell_wire[692];							inform_R[698][6] = r_cell_wire[693];							inform_R[667][6] = r_cell_wire[694];							inform_R[699][6] = r_cell_wire[695];							inform_R[668][6] = r_cell_wire[696];							inform_R[700][6] = r_cell_wire[697];							inform_R[669][6] = r_cell_wire[698];							inform_R[701][6] = r_cell_wire[699];							inform_R[670][6] = r_cell_wire[700];							inform_R[702][6] = r_cell_wire[701];							inform_R[671][6] = r_cell_wire[702];							inform_R[703][6] = r_cell_wire[703];							inform_R[704][6] = r_cell_wire[704];							inform_R[736][6] = r_cell_wire[705];							inform_R[705][6] = r_cell_wire[706];							inform_R[737][6] = r_cell_wire[707];							inform_R[706][6] = r_cell_wire[708];							inform_R[738][6] = r_cell_wire[709];							inform_R[707][6] = r_cell_wire[710];							inform_R[739][6] = r_cell_wire[711];							inform_R[708][6] = r_cell_wire[712];							inform_R[740][6] = r_cell_wire[713];							inform_R[709][6] = r_cell_wire[714];							inform_R[741][6] = r_cell_wire[715];							inform_R[710][6] = r_cell_wire[716];							inform_R[742][6] = r_cell_wire[717];							inform_R[711][6] = r_cell_wire[718];							inform_R[743][6] = r_cell_wire[719];							inform_R[712][6] = r_cell_wire[720];							inform_R[744][6] = r_cell_wire[721];							inform_R[713][6] = r_cell_wire[722];							inform_R[745][6] = r_cell_wire[723];							inform_R[714][6] = r_cell_wire[724];							inform_R[746][6] = r_cell_wire[725];							inform_R[715][6] = r_cell_wire[726];							inform_R[747][6] = r_cell_wire[727];							inform_R[716][6] = r_cell_wire[728];							inform_R[748][6] = r_cell_wire[729];							inform_R[717][6] = r_cell_wire[730];							inform_R[749][6] = r_cell_wire[731];							inform_R[718][6] = r_cell_wire[732];							inform_R[750][6] = r_cell_wire[733];							inform_R[719][6] = r_cell_wire[734];							inform_R[751][6] = r_cell_wire[735];							inform_R[720][6] = r_cell_wire[736];							inform_R[752][6] = r_cell_wire[737];							inform_R[721][6] = r_cell_wire[738];							inform_R[753][6] = r_cell_wire[739];							inform_R[722][6] = r_cell_wire[740];							inform_R[754][6] = r_cell_wire[741];							inform_R[723][6] = r_cell_wire[742];							inform_R[755][6] = r_cell_wire[743];							inform_R[724][6] = r_cell_wire[744];							inform_R[756][6] = r_cell_wire[745];							inform_R[725][6] = r_cell_wire[746];							inform_R[757][6] = r_cell_wire[747];							inform_R[726][6] = r_cell_wire[748];							inform_R[758][6] = r_cell_wire[749];							inform_R[727][6] = r_cell_wire[750];							inform_R[759][6] = r_cell_wire[751];							inform_R[728][6] = r_cell_wire[752];							inform_R[760][6] = r_cell_wire[753];							inform_R[729][6] = r_cell_wire[754];							inform_R[761][6] = r_cell_wire[755];							inform_R[730][6] = r_cell_wire[756];							inform_R[762][6] = r_cell_wire[757];							inform_R[731][6] = r_cell_wire[758];							inform_R[763][6] = r_cell_wire[759];							inform_R[732][6] = r_cell_wire[760];							inform_R[764][6] = r_cell_wire[761];							inform_R[733][6] = r_cell_wire[762];							inform_R[765][6] = r_cell_wire[763];							inform_R[734][6] = r_cell_wire[764];							inform_R[766][6] = r_cell_wire[765];							inform_R[735][6] = r_cell_wire[766];							inform_R[767][6] = r_cell_wire[767];							inform_R[768][6] = r_cell_wire[768];							inform_R[800][6] = r_cell_wire[769];							inform_R[769][6] = r_cell_wire[770];							inform_R[801][6] = r_cell_wire[771];							inform_R[770][6] = r_cell_wire[772];							inform_R[802][6] = r_cell_wire[773];							inform_R[771][6] = r_cell_wire[774];							inform_R[803][6] = r_cell_wire[775];							inform_R[772][6] = r_cell_wire[776];							inform_R[804][6] = r_cell_wire[777];							inform_R[773][6] = r_cell_wire[778];							inform_R[805][6] = r_cell_wire[779];							inform_R[774][6] = r_cell_wire[780];							inform_R[806][6] = r_cell_wire[781];							inform_R[775][6] = r_cell_wire[782];							inform_R[807][6] = r_cell_wire[783];							inform_R[776][6] = r_cell_wire[784];							inform_R[808][6] = r_cell_wire[785];							inform_R[777][6] = r_cell_wire[786];							inform_R[809][6] = r_cell_wire[787];							inform_R[778][6] = r_cell_wire[788];							inform_R[810][6] = r_cell_wire[789];							inform_R[779][6] = r_cell_wire[790];							inform_R[811][6] = r_cell_wire[791];							inform_R[780][6] = r_cell_wire[792];							inform_R[812][6] = r_cell_wire[793];							inform_R[781][6] = r_cell_wire[794];							inform_R[813][6] = r_cell_wire[795];							inform_R[782][6] = r_cell_wire[796];							inform_R[814][6] = r_cell_wire[797];							inform_R[783][6] = r_cell_wire[798];							inform_R[815][6] = r_cell_wire[799];							inform_R[784][6] = r_cell_wire[800];							inform_R[816][6] = r_cell_wire[801];							inform_R[785][6] = r_cell_wire[802];							inform_R[817][6] = r_cell_wire[803];							inform_R[786][6] = r_cell_wire[804];							inform_R[818][6] = r_cell_wire[805];							inform_R[787][6] = r_cell_wire[806];							inform_R[819][6] = r_cell_wire[807];							inform_R[788][6] = r_cell_wire[808];							inform_R[820][6] = r_cell_wire[809];							inform_R[789][6] = r_cell_wire[810];							inform_R[821][6] = r_cell_wire[811];							inform_R[790][6] = r_cell_wire[812];							inform_R[822][6] = r_cell_wire[813];							inform_R[791][6] = r_cell_wire[814];							inform_R[823][6] = r_cell_wire[815];							inform_R[792][6] = r_cell_wire[816];							inform_R[824][6] = r_cell_wire[817];							inform_R[793][6] = r_cell_wire[818];							inform_R[825][6] = r_cell_wire[819];							inform_R[794][6] = r_cell_wire[820];							inform_R[826][6] = r_cell_wire[821];							inform_R[795][6] = r_cell_wire[822];							inform_R[827][6] = r_cell_wire[823];							inform_R[796][6] = r_cell_wire[824];							inform_R[828][6] = r_cell_wire[825];							inform_R[797][6] = r_cell_wire[826];							inform_R[829][6] = r_cell_wire[827];							inform_R[798][6] = r_cell_wire[828];							inform_R[830][6] = r_cell_wire[829];							inform_R[799][6] = r_cell_wire[830];							inform_R[831][6] = r_cell_wire[831];							inform_R[832][6] = r_cell_wire[832];							inform_R[864][6] = r_cell_wire[833];							inform_R[833][6] = r_cell_wire[834];							inform_R[865][6] = r_cell_wire[835];							inform_R[834][6] = r_cell_wire[836];							inform_R[866][6] = r_cell_wire[837];							inform_R[835][6] = r_cell_wire[838];							inform_R[867][6] = r_cell_wire[839];							inform_R[836][6] = r_cell_wire[840];							inform_R[868][6] = r_cell_wire[841];							inform_R[837][6] = r_cell_wire[842];							inform_R[869][6] = r_cell_wire[843];							inform_R[838][6] = r_cell_wire[844];							inform_R[870][6] = r_cell_wire[845];							inform_R[839][6] = r_cell_wire[846];							inform_R[871][6] = r_cell_wire[847];							inform_R[840][6] = r_cell_wire[848];							inform_R[872][6] = r_cell_wire[849];							inform_R[841][6] = r_cell_wire[850];							inform_R[873][6] = r_cell_wire[851];							inform_R[842][6] = r_cell_wire[852];							inform_R[874][6] = r_cell_wire[853];							inform_R[843][6] = r_cell_wire[854];							inform_R[875][6] = r_cell_wire[855];							inform_R[844][6] = r_cell_wire[856];							inform_R[876][6] = r_cell_wire[857];							inform_R[845][6] = r_cell_wire[858];							inform_R[877][6] = r_cell_wire[859];							inform_R[846][6] = r_cell_wire[860];							inform_R[878][6] = r_cell_wire[861];							inform_R[847][6] = r_cell_wire[862];							inform_R[879][6] = r_cell_wire[863];							inform_R[848][6] = r_cell_wire[864];							inform_R[880][6] = r_cell_wire[865];							inform_R[849][6] = r_cell_wire[866];							inform_R[881][6] = r_cell_wire[867];							inform_R[850][6] = r_cell_wire[868];							inform_R[882][6] = r_cell_wire[869];							inform_R[851][6] = r_cell_wire[870];							inform_R[883][6] = r_cell_wire[871];							inform_R[852][6] = r_cell_wire[872];							inform_R[884][6] = r_cell_wire[873];							inform_R[853][6] = r_cell_wire[874];							inform_R[885][6] = r_cell_wire[875];							inform_R[854][6] = r_cell_wire[876];							inform_R[886][6] = r_cell_wire[877];							inform_R[855][6] = r_cell_wire[878];							inform_R[887][6] = r_cell_wire[879];							inform_R[856][6] = r_cell_wire[880];							inform_R[888][6] = r_cell_wire[881];							inform_R[857][6] = r_cell_wire[882];							inform_R[889][6] = r_cell_wire[883];							inform_R[858][6] = r_cell_wire[884];							inform_R[890][6] = r_cell_wire[885];							inform_R[859][6] = r_cell_wire[886];							inform_R[891][6] = r_cell_wire[887];							inform_R[860][6] = r_cell_wire[888];							inform_R[892][6] = r_cell_wire[889];							inform_R[861][6] = r_cell_wire[890];							inform_R[893][6] = r_cell_wire[891];							inform_R[862][6] = r_cell_wire[892];							inform_R[894][6] = r_cell_wire[893];							inform_R[863][6] = r_cell_wire[894];							inform_R[895][6] = r_cell_wire[895];							inform_R[896][6] = r_cell_wire[896];							inform_R[928][6] = r_cell_wire[897];							inform_R[897][6] = r_cell_wire[898];							inform_R[929][6] = r_cell_wire[899];							inform_R[898][6] = r_cell_wire[900];							inform_R[930][6] = r_cell_wire[901];							inform_R[899][6] = r_cell_wire[902];							inform_R[931][6] = r_cell_wire[903];							inform_R[900][6] = r_cell_wire[904];							inform_R[932][6] = r_cell_wire[905];							inform_R[901][6] = r_cell_wire[906];							inform_R[933][6] = r_cell_wire[907];							inform_R[902][6] = r_cell_wire[908];							inform_R[934][6] = r_cell_wire[909];							inform_R[903][6] = r_cell_wire[910];							inform_R[935][6] = r_cell_wire[911];							inform_R[904][6] = r_cell_wire[912];							inform_R[936][6] = r_cell_wire[913];							inform_R[905][6] = r_cell_wire[914];							inform_R[937][6] = r_cell_wire[915];							inform_R[906][6] = r_cell_wire[916];							inform_R[938][6] = r_cell_wire[917];							inform_R[907][6] = r_cell_wire[918];							inform_R[939][6] = r_cell_wire[919];							inform_R[908][6] = r_cell_wire[920];							inform_R[940][6] = r_cell_wire[921];							inform_R[909][6] = r_cell_wire[922];							inform_R[941][6] = r_cell_wire[923];							inform_R[910][6] = r_cell_wire[924];							inform_R[942][6] = r_cell_wire[925];							inform_R[911][6] = r_cell_wire[926];							inform_R[943][6] = r_cell_wire[927];							inform_R[912][6] = r_cell_wire[928];							inform_R[944][6] = r_cell_wire[929];							inform_R[913][6] = r_cell_wire[930];							inform_R[945][6] = r_cell_wire[931];							inform_R[914][6] = r_cell_wire[932];							inform_R[946][6] = r_cell_wire[933];							inform_R[915][6] = r_cell_wire[934];							inform_R[947][6] = r_cell_wire[935];							inform_R[916][6] = r_cell_wire[936];							inform_R[948][6] = r_cell_wire[937];							inform_R[917][6] = r_cell_wire[938];							inform_R[949][6] = r_cell_wire[939];							inform_R[918][6] = r_cell_wire[940];							inform_R[950][6] = r_cell_wire[941];							inform_R[919][6] = r_cell_wire[942];							inform_R[951][6] = r_cell_wire[943];							inform_R[920][6] = r_cell_wire[944];							inform_R[952][6] = r_cell_wire[945];							inform_R[921][6] = r_cell_wire[946];							inform_R[953][6] = r_cell_wire[947];							inform_R[922][6] = r_cell_wire[948];							inform_R[954][6] = r_cell_wire[949];							inform_R[923][6] = r_cell_wire[950];							inform_R[955][6] = r_cell_wire[951];							inform_R[924][6] = r_cell_wire[952];							inform_R[956][6] = r_cell_wire[953];							inform_R[925][6] = r_cell_wire[954];							inform_R[957][6] = r_cell_wire[955];							inform_R[926][6] = r_cell_wire[956];							inform_R[958][6] = r_cell_wire[957];							inform_R[927][6] = r_cell_wire[958];							inform_R[959][6] = r_cell_wire[959];							inform_R[960][6] = r_cell_wire[960];							inform_R[992][6] = r_cell_wire[961];							inform_R[961][6] = r_cell_wire[962];							inform_R[993][6] = r_cell_wire[963];							inform_R[962][6] = r_cell_wire[964];							inform_R[994][6] = r_cell_wire[965];							inform_R[963][6] = r_cell_wire[966];							inform_R[995][6] = r_cell_wire[967];							inform_R[964][6] = r_cell_wire[968];							inform_R[996][6] = r_cell_wire[969];							inform_R[965][6] = r_cell_wire[970];							inform_R[997][6] = r_cell_wire[971];							inform_R[966][6] = r_cell_wire[972];							inform_R[998][6] = r_cell_wire[973];							inform_R[967][6] = r_cell_wire[974];							inform_R[999][6] = r_cell_wire[975];							inform_R[968][6] = r_cell_wire[976];							inform_R[1000][6] = r_cell_wire[977];							inform_R[969][6] = r_cell_wire[978];							inform_R[1001][6] = r_cell_wire[979];							inform_R[970][6] = r_cell_wire[980];							inform_R[1002][6] = r_cell_wire[981];							inform_R[971][6] = r_cell_wire[982];							inform_R[1003][6] = r_cell_wire[983];							inform_R[972][6] = r_cell_wire[984];							inform_R[1004][6] = r_cell_wire[985];							inform_R[973][6] = r_cell_wire[986];							inform_R[1005][6] = r_cell_wire[987];							inform_R[974][6] = r_cell_wire[988];							inform_R[1006][6] = r_cell_wire[989];							inform_R[975][6] = r_cell_wire[990];							inform_R[1007][6] = r_cell_wire[991];							inform_R[976][6] = r_cell_wire[992];							inform_R[1008][6] = r_cell_wire[993];							inform_R[977][6] = r_cell_wire[994];							inform_R[1009][6] = r_cell_wire[995];							inform_R[978][6] = r_cell_wire[996];							inform_R[1010][6] = r_cell_wire[997];							inform_R[979][6] = r_cell_wire[998];							inform_R[1011][6] = r_cell_wire[999];							inform_R[980][6] = r_cell_wire[1000];							inform_R[1012][6] = r_cell_wire[1001];							inform_R[981][6] = r_cell_wire[1002];							inform_R[1013][6] = r_cell_wire[1003];							inform_R[982][6] = r_cell_wire[1004];							inform_R[1014][6] = r_cell_wire[1005];							inform_R[983][6] = r_cell_wire[1006];							inform_R[1015][6] = r_cell_wire[1007];							inform_R[984][6] = r_cell_wire[1008];							inform_R[1016][6] = r_cell_wire[1009];							inform_R[985][6] = r_cell_wire[1010];							inform_R[1017][6] = r_cell_wire[1011];							inform_R[986][6] = r_cell_wire[1012];							inform_R[1018][6] = r_cell_wire[1013];							inform_R[987][6] = r_cell_wire[1014];							inform_R[1019][6] = r_cell_wire[1015];							inform_R[988][6] = r_cell_wire[1016];							inform_R[1020][6] = r_cell_wire[1017];							inform_R[989][6] = r_cell_wire[1018];							inform_R[1021][6] = r_cell_wire[1019];							inform_R[990][6] = r_cell_wire[1020];							inform_R[1022][6] = r_cell_wire[1021];							inform_R[991][6] = r_cell_wire[1022];							inform_R[1023][6] = r_cell_wire[1023];							inform_L[0][5] = l_cell_wire[0];							inform_L[32][5] = l_cell_wire[1];							inform_L[1][5] = l_cell_wire[2];							inform_L[33][5] = l_cell_wire[3];							inform_L[2][5] = l_cell_wire[4];							inform_L[34][5] = l_cell_wire[5];							inform_L[3][5] = l_cell_wire[6];							inform_L[35][5] = l_cell_wire[7];							inform_L[4][5] = l_cell_wire[8];							inform_L[36][5] = l_cell_wire[9];							inform_L[5][5] = l_cell_wire[10];							inform_L[37][5] = l_cell_wire[11];							inform_L[6][5] = l_cell_wire[12];							inform_L[38][5] = l_cell_wire[13];							inform_L[7][5] = l_cell_wire[14];							inform_L[39][5] = l_cell_wire[15];							inform_L[8][5] = l_cell_wire[16];							inform_L[40][5] = l_cell_wire[17];							inform_L[9][5] = l_cell_wire[18];							inform_L[41][5] = l_cell_wire[19];							inform_L[10][5] = l_cell_wire[20];							inform_L[42][5] = l_cell_wire[21];							inform_L[11][5] = l_cell_wire[22];							inform_L[43][5] = l_cell_wire[23];							inform_L[12][5] = l_cell_wire[24];							inform_L[44][5] = l_cell_wire[25];							inform_L[13][5] = l_cell_wire[26];							inform_L[45][5] = l_cell_wire[27];							inform_L[14][5] = l_cell_wire[28];							inform_L[46][5] = l_cell_wire[29];							inform_L[15][5] = l_cell_wire[30];							inform_L[47][5] = l_cell_wire[31];							inform_L[16][5] = l_cell_wire[32];							inform_L[48][5] = l_cell_wire[33];							inform_L[17][5] = l_cell_wire[34];							inform_L[49][5] = l_cell_wire[35];							inform_L[18][5] = l_cell_wire[36];							inform_L[50][5] = l_cell_wire[37];							inform_L[19][5] = l_cell_wire[38];							inform_L[51][5] = l_cell_wire[39];							inform_L[20][5] = l_cell_wire[40];							inform_L[52][5] = l_cell_wire[41];							inform_L[21][5] = l_cell_wire[42];							inform_L[53][5] = l_cell_wire[43];							inform_L[22][5] = l_cell_wire[44];							inform_L[54][5] = l_cell_wire[45];							inform_L[23][5] = l_cell_wire[46];							inform_L[55][5] = l_cell_wire[47];							inform_L[24][5] = l_cell_wire[48];							inform_L[56][5] = l_cell_wire[49];							inform_L[25][5] = l_cell_wire[50];							inform_L[57][5] = l_cell_wire[51];							inform_L[26][5] = l_cell_wire[52];							inform_L[58][5] = l_cell_wire[53];							inform_L[27][5] = l_cell_wire[54];							inform_L[59][5] = l_cell_wire[55];							inform_L[28][5] = l_cell_wire[56];							inform_L[60][5] = l_cell_wire[57];							inform_L[29][5] = l_cell_wire[58];							inform_L[61][5] = l_cell_wire[59];							inform_L[30][5] = l_cell_wire[60];							inform_L[62][5] = l_cell_wire[61];							inform_L[31][5] = l_cell_wire[62];							inform_L[63][5] = l_cell_wire[63];							inform_L[64][5] = l_cell_wire[64];							inform_L[96][5] = l_cell_wire[65];							inform_L[65][5] = l_cell_wire[66];							inform_L[97][5] = l_cell_wire[67];							inform_L[66][5] = l_cell_wire[68];							inform_L[98][5] = l_cell_wire[69];							inform_L[67][5] = l_cell_wire[70];							inform_L[99][5] = l_cell_wire[71];							inform_L[68][5] = l_cell_wire[72];							inform_L[100][5] = l_cell_wire[73];							inform_L[69][5] = l_cell_wire[74];							inform_L[101][5] = l_cell_wire[75];							inform_L[70][5] = l_cell_wire[76];							inform_L[102][5] = l_cell_wire[77];							inform_L[71][5] = l_cell_wire[78];							inform_L[103][5] = l_cell_wire[79];							inform_L[72][5] = l_cell_wire[80];							inform_L[104][5] = l_cell_wire[81];							inform_L[73][5] = l_cell_wire[82];							inform_L[105][5] = l_cell_wire[83];							inform_L[74][5] = l_cell_wire[84];							inform_L[106][5] = l_cell_wire[85];							inform_L[75][5] = l_cell_wire[86];							inform_L[107][5] = l_cell_wire[87];							inform_L[76][5] = l_cell_wire[88];							inform_L[108][5] = l_cell_wire[89];							inform_L[77][5] = l_cell_wire[90];							inform_L[109][5] = l_cell_wire[91];							inform_L[78][5] = l_cell_wire[92];							inform_L[110][5] = l_cell_wire[93];							inform_L[79][5] = l_cell_wire[94];							inform_L[111][5] = l_cell_wire[95];							inform_L[80][5] = l_cell_wire[96];							inform_L[112][5] = l_cell_wire[97];							inform_L[81][5] = l_cell_wire[98];							inform_L[113][5] = l_cell_wire[99];							inform_L[82][5] = l_cell_wire[100];							inform_L[114][5] = l_cell_wire[101];							inform_L[83][5] = l_cell_wire[102];							inform_L[115][5] = l_cell_wire[103];							inform_L[84][5] = l_cell_wire[104];							inform_L[116][5] = l_cell_wire[105];							inform_L[85][5] = l_cell_wire[106];							inform_L[117][5] = l_cell_wire[107];							inform_L[86][5] = l_cell_wire[108];							inform_L[118][5] = l_cell_wire[109];							inform_L[87][5] = l_cell_wire[110];							inform_L[119][5] = l_cell_wire[111];							inform_L[88][5] = l_cell_wire[112];							inform_L[120][5] = l_cell_wire[113];							inform_L[89][5] = l_cell_wire[114];							inform_L[121][5] = l_cell_wire[115];							inform_L[90][5] = l_cell_wire[116];							inform_L[122][5] = l_cell_wire[117];							inform_L[91][5] = l_cell_wire[118];							inform_L[123][5] = l_cell_wire[119];							inform_L[92][5] = l_cell_wire[120];							inform_L[124][5] = l_cell_wire[121];							inform_L[93][5] = l_cell_wire[122];							inform_L[125][5] = l_cell_wire[123];							inform_L[94][5] = l_cell_wire[124];							inform_L[126][5] = l_cell_wire[125];							inform_L[95][5] = l_cell_wire[126];							inform_L[127][5] = l_cell_wire[127];							inform_L[128][5] = l_cell_wire[128];							inform_L[160][5] = l_cell_wire[129];							inform_L[129][5] = l_cell_wire[130];							inform_L[161][5] = l_cell_wire[131];							inform_L[130][5] = l_cell_wire[132];							inform_L[162][5] = l_cell_wire[133];							inform_L[131][5] = l_cell_wire[134];							inform_L[163][5] = l_cell_wire[135];							inform_L[132][5] = l_cell_wire[136];							inform_L[164][5] = l_cell_wire[137];							inform_L[133][5] = l_cell_wire[138];							inform_L[165][5] = l_cell_wire[139];							inform_L[134][5] = l_cell_wire[140];							inform_L[166][5] = l_cell_wire[141];							inform_L[135][5] = l_cell_wire[142];							inform_L[167][5] = l_cell_wire[143];							inform_L[136][5] = l_cell_wire[144];							inform_L[168][5] = l_cell_wire[145];							inform_L[137][5] = l_cell_wire[146];							inform_L[169][5] = l_cell_wire[147];							inform_L[138][5] = l_cell_wire[148];							inform_L[170][5] = l_cell_wire[149];							inform_L[139][5] = l_cell_wire[150];							inform_L[171][5] = l_cell_wire[151];							inform_L[140][5] = l_cell_wire[152];							inform_L[172][5] = l_cell_wire[153];							inform_L[141][5] = l_cell_wire[154];							inform_L[173][5] = l_cell_wire[155];							inform_L[142][5] = l_cell_wire[156];							inform_L[174][5] = l_cell_wire[157];							inform_L[143][5] = l_cell_wire[158];							inform_L[175][5] = l_cell_wire[159];							inform_L[144][5] = l_cell_wire[160];							inform_L[176][5] = l_cell_wire[161];							inform_L[145][5] = l_cell_wire[162];							inform_L[177][5] = l_cell_wire[163];							inform_L[146][5] = l_cell_wire[164];							inform_L[178][5] = l_cell_wire[165];							inform_L[147][5] = l_cell_wire[166];							inform_L[179][5] = l_cell_wire[167];							inform_L[148][5] = l_cell_wire[168];							inform_L[180][5] = l_cell_wire[169];							inform_L[149][5] = l_cell_wire[170];							inform_L[181][5] = l_cell_wire[171];							inform_L[150][5] = l_cell_wire[172];							inform_L[182][5] = l_cell_wire[173];							inform_L[151][5] = l_cell_wire[174];							inform_L[183][5] = l_cell_wire[175];							inform_L[152][5] = l_cell_wire[176];							inform_L[184][5] = l_cell_wire[177];							inform_L[153][5] = l_cell_wire[178];							inform_L[185][5] = l_cell_wire[179];							inform_L[154][5] = l_cell_wire[180];							inform_L[186][5] = l_cell_wire[181];							inform_L[155][5] = l_cell_wire[182];							inform_L[187][5] = l_cell_wire[183];							inform_L[156][5] = l_cell_wire[184];							inform_L[188][5] = l_cell_wire[185];							inform_L[157][5] = l_cell_wire[186];							inform_L[189][5] = l_cell_wire[187];							inform_L[158][5] = l_cell_wire[188];							inform_L[190][5] = l_cell_wire[189];							inform_L[159][5] = l_cell_wire[190];							inform_L[191][5] = l_cell_wire[191];							inform_L[192][5] = l_cell_wire[192];							inform_L[224][5] = l_cell_wire[193];							inform_L[193][5] = l_cell_wire[194];							inform_L[225][5] = l_cell_wire[195];							inform_L[194][5] = l_cell_wire[196];							inform_L[226][5] = l_cell_wire[197];							inform_L[195][5] = l_cell_wire[198];							inform_L[227][5] = l_cell_wire[199];							inform_L[196][5] = l_cell_wire[200];							inform_L[228][5] = l_cell_wire[201];							inform_L[197][5] = l_cell_wire[202];							inform_L[229][5] = l_cell_wire[203];							inform_L[198][5] = l_cell_wire[204];							inform_L[230][5] = l_cell_wire[205];							inform_L[199][5] = l_cell_wire[206];							inform_L[231][5] = l_cell_wire[207];							inform_L[200][5] = l_cell_wire[208];							inform_L[232][5] = l_cell_wire[209];							inform_L[201][5] = l_cell_wire[210];							inform_L[233][5] = l_cell_wire[211];							inform_L[202][5] = l_cell_wire[212];							inform_L[234][5] = l_cell_wire[213];							inform_L[203][5] = l_cell_wire[214];							inform_L[235][5] = l_cell_wire[215];							inform_L[204][5] = l_cell_wire[216];							inform_L[236][5] = l_cell_wire[217];							inform_L[205][5] = l_cell_wire[218];							inform_L[237][5] = l_cell_wire[219];							inform_L[206][5] = l_cell_wire[220];							inform_L[238][5] = l_cell_wire[221];							inform_L[207][5] = l_cell_wire[222];							inform_L[239][5] = l_cell_wire[223];							inform_L[208][5] = l_cell_wire[224];							inform_L[240][5] = l_cell_wire[225];							inform_L[209][5] = l_cell_wire[226];							inform_L[241][5] = l_cell_wire[227];							inform_L[210][5] = l_cell_wire[228];							inform_L[242][5] = l_cell_wire[229];							inform_L[211][5] = l_cell_wire[230];							inform_L[243][5] = l_cell_wire[231];							inform_L[212][5] = l_cell_wire[232];							inform_L[244][5] = l_cell_wire[233];							inform_L[213][5] = l_cell_wire[234];							inform_L[245][5] = l_cell_wire[235];							inform_L[214][5] = l_cell_wire[236];							inform_L[246][5] = l_cell_wire[237];							inform_L[215][5] = l_cell_wire[238];							inform_L[247][5] = l_cell_wire[239];							inform_L[216][5] = l_cell_wire[240];							inform_L[248][5] = l_cell_wire[241];							inform_L[217][5] = l_cell_wire[242];							inform_L[249][5] = l_cell_wire[243];							inform_L[218][5] = l_cell_wire[244];							inform_L[250][5] = l_cell_wire[245];							inform_L[219][5] = l_cell_wire[246];							inform_L[251][5] = l_cell_wire[247];							inform_L[220][5] = l_cell_wire[248];							inform_L[252][5] = l_cell_wire[249];							inform_L[221][5] = l_cell_wire[250];							inform_L[253][5] = l_cell_wire[251];							inform_L[222][5] = l_cell_wire[252];							inform_L[254][5] = l_cell_wire[253];							inform_L[223][5] = l_cell_wire[254];							inform_L[255][5] = l_cell_wire[255];							inform_L[256][5] = l_cell_wire[256];							inform_L[288][5] = l_cell_wire[257];							inform_L[257][5] = l_cell_wire[258];							inform_L[289][5] = l_cell_wire[259];							inform_L[258][5] = l_cell_wire[260];							inform_L[290][5] = l_cell_wire[261];							inform_L[259][5] = l_cell_wire[262];							inform_L[291][5] = l_cell_wire[263];							inform_L[260][5] = l_cell_wire[264];							inform_L[292][5] = l_cell_wire[265];							inform_L[261][5] = l_cell_wire[266];							inform_L[293][5] = l_cell_wire[267];							inform_L[262][5] = l_cell_wire[268];							inform_L[294][5] = l_cell_wire[269];							inform_L[263][5] = l_cell_wire[270];							inform_L[295][5] = l_cell_wire[271];							inform_L[264][5] = l_cell_wire[272];							inform_L[296][5] = l_cell_wire[273];							inform_L[265][5] = l_cell_wire[274];							inform_L[297][5] = l_cell_wire[275];							inform_L[266][5] = l_cell_wire[276];							inform_L[298][5] = l_cell_wire[277];							inform_L[267][5] = l_cell_wire[278];							inform_L[299][5] = l_cell_wire[279];							inform_L[268][5] = l_cell_wire[280];							inform_L[300][5] = l_cell_wire[281];							inform_L[269][5] = l_cell_wire[282];							inform_L[301][5] = l_cell_wire[283];							inform_L[270][5] = l_cell_wire[284];							inform_L[302][5] = l_cell_wire[285];							inform_L[271][5] = l_cell_wire[286];							inform_L[303][5] = l_cell_wire[287];							inform_L[272][5] = l_cell_wire[288];							inform_L[304][5] = l_cell_wire[289];							inform_L[273][5] = l_cell_wire[290];							inform_L[305][5] = l_cell_wire[291];							inform_L[274][5] = l_cell_wire[292];							inform_L[306][5] = l_cell_wire[293];							inform_L[275][5] = l_cell_wire[294];							inform_L[307][5] = l_cell_wire[295];							inform_L[276][5] = l_cell_wire[296];							inform_L[308][5] = l_cell_wire[297];							inform_L[277][5] = l_cell_wire[298];							inform_L[309][5] = l_cell_wire[299];							inform_L[278][5] = l_cell_wire[300];							inform_L[310][5] = l_cell_wire[301];							inform_L[279][5] = l_cell_wire[302];							inform_L[311][5] = l_cell_wire[303];							inform_L[280][5] = l_cell_wire[304];							inform_L[312][5] = l_cell_wire[305];							inform_L[281][5] = l_cell_wire[306];							inform_L[313][5] = l_cell_wire[307];							inform_L[282][5] = l_cell_wire[308];							inform_L[314][5] = l_cell_wire[309];							inform_L[283][5] = l_cell_wire[310];							inform_L[315][5] = l_cell_wire[311];							inform_L[284][5] = l_cell_wire[312];							inform_L[316][5] = l_cell_wire[313];							inform_L[285][5] = l_cell_wire[314];							inform_L[317][5] = l_cell_wire[315];							inform_L[286][5] = l_cell_wire[316];							inform_L[318][5] = l_cell_wire[317];							inform_L[287][5] = l_cell_wire[318];							inform_L[319][5] = l_cell_wire[319];							inform_L[320][5] = l_cell_wire[320];							inform_L[352][5] = l_cell_wire[321];							inform_L[321][5] = l_cell_wire[322];							inform_L[353][5] = l_cell_wire[323];							inform_L[322][5] = l_cell_wire[324];							inform_L[354][5] = l_cell_wire[325];							inform_L[323][5] = l_cell_wire[326];							inform_L[355][5] = l_cell_wire[327];							inform_L[324][5] = l_cell_wire[328];							inform_L[356][5] = l_cell_wire[329];							inform_L[325][5] = l_cell_wire[330];							inform_L[357][5] = l_cell_wire[331];							inform_L[326][5] = l_cell_wire[332];							inform_L[358][5] = l_cell_wire[333];							inform_L[327][5] = l_cell_wire[334];							inform_L[359][5] = l_cell_wire[335];							inform_L[328][5] = l_cell_wire[336];							inform_L[360][5] = l_cell_wire[337];							inform_L[329][5] = l_cell_wire[338];							inform_L[361][5] = l_cell_wire[339];							inform_L[330][5] = l_cell_wire[340];							inform_L[362][5] = l_cell_wire[341];							inform_L[331][5] = l_cell_wire[342];							inform_L[363][5] = l_cell_wire[343];							inform_L[332][5] = l_cell_wire[344];							inform_L[364][5] = l_cell_wire[345];							inform_L[333][5] = l_cell_wire[346];							inform_L[365][5] = l_cell_wire[347];							inform_L[334][5] = l_cell_wire[348];							inform_L[366][5] = l_cell_wire[349];							inform_L[335][5] = l_cell_wire[350];							inform_L[367][5] = l_cell_wire[351];							inform_L[336][5] = l_cell_wire[352];							inform_L[368][5] = l_cell_wire[353];							inform_L[337][5] = l_cell_wire[354];							inform_L[369][5] = l_cell_wire[355];							inform_L[338][5] = l_cell_wire[356];							inform_L[370][5] = l_cell_wire[357];							inform_L[339][5] = l_cell_wire[358];							inform_L[371][5] = l_cell_wire[359];							inform_L[340][5] = l_cell_wire[360];							inform_L[372][5] = l_cell_wire[361];							inform_L[341][5] = l_cell_wire[362];							inform_L[373][5] = l_cell_wire[363];							inform_L[342][5] = l_cell_wire[364];							inform_L[374][5] = l_cell_wire[365];							inform_L[343][5] = l_cell_wire[366];							inform_L[375][5] = l_cell_wire[367];							inform_L[344][5] = l_cell_wire[368];							inform_L[376][5] = l_cell_wire[369];							inform_L[345][5] = l_cell_wire[370];							inform_L[377][5] = l_cell_wire[371];							inform_L[346][5] = l_cell_wire[372];							inform_L[378][5] = l_cell_wire[373];							inform_L[347][5] = l_cell_wire[374];							inform_L[379][5] = l_cell_wire[375];							inform_L[348][5] = l_cell_wire[376];							inform_L[380][5] = l_cell_wire[377];							inform_L[349][5] = l_cell_wire[378];							inform_L[381][5] = l_cell_wire[379];							inform_L[350][5] = l_cell_wire[380];							inform_L[382][5] = l_cell_wire[381];							inform_L[351][5] = l_cell_wire[382];							inform_L[383][5] = l_cell_wire[383];							inform_L[384][5] = l_cell_wire[384];							inform_L[416][5] = l_cell_wire[385];							inform_L[385][5] = l_cell_wire[386];							inform_L[417][5] = l_cell_wire[387];							inform_L[386][5] = l_cell_wire[388];							inform_L[418][5] = l_cell_wire[389];							inform_L[387][5] = l_cell_wire[390];							inform_L[419][5] = l_cell_wire[391];							inform_L[388][5] = l_cell_wire[392];							inform_L[420][5] = l_cell_wire[393];							inform_L[389][5] = l_cell_wire[394];							inform_L[421][5] = l_cell_wire[395];							inform_L[390][5] = l_cell_wire[396];							inform_L[422][5] = l_cell_wire[397];							inform_L[391][5] = l_cell_wire[398];							inform_L[423][5] = l_cell_wire[399];							inform_L[392][5] = l_cell_wire[400];							inform_L[424][5] = l_cell_wire[401];							inform_L[393][5] = l_cell_wire[402];							inform_L[425][5] = l_cell_wire[403];							inform_L[394][5] = l_cell_wire[404];							inform_L[426][5] = l_cell_wire[405];							inform_L[395][5] = l_cell_wire[406];							inform_L[427][5] = l_cell_wire[407];							inform_L[396][5] = l_cell_wire[408];							inform_L[428][5] = l_cell_wire[409];							inform_L[397][5] = l_cell_wire[410];							inform_L[429][5] = l_cell_wire[411];							inform_L[398][5] = l_cell_wire[412];							inform_L[430][5] = l_cell_wire[413];							inform_L[399][5] = l_cell_wire[414];							inform_L[431][5] = l_cell_wire[415];							inform_L[400][5] = l_cell_wire[416];							inform_L[432][5] = l_cell_wire[417];							inform_L[401][5] = l_cell_wire[418];							inform_L[433][5] = l_cell_wire[419];							inform_L[402][5] = l_cell_wire[420];							inform_L[434][5] = l_cell_wire[421];							inform_L[403][5] = l_cell_wire[422];							inform_L[435][5] = l_cell_wire[423];							inform_L[404][5] = l_cell_wire[424];							inform_L[436][5] = l_cell_wire[425];							inform_L[405][5] = l_cell_wire[426];							inform_L[437][5] = l_cell_wire[427];							inform_L[406][5] = l_cell_wire[428];							inform_L[438][5] = l_cell_wire[429];							inform_L[407][5] = l_cell_wire[430];							inform_L[439][5] = l_cell_wire[431];							inform_L[408][5] = l_cell_wire[432];							inform_L[440][5] = l_cell_wire[433];							inform_L[409][5] = l_cell_wire[434];							inform_L[441][5] = l_cell_wire[435];							inform_L[410][5] = l_cell_wire[436];							inform_L[442][5] = l_cell_wire[437];							inform_L[411][5] = l_cell_wire[438];							inform_L[443][5] = l_cell_wire[439];							inform_L[412][5] = l_cell_wire[440];							inform_L[444][5] = l_cell_wire[441];							inform_L[413][5] = l_cell_wire[442];							inform_L[445][5] = l_cell_wire[443];							inform_L[414][5] = l_cell_wire[444];							inform_L[446][5] = l_cell_wire[445];							inform_L[415][5] = l_cell_wire[446];							inform_L[447][5] = l_cell_wire[447];							inform_L[448][5] = l_cell_wire[448];							inform_L[480][5] = l_cell_wire[449];							inform_L[449][5] = l_cell_wire[450];							inform_L[481][5] = l_cell_wire[451];							inform_L[450][5] = l_cell_wire[452];							inform_L[482][5] = l_cell_wire[453];							inform_L[451][5] = l_cell_wire[454];							inform_L[483][5] = l_cell_wire[455];							inform_L[452][5] = l_cell_wire[456];							inform_L[484][5] = l_cell_wire[457];							inform_L[453][5] = l_cell_wire[458];							inform_L[485][5] = l_cell_wire[459];							inform_L[454][5] = l_cell_wire[460];							inform_L[486][5] = l_cell_wire[461];							inform_L[455][5] = l_cell_wire[462];							inform_L[487][5] = l_cell_wire[463];							inform_L[456][5] = l_cell_wire[464];							inform_L[488][5] = l_cell_wire[465];							inform_L[457][5] = l_cell_wire[466];							inform_L[489][5] = l_cell_wire[467];							inform_L[458][5] = l_cell_wire[468];							inform_L[490][5] = l_cell_wire[469];							inform_L[459][5] = l_cell_wire[470];							inform_L[491][5] = l_cell_wire[471];							inform_L[460][5] = l_cell_wire[472];							inform_L[492][5] = l_cell_wire[473];							inform_L[461][5] = l_cell_wire[474];							inform_L[493][5] = l_cell_wire[475];							inform_L[462][5] = l_cell_wire[476];							inform_L[494][5] = l_cell_wire[477];							inform_L[463][5] = l_cell_wire[478];							inform_L[495][5] = l_cell_wire[479];							inform_L[464][5] = l_cell_wire[480];							inform_L[496][5] = l_cell_wire[481];							inform_L[465][5] = l_cell_wire[482];							inform_L[497][5] = l_cell_wire[483];							inform_L[466][5] = l_cell_wire[484];							inform_L[498][5] = l_cell_wire[485];							inform_L[467][5] = l_cell_wire[486];							inform_L[499][5] = l_cell_wire[487];							inform_L[468][5] = l_cell_wire[488];							inform_L[500][5] = l_cell_wire[489];							inform_L[469][5] = l_cell_wire[490];							inform_L[501][5] = l_cell_wire[491];							inform_L[470][5] = l_cell_wire[492];							inform_L[502][5] = l_cell_wire[493];							inform_L[471][5] = l_cell_wire[494];							inform_L[503][5] = l_cell_wire[495];							inform_L[472][5] = l_cell_wire[496];							inform_L[504][5] = l_cell_wire[497];							inform_L[473][5] = l_cell_wire[498];							inform_L[505][5] = l_cell_wire[499];							inform_L[474][5] = l_cell_wire[500];							inform_L[506][5] = l_cell_wire[501];							inform_L[475][5] = l_cell_wire[502];							inform_L[507][5] = l_cell_wire[503];							inform_L[476][5] = l_cell_wire[504];							inform_L[508][5] = l_cell_wire[505];							inform_L[477][5] = l_cell_wire[506];							inform_L[509][5] = l_cell_wire[507];							inform_L[478][5] = l_cell_wire[508];							inform_L[510][5] = l_cell_wire[509];							inform_L[479][5] = l_cell_wire[510];							inform_L[511][5] = l_cell_wire[511];							inform_L[512][5] = l_cell_wire[512];							inform_L[544][5] = l_cell_wire[513];							inform_L[513][5] = l_cell_wire[514];							inform_L[545][5] = l_cell_wire[515];							inform_L[514][5] = l_cell_wire[516];							inform_L[546][5] = l_cell_wire[517];							inform_L[515][5] = l_cell_wire[518];							inform_L[547][5] = l_cell_wire[519];							inform_L[516][5] = l_cell_wire[520];							inform_L[548][5] = l_cell_wire[521];							inform_L[517][5] = l_cell_wire[522];							inform_L[549][5] = l_cell_wire[523];							inform_L[518][5] = l_cell_wire[524];							inform_L[550][5] = l_cell_wire[525];							inform_L[519][5] = l_cell_wire[526];							inform_L[551][5] = l_cell_wire[527];							inform_L[520][5] = l_cell_wire[528];							inform_L[552][5] = l_cell_wire[529];							inform_L[521][5] = l_cell_wire[530];							inform_L[553][5] = l_cell_wire[531];							inform_L[522][5] = l_cell_wire[532];							inform_L[554][5] = l_cell_wire[533];							inform_L[523][5] = l_cell_wire[534];							inform_L[555][5] = l_cell_wire[535];							inform_L[524][5] = l_cell_wire[536];							inform_L[556][5] = l_cell_wire[537];							inform_L[525][5] = l_cell_wire[538];							inform_L[557][5] = l_cell_wire[539];							inform_L[526][5] = l_cell_wire[540];							inform_L[558][5] = l_cell_wire[541];							inform_L[527][5] = l_cell_wire[542];							inform_L[559][5] = l_cell_wire[543];							inform_L[528][5] = l_cell_wire[544];							inform_L[560][5] = l_cell_wire[545];							inform_L[529][5] = l_cell_wire[546];							inform_L[561][5] = l_cell_wire[547];							inform_L[530][5] = l_cell_wire[548];							inform_L[562][5] = l_cell_wire[549];							inform_L[531][5] = l_cell_wire[550];							inform_L[563][5] = l_cell_wire[551];							inform_L[532][5] = l_cell_wire[552];							inform_L[564][5] = l_cell_wire[553];							inform_L[533][5] = l_cell_wire[554];							inform_L[565][5] = l_cell_wire[555];							inform_L[534][5] = l_cell_wire[556];							inform_L[566][5] = l_cell_wire[557];							inform_L[535][5] = l_cell_wire[558];							inform_L[567][5] = l_cell_wire[559];							inform_L[536][5] = l_cell_wire[560];							inform_L[568][5] = l_cell_wire[561];							inform_L[537][5] = l_cell_wire[562];							inform_L[569][5] = l_cell_wire[563];							inform_L[538][5] = l_cell_wire[564];							inform_L[570][5] = l_cell_wire[565];							inform_L[539][5] = l_cell_wire[566];							inform_L[571][5] = l_cell_wire[567];							inform_L[540][5] = l_cell_wire[568];							inform_L[572][5] = l_cell_wire[569];							inform_L[541][5] = l_cell_wire[570];							inform_L[573][5] = l_cell_wire[571];							inform_L[542][5] = l_cell_wire[572];							inform_L[574][5] = l_cell_wire[573];							inform_L[543][5] = l_cell_wire[574];							inform_L[575][5] = l_cell_wire[575];							inform_L[576][5] = l_cell_wire[576];							inform_L[608][5] = l_cell_wire[577];							inform_L[577][5] = l_cell_wire[578];							inform_L[609][5] = l_cell_wire[579];							inform_L[578][5] = l_cell_wire[580];							inform_L[610][5] = l_cell_wire[581];							inform_L[579][5] = l_cell_wire[582];							inform_L[611][5] = l_cell_wire[583];							inform_L[580][5] = l_cell_wire[584];							inform_L[612][5] = l_cell_wire[585];							inform_L[581][5] = l_cell_wire[586];							inform_L[613][5] = l_cell_wire[587];							inform_L[582][5] = l_cell_wire[588];							inform_L[614][5] = l_cell_wire[589];							inform_L[583][5] = l_cell_wire[590];							inform_L[615][5] = l_cell_wire[591];							inform_L[584][5] = l_cell_wire[592];							inform_L[616][5] = l_cell_wire[593];							inform_L[585][5] = l_cell_wire[594];							inform_L[617][5] = l_cell_wire[595];							inform_L[586][5] = l_cell_wire[596];							inform_L[618][5] = l_cell_wire[597];							inform_L[587][5] = l_cell_wire[598];							inform_L[619][5] = l_cell_wire[599];							inform_L[588][5] = l_cell_wire[600];							inform_L[620][5] = l_cell_wire[601];							inform_L[589][5] = l_cell_wire[602];							inform_L[621][5] = l_cell_wire[603];							inform_L[590][5] = l_cell_wire[604];							inform_L[622][5] = l_cell_wire[605];							inform_L[591][5] = l_cell_wire[606];							inform_L[623][5] = l_cell_wire[607];							inform_L[592][5] = l_cell_wire[608];							inform_L[624][5] = l_cell_wire[609];							inform_L[593][5] = l_cell_wire[610];							inform_L[625][5] = l_cell_wire[611];							inform_L[594][5] = l_cell_wire[612];							inform_L[626][5] = l_cell_wire[613];							inform_L[595][5] = l_cell_wire[614];							inform_L[627][5] = l_cell_wire[615];							inform_L[596][5] = l_cell_wire[616];							inform_L[628][5] = l_cell_wire[617];							inform_L[597][5] = l_cell_wire[618];							inform_L[629][5] = l_cell_wire[619];							inform_L[598][5] = l_cell_wire[620];							inform_L[630][5] = l_cell_wire[621];							inform_L[599][5] = l_cell_wire[622];							inform_L[631][5] = l_cell_wire[623];							inform_L[600][5] = l_cell_wire[624];							inform_L[632][5] = l_cell_wire[625];							inform_L[601][5] = l_cell_wire[626];							inform_L[633][5] = l_cell_wire[627];							inform_L[602][5] = l_cell_wire[628];							inform_L[634][5] = l_cell_wire[629];							inform_L[603][5] = l_cell_wire[630];							inform_L[635][5] = l_cell_wire[631];							inform_L[604][5] = l_cell_wire[632];							inform_L[636][5] = l_cell_wire[633];							inform_L[605][5] = l_cell_wire[634];							inform_L[637][5] = l_cell_wire[635];							inform_L[606][5] = l_cell_wire[636];							inform_L[638][5] = l_cell_wire[637];							inform_L[607][5] = l_cell_wire[638];							inform_L[639][5] = l_cell_wire[639];							inform_L[640][5] = l_cell_wire[640];							inform_L[672][5] = l_cell_wire[641];							inform_L[641][5] = l_cell_wire[642];							inform_L[673][5] = l_cell_wire[643];							inform_L[642][5] = l_cell_wire[644];							inform_L[674][5] = l_cell_wire[645];							inform_L[643][5] = l_cell_wire[646];							inform_L[675][5] = l_cell_wire[647];							inform_L[644][5] = l_cell_wire[648];							inform_L[676][5] = l_cell_wire[649];							inform_L[645][5] = l_cell_wire[650];							inform_L[677][5] = l_cell_wire[651];							inform_L[646][5] = l_cell_wire[652];							inform_L[678][5] = l_cell_wire[653];							inform_L[647][5] = l_cell_wire[654];							inform_L[679][5] = l_cell_wire[655];							inform_L[648][5] = l_cell_wire[656];							inform_L[680][5] = l_cell_wire[657];							inform_L[649][5] = l_cell_wire[658];							inform_L[681][5] = l_cell_wire[659];							inform_L[650][5] = l_cell_wire[660];							inform_L[682][5] = l_cell_wire[661];							inform_L[651][5] = l_cell_wire[662];							inform_L[683][5] = l_cell_wire[663];							inform_L[652][5] = l_cell_wire[664];							inform_L[684][5] = l_cell_wire[665];							inform_L[653][5] = l_cell_wire[666];							inform_L[685][5] = l_cell_wire[667];							inform_L[654][5] = l_cell_wire[668];							inform_L[686][5] = l_cell_wire[669];							inform_L[655][5] = l_cell_wire[670];							inform_L[687][5] = l_cell_wire[671];							inform_L[656][5] = l_cell_wire[672];							inform_L[688][5] = l_cell_wire[673];							inform_L[657][5] = l_cell_wire[674];							inform_L[689][5] = l_cell_wire[675];							inform_L[658][5] = l_cell_wire[676];							inform_L[690][5] = l_cell_wire[677];							inform_L[659][5] = l_cell_wire[678];							inform_L[691][5] = l_cell_wire[679];							inform_L[660][5] = l_cell_wire[680];							inform_L[692][5] = l_cell_wire[681];							inform_L[661][5] = l_cell_wire[682];							inform_L[693][5] = l_cell_wire[683];							inform_L[662][5] = l_cell_wire[684];							inform_L[694][5] = l_cell_wire[685];							inform_L[663][5] = l_cell_wire[686];							inform_L[695][5] = l_cell_wire[687];							inform_L[664][5] = l_cell_wire[688];							inform_L[696][5] = l_cell_wire[689];							inform_L[665][5] = l_cell_wire[690];							inform_L[697][5] = l_cell_wire[691];							inform_L[666][5] = l_cell_wire[692];							inform_L[698][5] = l_cell_wire[693];							inform_L[667][5] = l_cell_wire[694];							inform_L[699][5] = l_cell_wire[695];							inform_L[668][5] = l_cell_wire[696];							inform_L[700][5] = l_cell_wire[697];							inform_L[669][5] = l_cell_wire[698];							inform_L[701][5] = l_cell_wire[699];							inform_L[670][5] = l_cell_wire[700];							inform_L[702][5] = l_cell_wire[701];							inform_L[671][5] = l_cell_wire[702];							inform_L[703][5] = l_cell_wire[703];							inform_L[704][5] = l_cell_wire[704];							inform_L[736][5] = l_cell_wire[705];							inform_L[705][5] = l_cell_wire[706];							inform_L[737][5] = l_cell_wire[707];							inform_L[706][5] = l_cell_wire[708];							inform_L[738][5] = l_cell_wire[709];							inform_L[707][5] = l_cell_wire[710];							inform_L[739][5] = l_cell_wire[711];							inform_L[708][5] = l_cell_wire[712];							inform_L[740][5] = l_cell_wire[713];							inform_L[709][5] = l_cell_wire[714];							inform_L[741][5] = l_cell_wire[715];							inform_L[710][5] = l_cell_wire[716];							inform_L[742][5] = l_cell_wire[717];							inform_L[711][5] = l_cell_wire[718];							inform_L[743][5] = l_cell_wire[719];							inform_L[712][5] = l_cell_wire[720];							inform_L[744][5] = l_cell_wire[721];							inform_L[713][5] = l_cell_wire[722];							inform_L[745][5] = l_cell_wire[723];							inform_L[714][5] = l_cell_wire[724];							inform_L[746][5] = l_cell_wire[725];							inform_L[715][5] = l_cell_wire[726];							inform_L[747][5] = l_cell_wire[727];							inform_L[716][5] = l_cell_wire[728];							inform_L[748][5] = l_cell_wire[729];							inform_L[717][5] = l_cell_wire[730];							inform_L[749][5] = l_cell_wire[731];							inform_L[718][5] = l_cell_wire[732];							inform_L[750][5] = l_cell_wire[733];							inform_L[719][5] = l_cell_wire[734];							inform_L[751][5] = l_cell_wire[735];							inform_L[720][5] = l_cell_wire[736];							inform_L[752][5] = l_cell_wire[737];							inform_L[721][5] = l_cell_wire[738];							inform_L[753][5] = l_cell_wire[739];							inform_L[722][5] = l_cell_wire[740];							inform_L[754][5] = l_cell_wire[741];							inform_L[723][5] = l_cell_wire[742];							inform_L[755][5] = l_cell_wire[743];							inform_L[724][5] = l_cell_wire[744];							inform_L[756][5] = l_cell_wire[745];							inform_L[725][5] = l_cell_wire[746];							inform_L[757][5] = l_cell_wire[747];							inform_L[726][5] = l_cell_wire[748];							inform_L[758][5] = l_cell_wire[749];							inform_L[727][5] = l_cell_wire[750];							inform_L[759][5] = l_cell_wire[751];							inform_L[728][5] = l_cell_wire[752];							inform_L[760][5] = l_cell_wire[753];							inform_L[729][5] = l_cell_wire[754];							inform_L[761][5] = l_cell_wire[755];							inform_L[730][5] = l_cell_wire[756];							inform_L[762][5] = l_cell_wire[757];							inform_L[731][5] = l_cell_wire[758];							inform_L[763][5] = l_cell_wire[759];							inform_L[732][5] = l_cell_wire[760];							inform_L[764][5] = l_cell_wire[761];							inform_L[733][5] = l_cell_wire[762];							inform_L[765][5] = l_cell_wire[763];							inform_L[734][5] = l_cell_wire[764];							inform_L[766][5] = l_cell_wire[765];							inform_L[735][5] = l_cell_wire[766];							inform_L[767][5] = l_cell_wire[767];							inform_L[768][5] = l_cell_wire[768];							inform_L[800][5] = l_cell_wire[769];							inform_L[769][5] = l_cell_wire[770];							inform_L[801][5] = l_cell_wire[771];							inform_L[770][5] = l_cell_wire[772];							inform_L[802][5] = l_cell_wire[773];							inform_L[771][5] = l_cell_wire[774];							inform_L[803][5] = l_cell_wire[775];							inform_L[772][5] = l_cell_wire[776];							inform_L[804][5] = l_cell_wire[777];							inform_L[773][5] = l_cell_wire[778];							inform_L[805][5] = l_cell_wire[779];							inform_L[774][5] = l_cell_wire[780];							inform_L[806][5] = l_cell_wire[781];							inform_L[775][5] = l_cell_wire[782];							inform_L[807][5] = l_cell_wire[783];							inform_L[776][5] = l_cell_wire[784];							inform_L[808][5] = l_cell_wire[785];							inform_L[777][5] = l_cell_wire[786];							inform_L[809][5] = l_cell_wire[787];							inform_L[778][5] = l_cell_wire[788];							inform_L[810][5] = l_cell_wire[789];							inform_L[779][5] = l_cell_wire[790];							inform_L[811][5] = l_cell_wire[791];							inform_L[780][5] = l_cell_wire[792];							inform_L[812][5] = l_cell_wire[793];							inform_L[781][5] = l_cell_wire[794];							inform_L[813][5] = l_cell_wire[795];							inform_L[782][5] = l_cell_wire[796];							inform_L[814][5] = l_cell_wire[797];							inform_L[783][5] = l_cell_wire[798];							inform_L[815][5] = l_cell_wire[799];							inform_L[784][5] = l_cell_wire[800];							inform_L[816][5] = l_cell_wire[801];							inform_L[785][5] = l_cell_wire[802];							inform_L[817][5] = l_cell_wire[803];							inform_L[786][5] = l_cell_wire[804];							inform_L[818][5] = l_cell_wire[805];							inform_L[787][5] = l_cell_wire[806];							inform_L[819][5] = l_cell_wire[807];							inform_L[788][5] = l_cell_wire[808];							inform_L[820][5] = l_cell_wire[809];							inform_L[789][5] = l_cell_wire[810];							inform_L[821][5] = l_cell_wire[811];							inform_L[790][5] = l_cell_wire[812];							inform_L[822][5] = l_cell_wire[813];							inform_L[791][5] = l_cell_wire[814];							inform_L[823][5] = l_cell_wire[815];							inform_L[792][5] = l_cell_wire[816];							inform_L[824][5] = l_cell_wire[817];							inform_L[793][5] = l_cell_wire[818];							inform_L[825][5] = l_cell_wire[819];							inform_L[794][5] = l_cell_wire[820];							inform_L[826][5] = l_cell_wire[821];							inform_L[795][5] = l_cell_wire[822];							inform_L[827][5] = l_cell_wire[823];							inform_L[796][5] = l_cell_wire[824];							inform_L[828][5] = l_cell_wire[825];							inform_L[797][5] = l_cell_wire[826];							inform_L[829][5] = l_cell_wire[827];							inform_L[798][5] = l_cell_wire[828];							inform_L[830][5] = l_cell_wire[829];							inform_L[799][5] = l_cell_wire[830];							inform_L[831][5] = l_cell_wire[831];							inform_L[832][5] = l_cell_wire[832];							inform_L[864][5] = l_cell_wire[833];							inform_L[833][5] = l_cell_wire[834];							inform_L[865][5] = l_cell_wire[835];							inform_L[834][5] = l_cell_wire[836];							inform_L[866][5] = l_cell_wire[837];							inform_L[835][5] = l_cell_wire[838];							inform_L[867][5] = l_cell_wire[839];							inform_L[836][5] = l_cell_wire[840];							inform_L[868][5] = l_cell_wire[841];							inform_L[837][5] = l_cell_wire[842];							inform_L[869][5] = l_cell_wire[843];							inform_L[838][5] = l_cell_wire[844];							inform_L[870][5] = l_cell_wire[845];							inform_L[839][5] = l_cell_wire[846];							inform_L[871][5] = l_cell_wire[847];							inform_L[840][5] = l_cell_wire[848];							inform_L[872][5] = l_cell_wire[849];							inform_L[841][5] = l_cell_wire[850];							inform_L[873][5] = l_cell_wire[851];							inform_L[842][5] = l_cell_wire[852];							inform_L[874][5] = l_cell_wire[853];							inform_L[843][5] = l_cell_wire[854];							inform_L[875][5] = l_cell_wire[855];							inform_L[844][5] = l_cell_wire[856];							inform_L[876][5] = l_cell_wire[857];							inform_L[845][5] = l_cell_wire[858];							inform_L[877][5] = l_cell_wire[859];							inform_L[846][5] = l_cell_wire[860];							inform_L[878][5] = l_cell_wire[861];							inform_L[847][5] = l_cell_wire[862];							inform_L[879][5] = l_cell_wire[863];							inform_L[848][5] = l_cell_wire[864];							inform_L[880][5] = l_cell_wire[865];							inform_L[849][5] = l_cell_wire[866];							inform_L[881][5] = l_cell_wire[867];							inform_L[850][5] = l_cell_wire[868];							inform_L[882][5] = l_cell_wire[869];							inform_L[851][5] = l_cell_wire[870];							inform_L[883][5] = l_cell_wire[871];							inform_L[852][5] = l_cell_wire[872];							inform_L[884][5] = l_cell_wire[873];							inform_L[853][5] = l_cell_wire[874];							inform_L[885][5] = l_cell_wire[875];							inform_L[854][5] = l_cell_wire[876];							inform_L[886][5] = l_cell_wire[877];							inform_L[855][5] = l_cell_wire[878];							inform_L[887][5] = l_cell_wire[879];							inform_L[856][5] = l_cell_wire[880];							inform_L[888][5] = l_cell_wire[881];							inform_L[857][5] = l_cell_wire[882];							inform_L[889][5] = l_cell_wire[883];							inform_L[858][5] = l_cell_wire[884];							inform_L[890][5] = l_cell_wire[885];							inform_L[859][5] = l_cell_wire[886];							inform_L[891][5] = l_cell_wire[887];							inform_L[860][5] = l_cell_wire[888];							inform_L[892][5] = l_cell_wire[889];							inform_L[861][5] = l_cell_wire[890];							inform_L[893][5] = l_cell_wire[891];							inform_L[862][5] = l_cell_wire[892];							inform_L[894][5] = l_cell_wire[893];							inform_L[863][5] = l_cell_wire[894];							inform_L[895][5] = l_cell_wire[895];							inform_L[896][5] = l_cell_wire[896];							inform_L[928][5] = l_cell_wire[897];							inform_L[897][5] = l_cell_wire[898];							inform_L[929][5] = l_cell_wire[899];							inform_L[898][5] = l_cell_wire[900];							inform_L[930][5] = l_cell_wire[901];							inform_L[899][5] = l_cell_wire[902];							inform_L[931][5] = l_cell_wire[903];							inform_L[900][5] = l_cell_wire[904];							inform_L[932][5] = l_cell_wire[905];							inform_L[901][5] = l_cell_wire[906];							inform_L[933][5] = l_cell_wire[907];							inform_L[902][5] = l_cell_wire[908];							inform_L[934][5] = l_cell_wire[909];							inform_L[903][5] = l_cell_wire[910];							inform_L[935][5] = l_cell_wire[911];							inform_L[904][5] = l_cell_wire[912];							inform_L[936][5] = l_cell_wire[913];							inform_L[905][5] = l_cell_wire[914];							inform_L[937][5] = l_cell_wire[915];							inform_L[906][5] = l_cell_wire[916];							inform_L[938][5] = l_cell_wire[917];							inform_L[907][5] = l_cell_wire[918];							inform_L[939][5] = l_cell_wire[919];							inform_L[908][5] = l_cell_wire[920];							inform_L[940][5] = l_cell_wire[921];							inform_L[909][5] = l_cell_wire[922];							inform_L[941][5] = l_cell_wire[923];							inform_L[910][5] = l_cell_wire[924];							inform_L[942][5] = l_cell_wire[925];							inform_L[911][5] = l_cell_wire[926];							inform_L[943][5] = l_cell_wire[927];							inform_L[912][5] = l_cell_wire[928];							inform_L[944][5] = l_cell_wire[929];							inform_L[913][5] = l_cell_wire[930];							inform_L[945][5] = l_cell_wire[931];							inform_L[914][5] = l_cell_wire[932];							inform_L[946][5] = l_cell_wire[933];							inform_L[915][5] = l_cell_wire[934];							inform_L[947][5] = l_cell_wire[935];							inform_L[916][5] = l_cell_wire[936];							inform_L[948][5] = l_cell_wire[937];							inform_L[917][5] = l_cell_wire[938];							inform_L[949][5] = l_cell_wire[939];							inform_L[918][5] = l_cell_wire[940];							inform_L[950][5] = l_cell_wire[941];							inform_L[919][5] = l_cell_wire[942];							inform_L[951][5] = l_cell_wire[943];							inform_L[920][5] = l_cell_wire[944];							inform_L[952][5] = l_cell_wire[945];							inform_L[921][5] = l_cell_wire[946];							inform_L[953][5] = l_cell_wire[947];							inform_L[922][5] = l_cell_wire[948];							inform_L[954][5] = l_cell_wire[949];							inform_L[923][5] = l_cell_wire[950];							inform_L[955][5] = l_cell_wire[951];							inform_L[924][5] = l_cell_wire[952];							inform_L[956][5] = l_cell_wire[953];							inform_L[925][5] = l_cell_wire[954];							inform_L[957][5] = l_cell_wire[955];							inform_L[926][5] = l_cell_wire[956];							inform_L[958][5] = l_cell_wire[957];							inform_L[927][5] = l_cell_wire[958];							inform_L[959][5] = l_cell_wire[959];							inform_L[960][5] = l_cell_wire[960];							inform_L[992][5] = l_cell_wire[961];							inform_L[961][5] = l_cell_wire[962];							inform_L[993][5] = l_cell_wire[963];							inform_L[962][5] = l_cell_wire[964];							inform_L[994][5] = l_cell_wire[965];							inform_L[963][5] = l_cell_wire[966];							inform_L[995][5] = l_cell_wire[967];							inform_L[964][5] = l_cell_wire[968];							inform_L[996][5] = l_cell_wire[969];							inform_L[965][5] = l_cell_wire[970];							inform_L[997][5] = l_cell_wire[971];							inform_L[966][5] = l_cell_wire[972];							inform_L[998][5] = l_cell_wire[973];							inform_L[967][5] = l_cell_wire[974];							inform_L[999][5] = l_cell_wire[975];							inform_L[968][5] = l_cell_wire[976];							inform_L[1000][5] = l_cell_wire[977];							inform_L[969][5] = l_cell_wire[978];							inform_L[1001][5] = l_cell_wire[979];							inform_L[970][5] = l_cell_wire[980];							inform_L[1002][5] = l_cell_wire[981];							inform_L[971][5] = l_cell_wire[982];							inform_L[1003][5] = l_cell_wire[983];							inform_L[972][5] = l_cell_wire[984];							inform_L[1004][5] = l_cell_wire[985];							inform_L[973][5] = l_cell_wire[986];							inform_L[1005][5] = l_cell_wire[987];							inform_L[974][5] = l_cell_wire[988];							inform_L[1006][5] = l_cell_wire[989];							inform_L[975][5] = l_cell_wire[990];							inform_L[1007][5] = l_cell_wire[991];							inform_L[976][5] = l_cell_wire[992];							inform_L[1008][5] = l_cell_wire[993];							inform_L[977][5] = l_cell_wire[994];							inform_L[1009][5] = l_cell_wire[995];							inform_L[978][5] = l_cell_wire[996];							inform_L[1010][5] = l_cell_wire[997];							inform_L[979][5] = l_cell_wire[998];							inform_L[1011][5] = l_cell_wire[999];							inform_L[980][5] = l_cell_wire[1000];							inform_L[1012][5] = l_cell_wire[1001];							inform_L[981][5] = l_cell_wire[1002];							inform_L[1013][5] = l_cell_wire[1003];							inform_L[982][5] = l_cell_wire[1004];							inform_L[1014][5] = l_cell_wire[1005];							inform_L[983][5] = l_cell_wire[1006];							inform_L[1015][5] = l_cell_wire[1007];							inform_L[984][5] = l_cell_wire[1008];							inform_L[1016][5] = l_cell_wire[1009];							inform_L[985][5] = l_cell_wire[1010];							inform_L[1017][5] = l_cell_wire[1011];							inform_L[986][5] = l_cell_wire[1012];							inform_L[1018][5] = l_cell_wire[1013];							inform_L[987][5] = l_cell_wire[1014];							inform_L[1019][5] = l_cell_wire[1015];							inform_L[988][5] = l_cell_wire[1016];							inform_L[1020][5] = l_cell_wire[1017];							inform_L[989][5] = l_cell_wire[1018];							inform_L[1021][5] = l_cell_wire[1019];							inform_L[990][5] = l_cell_wire[1020];							inform_L[1022][5] = l_cell_wire[1021];							inform_L[991][5] = l_cell_wire[1022];							inform_L[1023][5] = l_cell_wire[1023];						end
						7:						begin							inform_R[0][7] = r_cell_wire[0];							inform_R[64][7] = r_cell_wire[1];							inform_R[1][7] = r_cell_wire[2];							inform_R[65][7] = r_cell_wire[3];							inform_R[2][7] = r_cell_wire[4];							inform_R[66][7] = r_cell_wire[5];							inform_R[3][7] = r_cell_wire[6];							inform_R[67][7] = r_cell_wire[7];							inform_R[4][7] = r_cell_wire[8];							inform_R[68][7] = r_cell_wire[9];							inform_R[5][7] = r_cell_wire[10];							inform_R[69][7] = r_cell_wire[11];							inform_R[6][7] = r_cell_wire[12];							inform_R[70][7] = r_cell_wire[13];							inform_R[7][7] = r_cell_wire[14];							inform_R[71][7] = r_cell_wire[15];							inform_R[8][7] = r_cell_wire[16];							inform_R[72][7] = r_cell_wire[17];							inform_R[9][7] = r_cell_wire[18];							inform_R[73][7] = r_cell_wire[19];							inform_R[10][7] = r_cell_wire[20];							inform_R[74][7] = r_cell_wire[21];							inform_R[11][7] = r_cell_wire[22];							inform_R[75][7] = r_cell_wire[23];							inform_R[12][7] = r_cell_wire[24];							inform_R[76][7] = r_cell_wire[25];							inform_R[13][7] = r_cell_wire[26];							inform_R[77][7] = r_cell_wire[27];							inform_R[14][7] = r_cell_wire[28];							inform_R[78][7] = r_cell_wire[29];							inform_R[15][7] = r_cell_wire[30];							inform_R[79][7] = r_cell_wire[31];							inform_R[16][7] = r_cell_wire[32];							inform_R[80][7] = r_cell_wire[33];							inform_R[17][7] = r_cell_wire[34];							inform_R[81][7] = r_cell_wire[35];							inform_R[18][7] = r_cell_wire[36];							inform_R[82][7] = r_cell_wire[37];							inform_R[19][7] = r_cell_wire[38];							inform_R[83][7] = r_cell_wire[39];							inform_R[20][7] = r_cell_wire[40];							inform_R[84][7] = r_cell_wire[41];							inform_R[21][7] = r_cell_wire[42];							inform_R[85][7] = r_cell_wire[43];							inform_R[22][7] = r_cell_wire[44];							inform_R[86][7] = r_cell_wire[45];							inform_R[23][7] = r_cell_wire[46];							inform_R[87][7] = r_cell_wire[47];							inform_R[24][7] = r_cell_wire[48];							inform_R[88][7] = r_cell_wire[49];							inform_R[25][7] = r_cell_wire[50];							inform_R[89][7] = r_cell_wire[51];							inform_R[26][7] = r_cell_wire[52];							inform_R[90][7] = r_cell_wire[53];							inform_R[27][7] = r_cell_wire[54];							inform_R[91][7] = r_cell_wire[55];							inform_R[28][7] = r_cell_wire[56];							inform_R[92][7] = r_cell_wire[57];							inform_R[29][7] = r_cell_wire[58];							inform_R[93][7] = r_cell_wire[59];							inform_R[30][7] = r_cell_wire[60];							inform_R[94][7] = r_cell_wire[61];							inform_R[31][7] = r_cell_wire[62];							inform_R[95][7] = r_cell_wire[63];							inform_R[32][7] = r_cell_wire[64];							inform_R[96][7] = r_cell_wire[65];							inform_R[33][7] = r_cell_wire[66];							inform_R[97][7] = r_cell_wire[67];							inform_R[34][7] = r_cell_wire[68];							inform_R[98][7] = r_cell_wire[69];							inform_R[35][7] = r_cell_wire[70];							inform_R[99][7] = r_cell_wire[71];							inform_R[36][7] = r_cell_wire[72];							inform_R[100][7] = r_cell_wire[73];							inform_R[37][7] = r_cell_wire[74];							inform_R[101][7] = r_cell_wire[75];							inform_R[38][7] = r_cell_wire[76];							inform_R[102][7] = r_cell_wire[77];							inform_R[39][7] = r_cell_wire[78];							inform_R[103][7] = r_cell_wire[79];							inform_R[40][7] = r_cell_wire[80];							inform_R[104][7] = r_cell_wire[81];							inform_R[41][7] = r_cell_wire[82];							inform_R[105][7] = r_cell_wire[83];							inform_R[42][7] = r_cell_wire[84];							inform_R[106][7] = r_cell_wire[85];							inform_R[43][7] = r_cell_wire[86];							inform_R[107][7] = r_cell_wire[87];							inform_R[44][7] = r_cell_wire[88];							inform_R[108][7] = r_cell_wire[89];							inform_R[45][7] = r_cell_wire[90];							inform_R[109][7] = r_cell_wire[91];							inform_R[46][7] = r_cell_wire[92];							inform_R[110][7] = r_cell_wire[93];							inform_R[47][7] = r_cell_wire[94];							inform_R[111][7] = r_cell_wire[95];							inform_R[48][7] = r_cell_wire[96];							inform_R[112][7] = r_cell_wire[97];							inform_R[49][7] = r_cell_wire[98];							inform_R[113][7] = r_cell_wire[99];							inform_R[50][7] = r_cell_wire[100];							inform_R[114][7] = r_cell_wire[101];							inform_R[51][7] = r_cell_wire[102];							inform_R[115][7] = r_cell_wire[103];							inform_R[52][7] = r_cell_wire[104];							inform_R[116][7] = r_cell_wire[105];							inform_R[53][7] = r_cell_wire[106];							inform_R[117][7] = r_cell_wire[107];							inform_R[54][7] = r_cell_wire[108];							inform_R[118][7] = r_cell_wire[109];							inform_R[55][7] = r_cell_wire[110];							inform_R[119][7] = r_cell_wire[111];							inform_R[56][7] = r_cell_wire[112];							inform_R[120][7] = r_cell_wire[113];							inform_R[57][7] = r_cell_wire[114];							inform_R[121][7] = r_cell_wire[115];							inform_R[58][7] = r_cell_wire[116];							inform_R[122][7] = r_cell_wire[117];							inform_R[59][7] = r_cell_wire[118];							inform_R[123][7] = r_cell_wire[119];							inform_R[60][7] = r_cell_wire[120];							inform_R[124][7] = r_cell_wire[121];							inform_R[61][7] = r_cell_wire[122];							inform_R[125][7] = r_cell_wire[123];							inform_R[62][7] = r_cell_wire[124];							inform_R[126][7] = r_cell_wire[125];							inform_R[63][7] = r_cell_wire[126];							inform_R[127][7] = r_cell_wire[127];							inform_R[128][7] = r_cell_wire[128];							inform_R[192][7] = r_cell_wire[129];							inform_R[129][7] = r_cell_wire[130];							inform_R[193][7] = r_cell_wire[131];							inform_R[130][7] = r_cell_wire[132];							inform_R[194][7] = r_cell_wire[133];							inform_R[131][7] = r_cell_wire[134];							inform_R[195][7] = r_cell_wire[135];							inform_R[132][7] = r_cell_wire[136];							inform_R[196][7] = r_cell_wire[137];							inform_R[133][7] = r_cell_wire[138];							inform_R[197][7] = r_cell_wire[139];							inform_R[134][7] = r_cell_wire[140];							inform_R[198][7] = r_cell_wire[141];							inform_R[135][7] = r_cell_wire[142];							inform_R[199][7] = r_cell_wire[143];							inform_R[136][7] = r_cell_wire[144];							inform_R[200][7] = r_cell_wire[145];							inform_R[137][7] = r_cell_wire[146];							inform_R[201][7] = r_cell_wire[147];							inform_R[138][7] = r_cell_wire[148];							inform_R[202][7] = r_cell_wire[149];							inform_R[139][7] = r_cell_wire[150];							inform_R[203][7] = r_cell_wire[151];							inform_R[140][7] = r_cell_wire[152];							inform_R[204][7] = r_cell_wire[153];							inform_R[141][7] = r_cell_wire[154];							inform_R[205][7] = r_cell_wire[155];							inform_R[142][7] = r_cell_wire[156];							inform_R[206][7] = r_cell_wire[157];							inform_R[143][7] = r_cell_wire[158];							inform_R[207][7] = r_cell_wire[159];							inform_R[144][7] = r_cell_wire[160];							inform_R[208][7] = r_cell_wire[161];							inform_R[145][7] = r_cell_wire[162];							inform_R[209][7] = r_cell_wire[163];							inform_R[146][7] = r_cell_wire[164];							inform_R[210][7] = r_cell_wire[165];							inform_R[147][7] = r_cell_wire[166];							inform_R[211][7] = r_cell_wire[167];							inform_R[148][7] = r_cell_wire[168];							inform_R[212][7] = r_cell_wire[169];							inform_R[149][7] = r_cell_wire[170];							inform_R[213][7] = r_cell_wire[171];							inform_R[150][7] = r_cell_wire[172];							inform_R[214][7] = r_cell_wire[173];							inform_R[151][7] = r_cell_wire[174];							inform_R[215][7] = r_cell_wire[175];							inform_R[152][7] = r_cell_wire[176];							inform_R[216][7] = r_cell_wire[177];							inform_R[153][7] = r_cell_wire[178];							inform_R[217][7] = r_cell_wire[179];							inform_R[154][7] = r_cell_wire[180];							inform_R[218][7] = r_cell_wire[181];							inform_R[155][7] = r_cell_wire[182];							inform_R[219][7] = r_cell_wire[183];							inform_R[156][7] = r_cell_wire[184];							inform_R[220][7] = r_cell_wire[185];							inform_R[157][7] = r_cell_wire[186];							inform_R[221][7] = r_cell_wire[187];							inform_R[158][7] = r_cell_wire[188];							inform_R[222][7] = r_cell_wire[189];							inform_R[159][7] = r_cell_wire[190];							inform_R[223][7] = r_cell_wire[191];							inform_R[160][7] = r_cell_wire[192];							inform_R[224][7] = r_cell_wire[193];							inform_R[161][7] = r_cell_wire[194];							inform_R[225][7] = r_cell_wire[195];							inform_R[162][7] = r_cell_wire[196];							inform_R[226][7] = r_cell_wire[197];							inform_R[163][7] = r_cell_wire[198];							inform_R[227][7] = r_cell_wire[199];							inform_R[164][7] = r_cell_wire[200];							inform_R[228][7] = r_cell_wire[201];							inform_R[165][7] = r_cell_wire[202];							inform_R[229][7] = r_cell_wire[203];							inform_R[166][7] = r_cell_wire[204];							inform_R[230][7] = r_cell_wire[205];							inform_R[167][7] = r_cell_wire[206];							inform_R[231][7] = r_cell_wire[207];							inform_R[168][7] = r_cell_wire[208];							inform_R[232][7] = r_cell_wire[209];							inform_R[169][7] = r_cell_wire[210];							inform_R[233][7] = r_cell_wire[211];							inform_R[170][7] = r_cell_wire[212];							inform_R[234][7] = r_cell_wire[213];							inform_R[171][7] = r_cell_wire[214];							inform_R[235][7] = r_cell_wire[215];							inform_R[172][7] = r_cell_wire[216];							inform_R[236][7] = r_cell_wire[217];							inform_R[173][7] = r_cell_wire[218];							inform_R[237][7] = r_cell_wire[219];							inform_R[174][7] = r_cell_wire[220];							inform_R[238][7] = r_cell_wire[221];							inform_R[175][7] = r_cell_wire[222];							inform_R[239][7] = r_cell_wire[223];							inform_R[176][7] = r_cell_wire[224];							inform_R[240][7] = r_cell_wire[225];							inform_R[177][7] = r_cell_wire[226];							inform_R[241][7] = r_cell_wire[227];							inform_R[178][7] = r_cell_wire[228];							inform_R[242][7] = r_cell_wire[229];							inform_R[179][7] = r_cell_wire[230];							inform_R[243][7] = r_cell_wire[231];							inform_R[180][7] = r_cell_wire[232];							inform_R[244][7] = r_cell_wire[233];							inform_R[181][7] = r_cell_wire[234];							inform_R[245][7] = r_cell_wire[235];							inform_R[182][7] = r_cell_wire[236];							inform_R[246][7] = r_cell_wire[237];							inform_R[183][7] = r_cell_wire[238];							inform_R[247][7] = r_cell_wire[239];							inform_R[184][7] = r_cell_wire[240];							inform_R[248][7] = r_cell_wire[241];							inform_R[185][7] = r_cell_wire[242];							inform_R[249][7] = r_cell_wire[243];							inform_R[186][7] = r_cell_wire[244];							inform_R[250][7] = r_cell_wire[245];							inform_R[187][7] = r_cell_wire[246];							inform_R[251][7] = r_cell_wire[247];							inform_R[188][7] = r_cell_wire[248];							inform_R[252][7] = r_cell_wire[249];							inform_R[189][7] = r_cell_wire[250];							inform_R[253][7] = r_cell_wire[251];							inform_R[190][7] = r_cell_wire[252];							inform_R[254][7] = r_cell_wire[253];							inform_R[191][7] = r_cell_wire[254];							inform_R[255][7] = r_cell_wire[255];							inform_R[256][7] = r_cell_wire[256];							inform_R[320][7] = r_cell_wire[257];							inform_R[257][7] = r_cell_wire[258];							inform_R[321][7] = r_cell_wire[259];							inform_R[258][7] = r_cell_wire[260];							inform_R[322][7] = r_cell_wire[261];							inform_R[259][7] = r_cell_wire[262];							inform_R[323][7] = r_cell_wire[263];							inform_R[260][7] = r_cell_wire[264];							inform_R[324][7] = r_cell_wire[265];							inform_R[261][7] = r_cell_wire[266];							inform_R[325][7] = r_cell_wire[267];							inform_R[262][7] = r_cell_wire[268];							inform_R[326][7] = r_cell_wire[269];							inform_R[263][7] = r_cell_wire[270];							inform_R[327][7] = r_cell_wire[271];							inform_R[264][7] = r_cell_wire[272];							inform_R[328][7] = r_cell_wire[273];							inform_R[265][7] = r_cell_wire[274];							inform_R[329][7] = r_cell_wire[275];							inform_R[266][7] = r_cell_wire[276];							inform_R[330][7] = r_cell_wire[277];							inform_R[267][7] = r_cell_wire[278];							inform_R[331][7] = r_cell_wire[279];							inform_R[268][7] = r_cell_wire[280];							inform_R[332][7] = r_cell_wire[281];							inform_R[269][7] = r_cell_wire[282];							inform_R[333][7] = r_cell_wire[283];							inform_R[270][7] = r_cell_wire[284];							inform_R[334][7] = r_cell_wire[285];							inform_R[271][7] = r_cell_wire[286];							inform_R[335][7] = r_cell_wire[287];							inform_R[272][7] = r_cell_wire[288];							inform_R[336][7] = r_cell_wire[289];							inform_R[273][7] = r_cell_wire[290];							inform_R[337][7] = r_cell_wire[291];							inform_R[274][7] = r_cell_wire[292];							inform_R[338][7] = r_cell_wire[293];							inform_R[275][7] = r_cell_wire[294];							inform_R[339][7] = r_cell_wire[295];							inform_R[276][7] = r_cell_wire[296];							inform_R[340][7] = r_cell_wire[297];							inform_R[277][7] = r_cell_wire[298];							inform_R[341][7] = r_cell_wire[299];							inform_R[278][7] = r_cell_wire[300];							inform_R[342][7] = r_cell_wire[301];							inform_R[279][7] = r_cell_wire[302];							inform_R[343][7] = r_cell_wire[303];							inform_R[280][7] = r_cell_wire[304];							inform_R[344][7] = r_cell_wire[305];							inform_R[281][7] = r_cell_wire[306];							inform_R[345][7] = r_cell_wire[307];							inform_R[282][7] = r_cell_wire[308];							inform_R[346][7] = r_cell_wire[309];							inform_R[283][7] = r_cell_wire[310];							inform_R[347][7] = r_cell_wire[311];							inform_R[284][7] = r_cell_wire[312];							inform_R[348][7] = r_cell_wire[313];							inform_R[285][7] = r_cell_wire[314];							inform_R[349][7] = r_cell_wire[315];							inform_R[286][7] = r_cell_wire[316];							inform_R[350][7] = r_cell_wire[317];							inform_R[287][7] = r_cell_wire[318];							inform_R[351][7] = r_cell_wire[319];							inform_R[288][7] = r_cell_wire[320];							inform_R[352][7] = r_cell_wire[321];							inform_R[289][7] = r_cell_wire[322];							inform_R[353][7] = r_cell_wire[323];							inform_R[290][7] = r_cell_wire[324];							inform_R[354][7] = r_cell_wire[325];							inform_R[291][7] = r_cell_wire[326];							inform_R[355][7] = r_cell_wire[327];							inform_R[292][7] = r_cell_wire[328];							inform_R[356][7] = r_cell_wire[329];							inform_R[293][7] = r_cell_wire[330];							inform_R[357][7] = r_cell_wire[331];							inform_R[294][7] = r_cell_wire[332];							inform_R[358][7] = r_cell_wire[333];							inform_R[295][7] = r_cell_wire[334];							inform_R[359][7] = r_cell_wire[335];							inform_R[296][7] = r_cell_wire[336];							inform_R[360][7] = r_cell_wire[337];							inform_R[297][7] = r_cell_wire[338];							inform_R[361][7] = r_cell_wire[339];							inform_R[298][7] = r_cell_wire[340];							inform_R[362][7] = r_cell_wire[341];							inform_R[299][7] = r_cell_wire[342];							inform_R[363][7] = r_cell_wire[343];							inform_R[300][7] = r_cell_wire[344];							inform_R[364][7] = r_cell_wire[345];							inform_R[301][7] = r_cell_wire[346];							inform_R[365][7] = r_cell_wire[347];							inform_R[302][7] = r_cell_wire[348];							inform_R[366][7] = r_cell_wire[349];							inform_R[303][7] = r_cell_wire[350];							inform_R[367][7] = r_cell_wire[351];							inform_R[304][7] = r_cell_wire[352];							inform_R[368][7] = r_cell_wire[353];							inform_R[305][7] = r_cell_wire[354];							inform_R[369][7] = r_cell_wire[355];							inform_R[306][7] = r_cell_wire[356];							inform_R[370][7] = r_cell_wire[357];							inform_R[307][7] = r_cell_wire[358];							inform_R[371][7] = r_cell_wire[359];							inform_R[308][7] = r_cell_wire[360];							inform_R[372][7] = r_cell_wire[361];							inform_R[309][7] = r_cell_wire[362];							inform_R[373][7] = r_cell_wire[363];							inform_R[310][7] = r_cell_wire[364];							inform_R[374][7] = r_cell_wire[365];							inform_R[311][7] = r_cell_wire[366];							inform_R[375][7] = r_cell_wire[367];							inform_R[312][7] = r_cell_wire[368];							inform_R[376][7] = r_cell_wire[369];							inform_R[313][7] = r_cell_wire[370];							inform_R[377][7] = r_cell_wire[371];							inform_R[314][7] = r_cell_wire[372];							inform_R[378][7] = r_cell_wire[373];							inform_R[315][7] = r_cell_wire[374];							inform_R[379][7] = r_cell_wire[375];							inform_R[316][7] = r_cell_wire[376];							inform_R[380][7] = r_cell_wire[377];							inform_R[317][7] = r_cell_wire[378];							inform_R[381][7] = r_cell_wire[379];							inform_R[318][7] = r_cell_wire[380];							inform_R[382][7] = r_cell_wire[381];							inform_R[319][7] = r_cell_wire[382];							inform_R[383][7] = r_cell_wire[383];							inform_R[384][7] = r_cell_wire[384];							inform_R[448][7] = r_cell_wire[385];							inform_R[385][7] = r_cell_wire[386];							inform_R[449][7] = r_cell_wire[387];							inform_R[386][7] = r_cell_wire[388];							inform_R[450][7] = r_cell_wire[389];							inform_R[387][7] = r_cell_wire[390];							inform_R[451][7] = r_cell_wire[391];							inform_R[388][7] = r_cell_wire[392];							inform_R[452][7] = r_cell_wire[393];							inform_R[389][7] = r_cell_wire[394];							inform_R[453][7] = r_cell_wire[395];							inform_R[390][7] = r_cell_wire[396];							inform_R[454][7] = r_cell_wire[397];							inform_R[391][7] = r_cell_wire[398];							inform_R[455][7] = r_cell_wire[399];							inform_R[392][7] = r_cell_wire[400];							inform_R[456][7] = r_cell_wire[401];							inform_R[393][7] = r_cell_wire[402];							inform_R[457][7] = r_cell_wire[403];							inform_R[394][7] = r_cell_wire[404];							inform_R[458][7] = r_cell_wire[405];							inform_R[395][7] = r_cell_wire[406];							inform_R[459][7] = r_cell_wire[407];							inform_R[396][7] = r_cell_wire[408];							inform_R[460][7] = r_cell_wire[409];							inform_R[397][7] = r_cell_wire[410];							inform_R[461][7] = r_cell_wire[411];							inform_R[398][7] = r_cell_wire[412];							inform_R[462][7] = r_cell_wire[413];							inform_R[399][7] = r_cell_wire[414];							inform_R[463][7] = r_cell_wire[415];							inform_R[400][7] = r_cell_wire[416];							inform_R[464][7] = r_cell_wire[417];							inform_R[401][7] = r_cell_wire[418];							inform_R[465][7] = r_cell_wire[419];							inform_R[402][7] = r_cell_wire[420];							inform_R[466][7] = r_cell_wire[421];							inform_R[403][7] = r_cell_wire[422];							inform_R[467][7] = r_cell_wire[423];							inform_R[404][7] = r_cell_wire[424];							inform_R[468][7] = r_cell_wire[425];							inform_R[405][7] = r_cell_wire[426];							inform_R[469][7] = r_cell_wire[427];							inform_R[406][7] = r_cell_wire[428];							inform_R[470][7] = r_cell_wire[429];							inform_R[407][7] = r_cell_wire[430];							inform_R[471][7] = r_cell_wire[431];							inform_R[408][7] = r_cell_wire[432];							inform_R[472][7] = r_cell_wire[433];							inform_R[409][7] = r_cell_wire[434];							inform_R[473][7] = r_cell_wire[435];							inform_R[410][7] = r_cell_wire[436];							inform_R[474][7] = r_cell_wire[437];							inform_R[411][7] = r_cell_wire[438];							inform_R[475][7] = r_cell_wire[439];							inform_R[412][7] = r_cell_wire[440];							inform_R[476][7] = r_cell_wire[441];							inform_R[413][7] = r_cell_wire[442];							inform_R[477][7] = r_cell_wire[443];							inform_R[414][7] = r_cell_wire[444];							inform_R[478][7] = r_cell_wire[445];							inform_R[415][7] = r_cell_wire[446];							inform_R[479][7] = r_cell_wire[447];							inform_R[416][7] = r_cell_wire[448];							inform_R[480][7] = r_cell_wire[449];							inform_R[417][7] = r_cell_wire[450];							inform_R[481][7] = r_cell_wire[451];							inform_R[418][7] = r_cell_wire[452];							inform_R[482][7] = r_cell_wire[453];							inform_R[419][7] = r_cell_wire[454];							inform_R[483][7] = r_cell_wire[455];							inform_R[420][7] = r_cell_wire[456];							inform_R[484][7] = r_cell_wire[457];							inform_R[421][7] = r_cell_wire[458];							inform_R[485][7] = r_cell_wire[459];							inform_R[422][7] = r_cell_wire[460];							inform_R[486][7] = r_cell_wire[461];							inform_R[423][7] = r_cell_wire[462];							inform_R[487][7] = r_cell_wire[463];							inform_R[424][7] = r_cell_wire[464];							inform_R[488][7] = r_cell_wire[465];							inform_R[425][7] = r_cell_wire[466];							inform_R[489][7] = r_cell_wire[467];							inform_R[426][7] = r_cell_wire[468];							inform_R[490][7] = r_cell_wire[469];							inform_R[427][7] = r_cell_wire[470];							inform_R[491][7] = r_cell_wire[471];							inform_R[428][7] = r_cell_wire[472];							inform_R[492][7] = r_cell_wire[473];							inform_R[429][7] = r_cell_wire[474];							inform_R[493][7] = r_cell_wire[475];							inform_R[430][7] = r_cell_wire[476];							inform_R[494][7] = r_cell_wire[477];							inform_R[431][7] = r_cell_wire[478];							inform_R[495][7] = r_cell_wire[479];							inform_R[432][7] = r_cell_wire[480];							inform_R[496][7] = r_cell_wire[481];							inform_R[433][7] = r_cell_wire[482];							inform_R[497][7] = r_cell_wire[483];							inform_R[434][7] = r_cell_wire[484];							inform_R[498][7] = r_cell_wire[485];							inform_R[435][7] = r_cell_wire[486];							inform_R[499][7] = r_cell_wire[487];							inform_R[436][7] = r_cell_wire[488];							inform_R[500][7] = r_cell_wire[489];							inform_R[437][7] = r_cell_wire[490];							inform_R[501][7] = r_cell_wire[491];							inform_R[438][7] = r_cell_wire[492];							inform_R[502][7] = r_cell_wire[493];							inform_R[439][7] = r_cell_wire[494];							inform_R[503][7] = r_cell_wire[495];							inform_R[440][7] = r_cell_wire[496];							inform_R[504][7] = r_cell_wire[497];							inform_R[441][7] = r_cell_wire[498];							inform_R[505][7] = r_cell_wire[499];							inform_R[442][7] = r_cell_wire[500];							inform_R[506][7] = r_cell_wire[501];							inform_R[443][7] = r_cell_wire[502];							inform_R[507][7] = r_cell_wire[503];							inform_R[444][7] = r_cell_wire[504];							inform_R[508][7] = r_cell_wire[505];							inform_R[445][7] = r_cell_wire[506];							inform_R[509][7] = r_cell_wire[507];							inform_R[446][7] = r_cell_wire[508];							inform_R[510][7] = r_cell_wire[509];							inform_R[447][7] = r_cell_wire[510];							inform_R[511][7] = r_cell_wire[511];							inform_R[512][7] = r_cell_wire[512];							inform_R[576][7] = r_cell_wire[513];							inform_R[513][7] = r_cell_wire[514];							inform_R[577][7] = r_cell_wire[515];							inform_R[514][7] = r_cell_wire[516];							inform_R[578][7] = r_cell_wire[517];							inform_R[515][7] = r_cell_wire[518];							inform_R[579][7] = r_cell_wire[519];							inform_R[516][7] = r_cell_wire[520];							inform_R[580][7] = r_cell_wire[521];							inform_R[517][7] = r_cell_wire[522];							inform_R[581][7] = r_cell_wire[523];							inform_R[518][7] = r_cell_wire[524];							inform_R[582][7] = r_cell_wire[525];							inform_R[519][7] = r_cell_wire[526];							inform_R[583][7] = r_cell_wire[527];							inform_R[520][7] = r_cell_wire[528];							inform_R[584][7] = r_cell_wire[529];							inform_R[521][7] = r_cell_wire[530];							inform_R[585][7] = r_cell_wire[531];							inform_R[522][7] = r_cell_wire[532];							inform_R[586][7] = r_cell_wire[533];							inform_R[523][7] = r_cell_wire[534];							inform_R[587][7] = r_cell_wire[535];							inform_R[524][7] = r_cell_wire[536];							inform_R[588][7] = r_cell_wire[537];							inform_R[525][7] = r_cell_wire[538];							inform_R[589][7] = r_cell_wire[539];							inform_R[526][7] = r_cell_wire[540];							inform_R[590][7] = r_cell_wire[541];							inform_R[527][7] = r_cell_wire[542];							inform_R[591][7] = r_cell_wire[543];							inform_R[528][7] = r_cell_wire[544];							inform_R[592][7] = r_cell_wire[545];							inform_R[529][7] = r_cell_wire[546];							inform_R[593][7] = r_cell_wire[547];							inform_R[530][7] = r_cell_wire[548];							inform_R[594][7] = r_cell_wire[549];							inform_R[531][7] = r_cell_wire[550];							inform_R[595][7] = r_cell_wire[551];							inform_R[532][7] = r_cell_wire[552];							inform_R[596][7] = r_cell_wire[553];							inform_R[533][7] = r_cell_wire[554];							inform_R[597][7] = r_cell_wire[555];							inform_R[534][7] = r_cell_wire[556];							inform_R[598][7] = r_cell_wire[557];							inform_R[535][7] = r_cell_wire[558];							inform_R[599][7] = r_cell_wire[559];							inform_R[536][7] = r_cell_wire[560];							inform_R[600][7] = r_cell_wire[561];							inform_R[537][7] = r_cell_wire[562];							inform_R[601][7] = r_cell_wire[563];							inform_R[538][7] = r_cell_wire[564];							inform_R[602][7] = r_cell_wire[565];							inform_R[539][7] = r_cell_wire[566];							inform_R[603][7] = r_cell_wire[567];							inform_R[540][7] = r_cell_wire[568];							inform_R[604][7] = r_cell_wire[569];							inform_R[541][7] = r_cell_wire[570];							inform_R[605][7] = r_cell_wire[571];							inform_R[542][7] = r_cell_wire[572];							inform_R[606][7] = r_cell_wire[573];							inform_R[543][7] = r_cell_wire[574];							inform_R[607][7] = r_cell_wire[575];							inform_R[544][7] = r_cell_wire[576];							inform_R[608][7] = r_cell_wire[577];							inform_R[545][7] = r_cell_wire[578];							inform_R[609][7] = r_cell_wire[579];							inform_R[546][7] = r_cell_wire[580];							inform_R[610][7] = r_cell_wire[581];							inform_R[547][7] = r_cell_wire[582];							inform_R[611][7] = r_cell_wire[583];							inform_R[548][7] = r_cell_wire[584];							inform_R[612][7] = r_cell_wire[585];							inform_R[549][7] = r_cell_wire[586];							inform_R[613][7] = r_cell_wire[587];							inform_R[550][7] = r_cell_wire[588];							inform_R[614][7] = r_cell_wire[589];							inform_R[551][7] = r_cell_wire[590];							inform_R[615][7] = r_cell_wire[591];							inform_R[552][7] = r_cell_wire[592];							inform_R[616][7] = r_cell_wire[593];							inform_R[553][7] = r_cell_wire[594];							inform_R[617][7] = r_cell_wire[595];							inform_R[554][7] = r_cell_wire[596];							inform_R[618][7] = r_cell_wire[597];							inform_R[555][7] = r_cell_wire[598];							inform_R[619][7] = r_cell_wire[599];							inform_R[556][7] = r_cell_wire[600];							inform_R[620][7] = r_cell_wire[601];							inform_R[557][7] = r_cell_wire[602];							inform_R[621][7] = r_cell_wire[603];							inform_R[558][7] = r_cell_wire[604];							inform_R[622][7] = r_cell_wire[605];							inform_R[559][7] = r_cell_wire[606];							inform_R[623][7] = r_cell_wire[607];							inform_R[560][7] = r_cell_wire[608];							inform_R[624][7] = r_cell_wire[609];							inform_R[561][7] = r_cell_wire[610];							inform_R[625][7] = r_cell_wire[611];							inform_R[562][7] = r_cell_wire[612];							inform_R[626][7] = r_cell_wire[613];							inform_R[563][7] = r_cell_wire[614];							inform_R[627][7] = r_cell_wire[615];							inform_R[564][7] = r_cell_wire[616];							inform_R[628][7] = r_cell_wire[617];							inform_R[565][7] = r_cell_wire[618];							inform_R[629][7] = r_cell_wire[619];							inform_R[566][7] = r_cell_wire[620];							inform_R[630][7] = r_cell_wire[621];							inform_R[567][7] = r_cell_wire[622];							inform_R[631][7] = r_cell_wire[623];							inform_R[568][7] = r_cell_wire[624];							inform_R[632][7] = r_cell_wire[625];							inform_R[569][7] = r_cell_wire[626];							inform_R[633][7] = r_cell_wire[627];							inform_R[570][7] = r_cell_wire[628];							inform_R[634][7] = r_cell_wire[629];							inform_R[571][7] = r_cell_wire[630];							inform_R[635][7] = r_cell_wire[631];							inform_R[572][7] = r_cell_wire[632];							inform_R[636][7] = r_cell_wire[633];							inform_R[573][7] = r_cell_wire[634];							inform_R[637][7] = r_cell_wire[635];							inform_R[574][7] = r_cell_wire[636];							inform_R[638][7] = r_cell_wire[637];							inform_R[575][7] = r_cell_wire[638];							inform_R[639][7] = r_cell_wire[639];							inform_R[640][7] = r_cell_wire[640];							inform_R[704][7] = r_cell_wire[641];							inform_R[641][7] = r_cell_wire[642];							inform_R[705][7] = r_cell_wire[643];							inform_R[642][7] = r_cell_wire[644];							inform_R[706][7] = r_cell_wire[645];							inform_R[643][7] = r_cell_wire[646];							inform_R[707][7] = r_cell_wire[647];							inform_R[644][7] = r_cell_wire[648];							inform_R[708][7] = r_cell_wire[649];							inform_R[645][7] = r_cell_wire[650];							inform_R[709][7] = r_cell_wire[651];							inform_R[646][7] = r_cell_wire[652];							inform_R[710][7] = r_cell_wire[653];							inform_R[647][7] = r_cell_wire[654];							inform_R[711][7] = r_cell_wire[655];							inform_R[648][7] = r_cell_wire[656];							inform_R[712][7] = r_cell_wire[657];							inform_R[649][7] = r_cell_wire[658];							inform_R[713][7] = r_cell_wire[659];							inform_R[650][7] = r_cell_wire[660];							inform_R[714][7] = r_cell_wire[661];							inform_R[651][7] = r_cell_wire[662];							inform_R[715][7] = r_cell_wire[663];							inform_R[652][7] = r_cell_wire[664];							inform_R[716][7] = r_cell_wire[665];							inform_R[653][7] = r_cell_wire[666];							inform_R[717][7] = r_cell_wire[667];							inform_R[654][7] = r_cell_wire[668];							inform_R[718][7] = r_cell_wire[669];							inform_R[655][7] = r_cell_wire[670];							inform_R[719][7] = r_cell_wire[671];							inform_R[656][7] = r_cell_wire[672];							inform_R[720][7] = r_cell_wire[673];							inform_R[657][7] = r_cell_wire[674];							inform_R[721][7] = r_cell_wire[675];							inform_R[658][7] = r_cell_wire[676];							inform_R[722][7] = r_cell_wire[677];							inform_R[659][7] = r_cell_wire[678];							inform_R[723][7] = r_cell_wire[679];							inform_R[660][7] = r_cell_wire[680];							inform_R[724][7] = r_cell_wire[681];							inform_R[661][7] = r_cell_wire[682];							inform_R[725][7] = r_cell_wire[683];							inform_R[662][7] = r_cell_wire[684];							inform_R[726][7] = r_cell_wire[685];							inform_R[663][7] = r_cell_wire[686];							inform_R[727][7] = r_cell_wire[687];							inform_R[664][7] = r_cell_wire[688];							inform_R[728][7] = r_cell_wire[689];							inform_R[665][7] = r_cell_wire[690];							inform_R[729][7] = r_cell_wire[691];							inform_R[666][7] = r_cell_wire[692];							inform_R[730][7] = r_cell_wire[693];							inform_R[667][7] = r_cell_wire[694];							inform_R[731][7] = r_cell_wire[695];							inform_R[668][7] = r_cell_wire[696];							inform_R[732][7] = r_cell_wire[697];							inform_R[669][7] = r_cell_wire[698];							inform_R[733][7] = r_cell_wire[699];							inform_R[670][7] = r_cell_wire[700];							inform_R[734][7] = r_cell_wire[701];							inform_R[671][7] = r_cell_wire[702];							inform_R[735][7] = r_cell_wire[703];							inform_R[672][7] = r_cell_wire[704];							inform_R[736][7] = r_cell_wire[705];							inform_R[673][7] = r_cell_wire[706];							inform_R[737][7] = r_cell_wire[707];							inform_R[674][7] = r_cell_wire[708];							inform_R[738][7] = r_cell_wire[709];							inform_R[675][7] = r_cell_wire[710];							inform_R[739][7] = r_cell_wire[711];							inform_R[676][7] = r_cell_wire[712];							inform_R[740][7] = r_cell_wire[713];							inform_R[677][7] = r_cell_wire[714];							inform_R[741][7] = r_cell_wire[715];							inform_R[678][7] = r_cell_wire[716];							inform_R[742][7] = r_cell_wire[717];							inform_R[679][7] = r_cell_wire[718];							inform_R[743][7] = r_cell_wire[719];							inform_R[680][7] = r_cell_wire[720];							inform_R[744][7] = r_cell_wire[721];							inform_R[681][7] = r_cell_wire[722];							inform_R[745][7] = r_cell_wire[723];							inform_R[682][7] = r_cell_wire[724];							inform_R[746][7] = r_cell_wire[725];							inform_R[683][7] = r_cell_wire[726];							inform_R[747][7] = r_cell_wire[727];							inform_R[684][7] = r_cell_wire[728];							inform_R[748][7] = r_cell_wire[729];							inform_R[685][7] = r_cell_wire[730];							inform_R[749][7] = r_cell_wire[731];							inform_R[686][7] = r_cell_wire[732];							inform_R[750][7] = r_cell_wire[733];							inform_R[687][7] = r_cell_wire[734];							inform_R[751][7] = r_cell_wire[735];							inform_R[688][7] = r_cell_wire[736];							inform_R[752][7] = r_cell_wire[737];							inform_R[689][7] = r_cell_wire[738];							inform_R[753][7] = r_cell_wire[739];							inform_R[690][7] = r_cell_wire[740];							inform_R[754][7] = r_cell_wire[741];							inform_R[691][7] = r_cell_wire[742];							inform_R[755][7] = r_cell_wire[743];							inform_R[692][7] = r_cell_wire[744];							inform_R[756][7] = r_cell_wire[745];							inform_R[693][7] = r_cell_wire[746];							inform_R[757][7] = r_cell_wire[747];							inform_R[694][7] = r_cell_wire[748];							inform_R[758][7] = r_cell_wire[749];							inform_R[695][7] = r_cell_wire[750];							inform_R[759][7] = r_cell_wire[751];							inform_R[696][7] = r_cell_wire[752];							inform_R[760][7] = r_cell_wire[753];							inform_R[697][7] = r_cell_wire[754];							inform_R[761][7] = r_cell_wire[755];							inform_R[698][7] = r_cell_wire[756];							inform_R[762][7] = r_cell_wire[757];							inform_R[699][7] = r_cell_wire[758];							inform_R[763][7] = r_cell_wire[759];							inform_R[700][7] = r_cell_wire[760];							inform_R[764][7] = r_cell_wire[761];							inform_R[701][7] = r_cell_wire[762];							inform_R[765][7] = r_cell_wire[763];							inform_R[702][7] = r_cell_wire[764];							inform_R[766][7] = r_cell_wire[765];							inform_R[703][7] = r_cell_wire[766];							inform_R[767][7] = r_cell_wire[767];							inform_R[768][7] = r_cell_wire[768];							inform_R[832][7] = r_cell_wire[769];							inform_R[769][7] = r_cell_wire[770];							inform_R[833][7] = r_cell_wire[771];							inform_R[770][7] = r_cell_wire[772];							inform_R[834][7] = r_cell_wire[773];							inform_R[771][7] = r_cell_wire[774];							inform_R[835][7] = r_cell_wire[775];							inform_R[772][7] = r_cell_wire[776];							inform_R[836][7] = r_cell_wire[777];							inform_R[773][7] = r_cell_wire[778];							inform_R[837][7] = r_cell_wire[779];							inform_R[774][7] = r_cell_wire[780];							inform_R[838][7] = r_cell_wire[781];							inform_R[775][7] = r_cell_wire[782];							inform_R[839][7] = r_cell_wire[783];							inform_R[776][7] = r_cell_wire[784];							inform_R[840][7] = r_cell_wire[785];							inform_R[777][7] = r_cell_wire[786];							inform_R[841][7] = r_cell_wire[787];							inform_R[778][7] = r_cell_wire[788];							inform_R[842][7] = r_cell_wire[789];							inform_R[779][7] = r_cell_wire[790];							inform_R[843][7] = r_cell_wire[791];							inform_R[780][7] = r_cell_wire[792];							inform_R[844][7] = r_cell_wire[793];							inform_R[781][7] = r_cell_wire[794];							inform_R[845][7] = r_cell_wire[795];							inform_R[782][7] = r_cell_wire[796];							inform_R[846][7] = r_cell_wire[797];							inform_R[783][7] = r_cell_wire[798];							inform_R[847][7] = r_cell_wire[799];							inform_R[784][7] = r_cell_wire[800];							inform_R[848][7] = r_cell_wire[801];							inform_R[785][7] = r_cell_wire[802];							inform_R[849][7] = r_cell_wire[803];							inform_R[786][7] = r_cell_wire[804];							inform_R[850][7] = r_cell_wire[805];							inform_R[787][7] = r_cell_wire[806];							inform_R[851][7] = r_cell_wire[807];							inform_R[788][7] = r_cell_wire[808];							inform_R[852][7] = r_cell_wire[809];							inform_R[789][7] = r_cell_wire[810];							inform_R[853][7] = r_cell_wire[811];							inform_R[790][7] = r_cell_wire[812];							inform_R[854][7] = r_cell_wire[813];							inform_R[791][7] = r_cell_wire[814];							inform_R[855][7] = r_cell_wire[815];							inform_R[792][7] = r_cell_wire[816];							inform_R[856][7] = r_cell_wire[817];							inform_R[793][7] = r_cell_wire[818];							inform_R[857][7] = r_cell_wire[819];							inform_R[794][7] = r_cell_wire[820];							inform_R[858][7] = r_cell_wire[821];							inform_R[795][7] = r_cell_wire[822];							inform_R[859][7] = r_cell_wire[823];							inform_R[796][7] = r_cell_wire[824];							inform_R[860][7] = r_cell_wire[825];							inform_R[797][7] = r_cell_wire[826];							inform_R[861][7] = r_cell_wire[827];							inform_R[798][7] = r_cell_wire[828];							inform_R[862][7] = r_cell_wire[829];							inform_R[799][7] = r_cell_wire[830];							inform_R[863][7] = r_cell_wire[831];							inform_R[800][7] = r_cell_wire[832];							inform_R[864][7] = r_cell_wire[833];							inform_R[801][7] = r_cell_wire[834];							inform_R[865][7] = r_cell_wire[835];							inform_R[802][7] = r_cell_wire[836];							inform_R[866][7] = r_cell_wire[837];							inform_R[803][7] = r_cell_wire[838];							inform_R[867][7] = r_cell_wire[839];							inform_R[804][7] = r_cell_wire[840];							inform_R[868][7] = r_cell_wire[841];							inform_R[805][7] = r_cell_wire[842];							inform_R[869][7] = r_cell_wire[843];							inform_R[806][7] = r_cell_wire[844];							inform_R[870][7] = r_cell_wire[845];							inform_R[807][7] = r_cell_wire[846];							inform_R[871][7] = r_cell_wire[847];							inform_R[808][7] = r_cell_wire[848];							inform_R[872][7] = r_cell_wire[849];							inform_R[809][7] = r_cell_wire[850];							inform_R[873][7] = r_cell_wire[851];							inform_R[810][7] = r_cell_wire[852];							inform_R[874][7] = r_cell_wire[853];							inform_R[811][7] = r_cell_wire[854];							inform_R[875][7] = r_cell_wire[855];							inform_R[812][7] = r_cell_wire[856];							inform_R[876][7] = r_cell_wire[857];							inform_R[813][7] = r_cell_wire[858];							inform_R[877][7] = r_cell_wire[859];							inform_R[814][7] = r_cell_wire[860];							inform_R[878][7] = r_cell_wire[861];							inform_R[815][7] = r_cell_wire[862];							inform_R[879][7] = r_cell_wire[863];							inform_R[816][7] = r_cell_wire[864];							inform_R[880][7] = r_cell_wire[865];							inform_R[817][7] = r_cell_wire[866];							inform_R[881][7] = r_cell_wire[867];							inform_R[818][7] = r_cell_wire[868];							inform_R[882][7] = r_cell_wire[869];							inform_R[819][7] = r_cell_wire[870];							inform_R[883][7] = r_cell_wire[871];							inform_R[820][7] = r_cell_wire[872];							inform_R[884][7] = r_cell_wire[873];							inform_R[821][7] = r_cell_wire[874];							inform_R[885][7] = r_cell_wire[875];							inform_R[822][7] = r_cell_wire[876];							inform_R[886][7] = r_cell_wire[877];							inform_R[823][7] = r_cell_wire[878];							inform_R[887][7] = r_cell_wire[879];							inform_R[824][7] = r_cell_wire[880];							inform_R[888][7] = r_cell_wire[881];							inform_R[825][7] = r_cell_wire[882];							inform_R[889][7] = r_cell_wire[883];							inform_R[826][7] = r_cell_wire[884];							inform_R[890][7] = r_cell_wire[885];							inform_R[827][7] = r_cell_wire[886];							inform_R[891][7] = r_cell_wire[887];							inform_R[828][7] = r_cell_wire[888];							inform_R[892][7] = r_cell_wire[889];							inform_R[829][7] = r_cell_wire[890];							inform_R[893][7] = r_cell_wire[891];							inform_R[830][7] = r_cell_wire[892];							inform_R[894][7] = r_cell_wire[893];							inform_R[831][7] = r_cell_wire[894];							inform_R[895][7] = r_cell_wire[895];							inform_R[896][7] = r_cell_wire[896];							inform_R[960][7] = r_cell_wire[897];							inform_R[897][7] = r_cell_wire[898];							inform_R[961][7] = r_cell_wire[899];							inform_R[898][7] = r_cell_wire[900];							inform_R[962][7] = r_cell_wire[901];							inform_R[899][7] = r_cell_wire[902];							inform_R[963][7] = r_cell_wire[903];							inform_R[900][7] = r_cell_wire[904];							inform_R[964][7] = r_cell_wire[905];							inform_R[901][7] = r_cell_wire[906];							inform_R[965][7] = r_cell_wire[907];							inform_R[902][7] = r_cell_wire[908];							inform_R[966][7] = r_cell_wire[909];							inform_R[903][7] = r_cell_wire[910];							inform_R[967][7] = r_cell_wire[911];							inform_R[904][7] = r_cell_wire[912];							inform_R[968][7] = r_cell_wire[913];							inform_R[905][7] = r_cell_wire[914];							inform_R[969][7] = r_cell_wire[915];							inform_R[906][7] = r_cell_wire[916];							inform_R[970][7] = r_cell_wire[917];							inform_R[907][7] = r_cell_wire[918];							inform_R[971][7] = r_cell_wire[919];							inform_R[908][7] = r_cell_wire[920];							inform_R[972][7] = r_cell_wire[921];							inform_R[909][7] = r_cell_wire[922];							inform_R[973][7] = r_cell_wire[923];							inform_R[910][7] = r_cell_wire[924];							inform_R[974][7] = r_cell_wire[925];							inform_R[911][7] = r_cell_wire[926];							inform_R[975][7] = r_cell_wire[927];							inform_R[912][7] = r_cell_wire[928];							inform_R[976][7] = r_cell_wire[929];							inform_R[913][7] = r_cell_wire[930];							inform_R[977][7] = r_cell_wire[931];							inform_R[914][7] = r_cell_wire[932];							inform_R[978][7] = r_cell_wire[933];							inform_R[915][7] = r_cell_wire[934];							inform_R[979][7] = r_cell_wire[935];							inform_R[916][7] = r_cell_wire[936];							inform_R[980][7] = r_cell_wire[937];							inform_R[917][7] = r_cell_wire[938];							inform_R[981][7] = r_cell_wire[939];							inform_R[918][7] = r_cell_wire[940];							inform_R[982][7] = r_cell_wire[941];							inform_R[919][7] = r_cell_wire[942];							inform_R[983][7] = r_cell_wire[943];							inform_R[920][7] = r_cell_wire[944];							inform_R[984][7] = r_cell_wire[945];							inform_R[921][7] = r_cell_wire[946];							inform_R[985][7] = r_cell_wire[947];							inform_R[922][7] = r_cell_wire[948];							inform_R[986][7] = r_cell_wire[949];							inform_R[923][7] = r_cell_wire[950];							inform_R[987][7] = r_cell_wire[951];							inform_R[924][7] = r_cell_wire[952];							inform_R[988][7] = r_cell_wire[953];							inform_R[925][7] = r_cell_wire[954];							inform_R[989][7] = r_cell_wire[955];							inform_R[926][7] = r_cell_wire[956];							inform_R[990][7] = r_cell_wire[957];							inform_R[927][7] = r_cell_wire[958];							inform_R[991][7] = r_cell_wire[959];							inform_R[928][7] = r_cell_wire[960];							inform_R[992][7] = r_cell_wire[961];							inform_R[929][7] = r_cell_wire[962];							inform_R[993][7] = r_cell_wire[963];							inform_R[930][7] = r_cell_wire[964];							inform_R[994][7] = r_cell_wire[965];							inform_R[931][7] = r_cell_wire[966];							inform_R[995][7] = r_cell_wire[967];							inform_R[932][7] = r_cell_wire[968];							inform_R[996][7] = r_cell_wire[969];							inform_R[933][7] = r_cell_wire[970];							inform_R[997][7] = r_cell_wire[971];							inform_R[934][7] = r_cell_wire[972];							inform_R[998][7] = r_cell_wire[973];							inform_R[935][7] = r_cell_wire[974];							inform_R[999][7] = r_cell_wire[975];							inform_R[936][7] = r_cell_wire[976];							inform_R[1000][7] = r_cell_wire[977];							inform_R[937][7] = r_cell_wire[978];							inform_R[1001][7] = r_cell_wire[979];							inform_R[938][7] = r_cell_wire[980];							inform_R[1002][7] = r_cell_wire[981];							inform_R[939][7] = r_cell_wire[982];							inform_R[1003][7] = r_cell_wire[983];							inform_R[940][7] = r_cell_wire[984];							inform_R[1004][7] = r_cell_wire[985];							inform_R[941][7] = r_cell_wire[986];							inform_R[1005][7] = r_cell_wire[987];							inform_R[942][7] = r_cell_wire[988];							inform_R[1006][7] = r_cell_wire[989];							inform_R[943][7] = r_cell_wire[990];							inform_R[1007][7] = r_cell_wire[991];							inform_R[944][7] = r_cell_wire[992];							inform_R[1008][7] = r_cell_wire[993];							inform_R[945][7] = r_cell_wire[994];							inform_R[1009][7] = r_cell_wire[995];							inform_R[946][7] = r_cell_wire[996];							inform_R[1010][7] = r_cell_wire[997];							inform_R[947][7] = r_cell_wire[998];							inform_R[1011][7] = r_cell_wire[999];							inform_R[948][7] = r_cell_wire[1000];							inform_R[1012][7] = r_cell_wire[1001];							inform_R[949][7] = r_cell_wire[1002];							inform_R[1013][7] = r_cell_wire[1003];							inform_R[950][7] = r_cell_wire[1004];							inform_R[1014][7] = r_cell_wire[1005];							inform_R[951][7] = r_cell_wire[1006];							inform_R[1015][7] = r_cell_wire[1007];							inform_R[952][7] = r_cell_wire[1008];							inform_R[1016][7] = r_cell_wire[1009];							inform_R[953][7] = r_cell_wire[1010];							inform_R[1017][7] = r_cell_wire[1011];							inform_R[954][7] = r_cell_wire[1012];							inform_R[1018][7] = r_cell_wire[1013];							inform_R[955][7] = r_cell_wire[1014];							inform_R[1019][7] = r_cell_wire[1015];							inform_R[956][7] = r_cell_wire[1016];							inform_R[1020][7] = r_cell_wire[1017];							inform_R[957][7] = r_cell_wire[1018];							inform_R[1021][7] = r_cell_wire[1019];							inform_R[958][7] = r_cell_wire[1020];							inform_R[1022][7] = r_cell_wire[1021];							inform_R[959][7] = r_cell_wire[1022];							inform_R[1023][7] = r_cell_wire[1023];							inform_L[0][6] = l_cell_wire[0];							inform_L[64][6] = l_cell_wire[1];							inform_L[1][6] = l_cell_wire[2];							inform_L[65][6] = l_cell_wire[3];							inform_L[2][6] = l_cell_wire[4];							inform_L[66][6] = l_cell_wire[5];							inform_L[3][6] = l_cell_wire[6];							inform_L[67][6] = l_cell_wire[7];							inform_L[4][6] = l_cell_wire[8];							inform_L[68][6] = l_cell_wire[9];							inform_L[5][6] = l_cell_wire[10];							inform_L[69][6] = l_cell_wire[11];							inform_L[6][6] = l_cell_wire[12];							inform_L[70][6] = l_cell_wire[13];							inform_L[7][6] = l_cell_wire[14];							inform_L[71][6] = l_cell_wire[15];							inform_L[8][6] = l_cell_wire[16];							inform_L[72][6] = l_cell_wire[17];							inform_L[9][6] = l_cell_wire[18];							inform_L[73][6] = l_cell_wire[19];							inform_L[10][6] = l_cell_wire[20];							inform_L[74][6] = l_cell_wire[21];							inform_L[11][6] = l_cell_wire[22];							inform_L[75][6] = l_cell_wire[23];							inform_L[12][6] = l_cell_wire[24];							inform_L[76][6] = l_cell_wire[25];							inform_L[13][6] = l_cell_wire[26];							inform_L[77][6] = l_cell_wire[27];							inform_L[14][6] = l_cell_wire[28];							inform_L[78][6] = l_cell_wire[29];							inform_L[15][6] = l_cell_wire[30];							inform_L[79][6] = l_cell_wire[31];							inform_L[16][6] = l_cell_wire[32];							inform_L[80][6] = l_cell_wire[33];							inform_L[17][6] = l_cell_wire[34];							inform_L[81][6] = l_cell_wire[35];							inform_L[18][6] = l_cell_wire[36];							inform_L[82][6] = l_cell_wire[37];							inform_L[19][6] = l_cell_wire[38];							inform_L[83][6] = l_cell_wire[39];							inform_L[20][6] = l_cell_wire[40];							inform_L[84][6] = l_cell_wire[41];							inform_L[21][6] = l_cell_wire[42];							inform_L[85][6] = l_cell_wire[43];							inform_L[22][6] = l_cell_wire[44];							inform_L[86][6] = l_cell_wire[45];							inform_L[23][6] = l_cell_wire[46];							inform_L[87][6] = l_cell_wire[47];							inform_L[24][6] = l_cell_wire[48];							inform_L[88][6] = l_cell_wire[49];							inform_L[25][6] = l_cell_wire[50];							inform_L[89][6] = l_cell_wire[51];							inform_L[26][6] = l_cell_wire[52];							inform_L[90][6] = l_cell_wire[53];							inform_L[27][6] = l_cell_wire[54];							inform_L[91][6] = l_cell_wire[55];							inform_L[28][6] = l_cell_wire[56];							inform_L[92][6] = l_cell_wire[57];							inform_L[29][6] = l_cell_wire[58];							inform_L[93][6] = l_cell_wire[59];							inform_L[30][6] = l_cell_wire[60];							inform_L[94][6] = l_cell_wire[61];							inform_L[31][6] = l_cell_wire[62];							inform_L[95][6] = l_cell_wire[63];							inform_L[32][6] = l_cell_wire[64];							inform_L[96][6] = l_cell_wire[65];							inform_L[33][6] = l_cell_wire[66];							inform_L[97][6] = l_cell_wire[67];							inform_L[34][6] = l_cell_wire[68];							inform_L[98][6] = l_cell_wire[69];							inform_L[35][6] = l_cell_wire[70];							inform_L[99][6] = l_cell_wire[71];							inform_L[36][6] = l_cell_wire[72];							inform_L[100][6] = l_cell_wire[73];							inform_L[37][6] = l_cell_wire[74];							inform_L[101][6] = l_cell_wire[75];							inform_L[38][6] = l_cell_wire[76];							inform_L[102][6] = l_cell_wire[77];							inform_L[39][6] = l_cell_wire[78];							inform_L[103][6] = l_cell_wire[79];							inform_L[40][6] = l_cell_wire[80];							inform_L[104][6] = l_cell_wire[81];							inform_L[41][6] = l_cell_wire[82];							inform_L[105][6] = l_cell_wire[83];							inform_L[42][6] = l_cell_wire[84];							inform_L[106][6] = l_cell_wire[85];							inform_L[43][6] = l_cell_wire[86];							inform_L[107][6] = l_cell_wire[87];							inform_L[44][6] = l_cell_wire[88];							inform_L[108][6] = l_cell_wire[89];							inform_L[45][6] = l_cell_wire[90];							inform_L[109][6] = l_cell_wire[91];							inform_L[46][6] = l_cell_wire[92];							inform_L[110][6] = l_cell_wire[93];							inform_L[47][6] = l_cell_wire[94];							inform_L[111][6] = l_cell_wire[95];							inform_L[48][6] = l_cell_wire[96];							inform_L[112][6] = l_cell_wire[97];							inform_L[49][6] = l_cell_wire[98];							inform_L[113][6] = l_cell_wire[99];							inform_L[50][6] = l_cell_wire[100];							inform_L[114][6] = l_cell_wire[101];							inform_L[51][6] = l_cell_wire[102];							inform_L[115][6] = l_cell_wire[103];							inform_L[52][6] = l_cell_wire[104];							inform_L[116][6] = l_cell_wire[105];							inform_L[53][6] = l_cell_wire[106];							inform_L[117][6] = l_cell_wire[107];							inform_L[54][6] = l_cell_wire[108];							inform_L[118][6] = l_cell_wire[109];							inform_L[55][6] = l_cell_wire[110];							inform_L[119][6] = l_cell_wire[111];							inform_L[56][6] = l_cell_wire[112];							inform_L[120][6] = l_cell_wire[113];							inform_L[57][6] = l_cell_wire[114];							inform_L[121][6] = l_cell_wire[115];							inform_L[58][6] = l_cell_wire[116];							inform_L[122][6] = l_cell_wire[117];							inform_L[59][6] = l_cell_wire[118];							inform_L[123][6] = l_cell_wire[119];							inform_L[60][6] = l_cell_wire[120];							inform_L[124][6] = l_cell_wire[121];							inform_L[61][6] = l_cell_wire[122];							inform_L[125][6] = l_cell_wire[123];							inform_L[62][6] = l_cell_wire[124];							inform_L[126][6] = l_cell_wire[125];							inform_L[63][6] = l_cell_wire[126];							inform_L[127][6] = l_cell_wire[127];							inform_L[128][6] = l_cell_wire[128];							inform_L[192][6] = l_cell_wire[129];							inform_L[129][6] = l_cell_wire[130];							inform_L[193][6] = l_cell_wire[131];							inform_L[130][6] = l_cell_wire[132];							inform_L[194][6] = l_cell_wire[133];							inform_L[131][6] = l_cell_wire[134];							inform_L[195][6] = l_cell_wire[135];							inform_L[132][6] = l_cell_wire[136];							inform_L[196][6] = l_cell_wire[137];							inform_L[133][6] = l_cell_wire[138];							inform_L[197][6] = l_cell_wire[139];							inform_L[134][6] = l_cell_wire[140];							inform_L[198][6] = l_cell_wire[141];							inform_L[135][6] = l_cell_wire[142];							inform_L[199][6] = l_cell_wire[143];							inform_L[136][6] = l_cell_wire[144];							inform_L[200][6] = l_cell_wire[145];							inform_L[137][6] = l_cell_wire[146];							inform_L[201][6] = l_cell_wire[147];							inform_L[138][6] = l_cell_wire[148];							inform_L[202][6] = l_cell_wire[149];							inform_L[139][6] = l_cell_wire[150];							inform_L[203][6] = l_cell_wire[151];							inform_L[140][6] = l_cell_wire[152];							inform_L[204][6] = l_cell_wire[153];							inform_L[141][6] = l_cell_wire[154];							inform_L[205][6] = l_cell_wire[155];							inform_L[142][6] = l_cell_wire[156];							inform_L[206][6] = l_cell_wire[157];							inform_L[143][6] = l_cell_wire[158];							inform_L[207][6] = l_cell_wire[159];							inform_L[144][6] = l_cell_wire[160];							inform_L[208][6] = l_cell_wire[161];							inform_L[145][6] = l_cell_wire[162];							inform_L[209][6] = l_cell_wire[163];							inform_L[146][6] = l_cell_wire[164];							inform_L[210][6] = l_cell_wire[165];							inform_L[147][6] = l_cell_wire[166];							inform_L[211][6] = l_cell_wire[167];							inform_L[148][6] = l_cell_wire[168];							inform_L[212][6] = l_cell_wire[169];							inform_L[149][6] = l_cell_wire[170];							inform_L[213][6] = l_cell_wire[171];							inform_L[150][6] = l_cell_wire[172];							inform_L[214][6] = l_cell_wire[173];							inform_L[151][6] = l_cell_wire[174];							inform_L[215][6] = l_cell_wire[175];							inform_L[152][6] = l_cell_wire[176];							inform_L[216][6] = l_cell_wire[177];							inform_L[153][6] = l_cell_wire[178];							inform_L[217][6] = l_cell_wire[179];							inform_L[154][6] = l_cell_wire[180];							inform_L[218][6] = l_cell_wire[181];							inform_L[155][6] = l_cell_wire[182];							inform_L[219][6] = l_cell_wire[183];							inform_L[156][6] = l_cell_wire[184];							inform_L[220][6] = l_cell_wire[185];							inform_L[157][6] = l_cell_wire[186];							inform_L[221][6] = l_cell_wire[187];							inform_L[158][6] = l_cell_wire[188];							inform_L[222][6] = l_cell_wire[189];							inform_L[159][6] = l_cell_wire[190];							inform_L[223][6] = l_cell_wire[191];							inform_L[160][6] = l_cell_wire[192];							inform_L[224][6] = l_cell_wire[193];							inform_L[161][6] = l_cell_wire[194];							inform_L[225][6] = l_cell_wire[195];							inform_L[162][6] = l_cell_wire[196];							inform_L[226][6] = l_cell_wire[197];							inform_L[163][6] = l_cell_wire[198];							inform_L[227][6] = l_cell_wire[199];							inform_L[164][6] = l_cell_wire[200];							inform_L[228][6] = l_cell_wire[201];							inform_L[165][6] = l_cell_wire[202];							inform_L[229][6] = l_cell_wire[203];							inform_L[166][6] = l_cell_wire[204];							inform_L[230][6] = l_cell_wire[205];							inform_L[167][6] = l_cell_wire[206];							inform_L[231][6] = l_cell_wire[207];							inform_L[168][6] = l_cell_wire[208];							inform_L[232][6] = l_cell_wire[209];							inform_L[169][6] = l_cell_wire[210];							inform_L[233][6] = l_cell_wire[211];							inform_L[170][6] = l_cell_wire[212];							inform_L[234][6] = l_cell_wire[213];							inform_L[171][6] = l_cell_wire[214];							inform_L[235][6] = l_cell_wire[215];							inform_L[172][6] = l_cell_wire[216];							inform_L[236][6] = l_cell_wire[217];							inform_L[173][6] = l_cell_wire[218];							inform_L[237][6] = l_cell_wire[219];							inform_L[174][6] = l_cell_wire[220];							inform_L[238][6] = l_cell_wire[221];							inform_L[175][6] = l_cell_wire[222];							inform_L[239][6] = l_cell_wire[223];							inform_L[176][6] = l_cell_wire[224];							inform_L[240][6] = l_cell_wire[225];							inform_L[177][6] = l_cell_wire[226];							inform_L[241][6] = l_cell_wire[227];							inform_L[178][6] = l_cell_wire[228];							inform_L[242][6] = l_cell_wire[229];							inform_L[179][6] = l_cell_wire[230];							inform_L[243][6] = l_cell_wire[231];							inform_L[180][6] = l_cell_wire[232];							inform_L[244][6] = l_cell_wire[233];							inform_L[181][6] = l_cell_wire[234];							inform_L[245][6] = l_cell_wire[235];							inform_L[182][6] = l_cell_wire[236];							inform_L[246][6] = l_cell_wire[237];							inform_L[183][6] = l_cell_wire[238];							inform_L[247][6] = l_cell_wire[239];							inform_L[184][6] = l_cell_wire[240];							inform_L[248][6] = l_cell_wire[241];							inform_L[185][6] = l_cell_wire[242];							inform_L[249][6] = l_cell_wire[243];							inform_L[186][6] = l_cell_wire[244];							inform_L[250][6] = l_cell_wire[245];							inform_L[187][6] = l_cell_wire[246];							inform_L[251][6] = l_cell_wire[247];							inform_L[188][6] = l_cell_wire[248];							inform_L[252][6] = l_cell_wire[249];							inform_L[189][6] = l_cell_wire[250];							inform_L[253][6] = l_cell_wire[251];							inform_L[190][6] = l_cell_wire[252];							inform_L[254][6] = l_cell_wire[253];							inform_L[191][6] = l_cell_wire[254];							inform_L[255][6] = l_cell_wire[255];							inform_L[256][6] = l_cell_wire[256];							inform_L[320][6] = l_cell_wire[257];							inform_L[257][6] = l_cell_wire[258];							inform_L[321][6] = l_cell_wire[259];							inform_L[258][6] = l_cell_wire[260];							inform_L[322][6] = l_cell_wire[261];							inform_L[259][6] = l_cell_wire[262];							inform_L[323][6] = l_cell_wire[263];							inform_L[260][6] = l_cell_wire[264];							inform_L[324][6] = l_cell_wire[265];							inform_L[261][6] = l_cell_wire[266];							inform_L[325][6] = l_cell_wire[267];							inform_L[262][6] = l_cell_wire[268];							inform_L[326][6] = l_cell_wire[269];							inform_L[263][6] = l_cell_wire[270];							inform_L[327][6] = l_cell_wire[271];							inform_L[264][6] = l_cell_wire[272];							inform_L[328][6] = l_cell_wire[273];							inform_L[265][6] = l_cell_wire[274];							inform_L[329][6] = l_cell_wire[275];							inform_L[266][6] = l_cell_wire[276];							inform_L[330][6] = l_cell_wire[277];							inform_L[267][6] = l_cell_wire[278];							inform_L[331][6] = l_cell_wire[279];							inform_L[268][6] = l_cell_wire[280];							inform_L[332][6] = l_cell_wire[281];							inform_L[269][6] = l_cell_wire[282];							inform_L[333][6] = l_cell_wire[283];							inform_L[270][6] = l_cell_wire[284];							inform_L[334][6] = l_cell_wire[285];							inform_L[271][6] = l_cell_wire[286];							inform_L[335][6] = l_cell_wire[287];							inform_L[272][6] = l_cell_wire[288];							inform_L[336][6] = l_cell_wire[289];							inform_L[273][6] = l_cell_wire[290];							inform_L[337][6] = l_cell_wire[291];							inform_L[274][6] = l_cell_wire[292];							inform_L[338][6] = l_cell_wire[293];							inform_L[275][6] = l_cell_wire[294];							inform_L[339][6] = l_cell_wire[295];							inform_L[276][6] = l_cell_wire[296];							inform_L[340][6] = l_cell_wire[297];							inform_L[277][6] = l_cell_wire[298];							inform_L[341][6] = l_cell_wire[299];							inform_L[278][6] = l_cell_wire[300];							inform_L[342][6] = l_cell_wire[301];							inform_L[279][6] = l_cell_wire[302];							inform_L[343][6] = l_cell_wire[303];							inform_L[280][6] = l_cell_wire[304];							inform_L[344][6] = l_cell_wire[305];							inform_L[281][6] = l_cell_wire[306];							inform_L[345][6] = l_cell_wire[307];							inform_L[282][6] = l_cell_wire[308];							inform_L[346][6] = l_cell_wire[309];							inform_L[283][6] = l_cell_wire[310];							inform_L[347][6] = l_cell_wire[311];							inform_L[284][6] = l_cell_wire[312];							inform_L[348][6] = l_cell_wire[313];							inform_L[285][6] = l_cell_wire[314];							inform_L[349][6] = l_cell_wire[315];							inform_L[286][6] = l_cell_wire[316];							inform_L[350][6] = l_cell_wire[317];							inform_L[287][6] = l_cell_wire[318];							inform_L[351][6] = l_cell_wire[319];							inform_L[288][6] = l_cell_wire[320];							inform_L[352][6] = l_cell_wire[321];							inform_L[289][6] = l_cell_wire[322];							inform_L[353][6] = l_cell_wire[323];							inform_L[290][6] = l_cell_wire[324];							inform_L[354][6] = l_cell_wire[325];							inform_L[291][6] = l_cell_wire[326];							inform_L[355][6] = l_cell_wire[327];							inform_L[292][6] = l_cell_wire[328];							inform_L[356][6] = l_cell_wire[329];							inform_L[293][6] = l_cell_wire[330];							inform_L[357][6] = l_cell_wire[331];							inform_L[294][6] = l_cell_wire[332];							inform_L[358][6] = l_cell_wire[333];							inform_L[295][6] = l_cell_wire[334];							inform_L[359][6] = l_cell_wire[335];							inform_L[296][6] = l_cell_wire[336];							inform_L[360][6] = l_cell_wire[337];							inform_L[297][6] = l_cell_wire[338];							inform_L[361][6] = l_cell_wire[339];							inform_L[298][6] = l_cell_wire[340];							inform_L[362][6] = l_cell_wire[341];							inform_L[299][6] = l_cell_wire[342];							inform_L[363][6] = l_cell_wire[343];							inform_L[300][6] = l_cell_wire[344];							inform_L[364][6] = l_cell_wire[345];							inform_L[301][6] = l_cell_wire[346];							inform_L[365][6] = l_cell_wire[347];							inform_L[302][6] = l_cell_wire[348];							inform_L[366][6] = l_cell_wire[349];							inform_L[303][6] = l_cell_wire[350];							inform_L[367][6] = l_cell_wire[351];							inform_L[304][6] = l_cell_wire[352];							inform_L[368][6] = l_cell_wire[353];							inform_L[305][6] = l_cell_wire[354];							inform_L[369][6] = l_cell_wire[355];							inform_L[306][6] = l_cell_wire[356];							inform_L[370][6] = l_cell_wire[357];							inform_L[307][6] = l_cell_wire[358];							inform_L[371][6] = l_cell_wire[359];							inform_L[308][6] = l_cell_wire[360];							inform_L[372][6] = l_cell_wire[361];							inform_L[309][6] = l_cell_wire[362];							inform_L[373][6] = l_cell_wire[363];							inform_L[310][6] = l_cell_wire[364];							inform_L[374][6] = l_cell_wire[365];							inform_L[311][6] = l_cell_wire[366];							inform_L[375][6] = l_cell_wire[367];							inform_L[312][6] = l_cell_wire[368];							inform_L[376][6] = l_cell_wire[369];							inform_L[313][6] = l_cell_wire[370];							inform_L[377][6] = l_cell_wire[371];							inform_L[314][6] = l_cell_wire[372];							inform_L[378][6] = l_cell_wire[373];							inform_L[315][6] = l_cell_wire[374];							inform_L[379][6] = l_cell_wire[375];							inform_L[316][6] = l_cell_wire[376];							inform_L[380][6] = l_cell_wire[377];							inform_L[317][6] = l_cell_wire[378];							inform_L[381][6] = l_cell_wire[379];							inform_L[318][6] = l_cell_wire[380];							inform_L[382][6] = l_cell_wire[381];							inform_L[319][6] = l_cell_wire[382];							inform_L[383][6] = l_cell_wire[383];							inform_L[384][6] = l_cell_wire[384];							inform_L[448][6] = l_cell_wire[385];							inform_L[385][6] = l_cell_wire[386];							inform_L[449][6] = l_cell_wire[387];							inform_L[386][6] = l_cell_wire[388];							inform_L[450][6] = l_cell_wire[389];							inform_L[387][6] = l_cell_wire[390];							inform_L[451][6] = l_cell_wire[391];							inform_L[388][6] = l_cell_wire[392];							inform_L[452][6] = l_cell_wire[393];							inform_L[389][6] = l_cell_wire[394];							inform_L[453][6] = l_cell_wire[395];							inform_L[390][6] = l_cell_wire[396];							inform_L[454][6] = l_cell_wire[397];							inform_L[391][6] = l_cell_wire[398];							inform_L[455][6] = l_cell_wire[399];							inform_L[392][6] = l_cell_wire[400];							inform_L[456][6] = l_cell_wire[401];							inform_L[393][6] = l_cell_wire[402];							inform_L[457][6] = l_cell_wire[403];							inform_L[394][6] = l_cell_wire[404];							inform_L[458][6] = l_cell_wire[405];							inform_L[395][6] = l_cell_wire[406];							inform_L[459][6] = l_cell_wire[407];							inform_L[396][6] = l_cell_wire[408];							inform_L[460][6] = l_cell_wire[409];							inform_L[397][6] = l_cell_wire[410];							inform_L[461][6] = l_cell_wire[411];							inform_L[398][6] = l_cell_wire[412];							inform_L[462][6] = l_cell_wire[413];							inform_L[399][6] = l_cell_wire[414];							inform_L[463][6] = l_cell_wire[415];							inform_L[400][6] = l_cell_wire[416];							inform_L[464][6] = l_cell_wire[417];							inform_L[401][6] = l_cell_wire[418];							inform_L[465][6] = l_cell_wire[419];							inform_L[402][6] = l_cell_wire[420];							inform_L[466][6] = l_cell_wire[421];							inform_L[403][6] = l_cell_wire[422];							inform_L[467][6] = l_cell_wire[423];							inform_L[404][6] = l_cell_wire[424];							inform_L[468][6] = l_cell_wire[425];							inform_L[405][6] = l_cell_wire[426];							inform_L[469][6] = l_cell_wire[427];							inform_L[406][6] = l_cell_wire[428];							inform_L[470][6] = l_cell_wire[429];							inform_L[407][6] = l_cell_wire[430];							inform_L[471][6] = l_cell_wire[431];							inform_L[408][6] = l_cell_wire[432];							inform_L[472][6] = l_cell_wire[433];							inform_L[409][6] = l_cell_wire[434];							inform_L[473][6] = l_cell_wire[435];							inform_L[410][6] = l_cell_wire[436];							inform_L[474][6] = l_cell_wire[437];							inform_L[411][6] = l_cell_wire[438];							inform_L[475][6] = l_cell_wire[439];							inform_L[412][6] = l_cell_wire[440];							inform_L[476][6] = l_cell_wire[441];							inform_L[413][6] = l_cell_wire[442];							inform_L[477][6] = l_cell_wire[443];							inform_L[414][6] = l_cell_wire[444];							inform_L[478][6] = l_cell_wire[445];							inform_L[415][6] = l_cell_wire[446];							inform_L[479][6] = l_cell_wire[447];							inform_L[416][6] = l_cell_wire[448];							inform_L[480][6] = l_cell_wire[449];							inform_L[417][6] = l_cell_wire[450];							inform_L[481][6] = l_cell_wire[451];							inform_L[418][6] = l_cell_wire[452];							inform_L[482][6] = l_cell_wire[453];							inform_L[419][6] = l_cell_wire[454];							inform_L[483][6] = l_cell_wire[455];							inform_L[420][6] = l_cell_wire[456];							inform_L[484][6] = l_cell_wire[457];							inform_L[421][6] = l_cell_wire[458];							inform_L[485][6] = l_cell_wire[459];							inform_L[422][6] = l_cell_wire[460];							inform_L[486][6] = l_cell_wire[461];							inform_L[423][6] = l_cell_wire[462];							inform_L[487][6] = l_cell_wire[463];							inform_L[424][6] = l_cell_wire[464];							inform_L[488][6] = l_cell_wire[465];							inform_L[425][6] = l_cell_wire[466];							inform_L[489][6] = l_cell_wire[467];							inform_L[426][6] = l_cell_wire[468];							inform_L[490][6] = l_cell_wire[469];							inform_L[427][6] = l_cell_wire[470];							inform_L[491][6] = l_cell_wire[471];							inform_L[428][6] = l_cell_wire[472];							inform_L[492][6] = l_cell_wire[473];							inform_L[429][6] = l_cell_wire[474];							inform_L[493][6] = l_cell_wire[475];							inform_L[430][6] = l_cell_wire[476];							inform_L[494][6] = l_cell_wire[477];							inform_L[431][6] = l_cell_wire[478];							inform_L[495][6] = l_cell_wire[479];							inform_L[432][6] = l_cell_wire[480];							inform_L[496][6] = l_cell_wire[481];							inform_L[433][6] = l_cell_wire[482];							inform_L[497][6] = l_cell_wire[483];							inform_L[434][6] = l_cell_wire[484];							inform_L[498][6] = l_cell_wire[485];							inform_L[435][6] = l_cell_wire[486];							inform_L[499][6] = l_cell_wire[487];							inform_L[436][6] = l_cell_wire[488];							inform_L[500][6] = l_cell_wire[489];							inform_L[437][6] = l_cell_wire[490];							inform_L[501][6] = l_cell_wire[491];							inform_L[438][6] = l_cell_wire[492];							inform_L[502][6] = l_cell_wire[493];							inform_L[439][6] = l_cell_wire[494];							inform_L[503][6] = l_cell_wire[495];							inform_L[440][6] = l_cell_wire[496];							inform_L[504][6] = l_cell_wire[497];							inform_L[441][6] = l_cell_wire[498];							inform_L[505][6] = l_cell_wire[499];							inform_L[442][6] = l_cell_wire[500];							inform_L[506][6] = l_cell_wire[501];							inform_L[443][6] = l_cell_wire[502];							inform_L[507][6] = l_cell_wire[503];							inform_L[444][6] = l_cell_wire[504];							inform_L[508][6] = l_cell_wire[505];							inform_L[445][6] = l_cell_wire[506];							inform_L[509][6] = l_cell_wire[507];							inform_L[446][6] = l_cell_wire[508];							inform_L[510][6] = l_cell_wire[509];							inform_L[447][6] = l_cell_wire[510];							inform_L[511][6] = l_cell_wire[511];							inform_L[512][6] = l_cell_wire[512];							inform_L[576][6] = l_cell_wire[513];							inform_L[513][6] = l_cell_wire[514];							inform_L[577][6] = l_cell_wire[515];							inform_L[514][6] = l_cell_wire[516];							inform_L[578][6] = l_cell_wire[517];							inform_L[515][6] = l_cell_wire[518];							inform_L[579][6] = l_cell_wire[519];							inform_L[516][6] = l_cell_wire[520];							inform_L[580][6] = l_cell_wire[521];							inform_L[517][6] = l_cell_wire[522];							inform_L[581][6] = l_cell_wire[523];							inform_L[518][6] = l_cell_wire[524];							inform_L[582][6] = l_cell_wire[525];							inform_L[519][6] = l_cell_wire[526];							inform_L[583][6] = l_cell_wire[527];							inform_L[520][6] = l_cell_wire[528];							inform_L[584][6] = l_cell_wire[529];							inform_L[521][6] = l_cell_wire[530];							inform_L[585][6] = l_cell_wire[531];							inform_L[522][6] = l_cell_wire[532];							inform_L[586][6] = l_cell_wire[533];							inform_L[523][6] = l_cell_wire[534];							inform_L[587][6] = l_cell_wire[535];							inform_L[524][6] = l_cell_wire[536];							inform_L[588][6] = l_cell_wire[537];							inform_L[525][6] = l_cell_wire[538];							inform_L[589][6] = l_cell_wire[539];							inform_L[526][6] = l_cell_wire[540];							inform_L[590][6] = l_cell_wire[541];							inform_L[527][6] = l_cell_wire[542];							inform_L[591][6] = l_cell_wire[543];							inform_L[528][6] = l_cell_wire[544];							inform_L[592][6] = l_cell_wire[545];							inform_L[529][6] = l_cell_wire[546];							inform_L[593][6] = l_cell_wire[547];							inform_L[530][6] = l_cell_wire[548];							inform_L[594][6] = l_cell_wire[549];							inform_L[531][6] = l_cell_wire[550];							inform_L[595][6] = l_cell_wire[551];							inform_L[532][6] = l_cell_wire[552];							inform_L[596][6] = l_cell_wire[553];							inform_L[533][6] = l_cell_wire[554];							inform_L[597][6] = l_cell_wire[555];							inform_L[534][6] = l_cell_wire[556];							inform_L[598][6] = l_cell_wire[557];							inform_L[535][6] = l_cell_wire[558];							inform_L[599][6] = l_cell_wire[559];							inform_L[536][6] = l_cell_wire[560];							inform_L[600][6] = l_cell_wire[561];							inform_L[537][6] = l_cell_wire[562];							inform_L[601][6] = l_cell_wire[563];							inform_L[538][6] = l_cell_wire[564];							inform_L[602][6] = l_cell_wire[565];							inform_L[539][6] = l_cell_wire[566];							inform_L[603][6] = l_cell_wire[567];							inform_L[540][6] = l_cell_wire[568];							inform_L[604][6] = l_cell_wire[569];							inform_L[541][6] = l_cell_wire[570];							inform_L[605][6] = l_cell_wire[571];							inform_L[542][6] = l_cell_wire[572];							inform_L[606][6] = l_cell_wire[573];							inform_L[543][6] = l_cell_wire[574];							inform_L[607][6] = l_cell_wire[575];							inform_L[544][6] = l_cell_wire[576];							inform_L[608][6] = l_cell_wire[577];							inform_L[545][6] = l_cell_wire[578];							inform_L[609][6] = l_cell_wire[579];							inform_L[546][6] = l_cell_wire[580];							inform_L[610][6] = l_cell_wire[581];							inform_L[547][6] = l_cell_wire[582];							inform_L[611][6] = l_cell_wire[583];							inform_L[548][6] = l_cell_wire[584];							inform_L[612][6] = l_cell_wire[585];							inform_L[549][6] = l_cell_wire[586];							inform_L[613][6] = l_cell_wire[587];							inform_L[550][6] = l_cell_wire[588];							inform_L[614][6] = l_cell_wire[589];							inform_L[551][6] = l_cell_wire[590];							inform_L[615][6] = l_cell_wire[591];							inform_L[552][6] = l_cell_wire[592];							inform_L[616][6] = l_cell_wire[593];							inform_L[553][6] = l_cell_wire[594];							inform_L[617][6] = l_cell_wire[595];							inform_L[554][6] = l_cell_wire[596];							inform_L[618][6] = l_cell_wire[597];							inform_L[555][6] = l_cell_wire[598];							inform_L[619][6] = l_cell_wire[599];							inform_L[556][6] = l_cell_wire[600];							inform_L[620][6] = l_cell_wire[601];							inform_L[557][6] = l_cell_wire[602];							inform_L[621][6] = l_cell_wire[603];							inform_L[558][6] = l_cell_wire[604];							inform_L[622][6] = l_cell_wire[605];							inform_L[559][6] = l_cell_wire[606];							inform_L[623][6] = l_cell_wire[607];							inform_L[560][6] = l_cell_wire[608];							inform_L[624][6] = l_cell_wire[609];							inform_L[561][6] = l_cell_wire[610];							inform_L[625][6] = l_cell_wire[611];							inform_L[562][6] = l_cell_wire[612];							inform_L[626][6] = l_cell_wire[613];							inform_L[563][6] = l_cell_wire[614];							inform_L[627][6] = l_cell_wire[615];							inform_L[564][6] = l_cell_wire[616];							inform_L[628][6] = l_cell_wire[617];							inform_L[565][6] = l_cell_wire[618];							inform_L[629][6] = l_cell_wire[619];							inform_L[566][6] = l_cell_wire[620];							inform_L[630][6] = l_cell_wire[621];							inform_L[567][6] = l_cell_wire[622];							inform_L[631][6] = l_cell_wire[623];							inform_L[568][6] = l_cell_wire[624];							inform_L[632][6] = l_cell_wire[625];							inform_L[569][6] = l_cell_wire[626];							inform_L[633][6] = l_cell_wire[627];							inform_L[570][6] = l_cell_wire[628];							inform_L[634][6] = l_cell_wire[629];							inform_L[571][6] = l_cell_wire[630];							inform_L[635][6] = l_cell_wire[631];							inform_L[572][6] = l_cell_wire[632];							inform_L[636][6] = l_cell_wire[633];							inform_L[573][6] = l_cell_wire[634];							inform_L[637][6] = l_cell_wire[635];							inform_L[574][6] = l_cell_wire[636];							inform_L[638][6] = l_cell_wire[637];							inform_L[575][6] = l_cell_wire[638];							inform_L[639][6] = l_cell_wire[639];							inform_L[640][6] = l_cell_wire[640];							inform_L[704][6] = l_cell_wire[641];							inform_L[641][6] = l_cell_wire[642];							inform_L[705][6] = l_cell_wire[643];							inform_L[642][6] = l_cell_wire[644];							inform_L[706][6] = l_cell_wire[645];							inform_L[643][6] = l_cell_wire[646];							inform_L[707][6] = l_cell_wire[647];							inform_L[644][6] = l_cell_wire[648];							inform_L[708][6] = l_cell_wire[649];							inform_L[645][6] = l_cell_wire[650];							inform_L[709][6] = l_cell_wire[651];							inform_L[646][6] = l_cell_wire[652];							inform_L[710][6] = l_cell_wire[653];							inform_L[647][6] = l_cell_wire[654];							inform_L[711][6] = l_cell_wire[655];							inform_L[648][6] = l_cell_wire[656];							inform_L[712][6] = l_cell_wire[657];							inform_L[649][6] = l_cell_wire[658];							inform_L[713][6] = l_cell_wire[659];							inform_L[650][6] = l_cell_wire[660];							inform_L[714][6] = l_cell_wire[661];							inform_L[651][6] = l_cell_wire[662];							inform_L[715][6] = l_cell_wire[663];							inform_L[652][6] = l_cell_wire[664];							inform_L[716][6] = l_cell_wire[665];							inform_L[653][6] = l_cell_wire[666];							inform_L[717][6] = l_cell_wire[667];							inform_L[654][6] = l_cell_wire[668];							inform_L[718][6] = l_cell_wire[669];							inform_L[655][6] = l_cell_wire[670];							inform_L[719][6] = l_cell_wire[671];							inform_L[656][6] = l_cell_wire[672];							inform_L[720][6] = l_cell_wire[673];							inform_L[657][6] = l_cell_wire[674];							inform_L[721][6] = l_cell_wire[675];							inform_L[658][6] = l_cell_wire[676];							inform_L[722][6] = l_cell_wire[677];							inform_L[659][6] = l_cell_wire[678];							inform_L[723][6] = l_cell_wire[679];							inform_L[660][6] = l_cell_wire[680];							inform_L[724][6] = l_cell_wire[681];							inform_L[661][6] = l_cell_wire[682];							inform_L[725][6] = l_cell_wire[683];							inform_L[662][6] = l_cell_wire[684];							inform_L[726][6] = l_cell_wire[685];							inform_L[663][6] = l_cell_wire[686];							inform_L[727][6] = l_cell_wire[687];							inform_L[664][6] = l_cell_wire[688];							inform_L[728][6] = l_cell_wire[689];							inform_L[665][6] = l_cell_wire[690];							inform_L[729][6] = l_cell_wire[691];							inform_L[666][6] = l_cell_wire[692];							inform_L[730][6] = l_cell_wire[693];							inform_L[667][6] = l_cell_wire[694];							inform_L[731][6] = l_cell_wire[695];							inform_L[668][6] = l_cell_wire[696];							inform_L[732][6] = l_cell_wire[697];							inform_L[669][6] = l_cell_wire[698];							inform_L[733][6] = l_cell_wire[699];							inform_L[670][6] = l_cell_wire[700];							inform_L[734][6] = l_cell_wire[701];							inform_L[671][6] = l_cell_wire[702];							inform_L[735][6] = l_cell_wire[703];							inform_L[672][6] = l_cell_wire[704];							inform_L[736][6] = l_cell_wire[705];							inform_L[673][6] = l_cell_wire[706];							inform_L[737][6] = l_cell_wire[707];							inform_L[674][6] = l_cell_wire[708];							inform_L[738][6] = l_cell_wire[709];							inform_L[675][6] = l_cell_wire[710];							inform_L[739][6] = l_cell_wire[711];							inform_L[676][6] = l_cell_wire[712];							inform_L[740][6] = l_cell_wire[713];							inform_L[677][6] = l_cell_wire[714];							inform_L[741][6] = l_cell_wire[715];							inform_L[678][6] = l_cell_wire[716];							inform_L[742][6] = l_cell_wire[717];							inform_L[679][6] = l_cell_wire[718];							inform_L[743][6] = l_cell_wire[719];							inform_L[680][6] = l_cell_wire[720];							inform_L[744][6] = l_cell_wire[721];							inform_L[681][6] = l_cell_wire[722];							inform_L[745][6] = l_cell_wire[723];							inform_L[682][6] = l_cell_wire[724];							inform_L[746][6] = l_cell_wire[725];							inform_L[683][6] = l_cell_wire[726];							inform_L[747][6] = l_cell_wire[727];							inform_L[684][6] = l_cell_wire[728];							inform_L[748][6] = l_cell_wire[729];							inform_L[685][6] = l_cell_wire[730];							inform_L[749][6] = l_cell_wire[731];							inform_L[686][6] = l_cell_wire[732];							inform_L[750][6] = l_cell_wire[733];							inform_L[687][6] = l_cell_wire[734];							inform_L[751][6] = l_cell_wire[735];							inform_L[688][6] = l_cell_wire[736];							inform_L[752][6] = l_cell_wire[737];							inform_L[689][6] = l_cell_wire[738];							inform_L[753][6] = l_cell_wire[739];							inform_L[690][6] = l_cell_wire[740];							inform_L[754][6] = l_cell_wire[741];							inform_L[691][6] = l_cell_wire[742];							inform_L[755][6] = l_cell_wire[743];							inform_L[692][6] = l_cell_wire[744];							inform_L[756][6] = l_cell_wire[745];							inform_L[693][6] = l_cell_wire[746];							inform_L[757][6] = l_cell_wire[747];							inform_L[694][6] = l_cell_wire[748];							inform_L[758][6] = l_cell_wire[749];							inform_L[695][6] = l_cell_wire[750];							inform_L[759][6] = l_cell_wire[751];							inform_L[696][6] = l_cell_wire[752];							inform_L[760][6] = l_cell_wire[753];							inform_L[697][6] = l_cell_wire[754];							inform_L[761][6] = l_cell_wire[755];							inform_L[698][6] = l_cell_wire[756];							inform_L[762][6] = l_cell_wire[757];							inform_L[699][6] = l_cell_wire[758];							inform_L[763][6] = l_cell_wire[759];							inform_L[700][6] = l_cell_wire[760];							inform_L[764][6] = l_cell_wire[761];							inform_L[701][6] = l_cell_wire[762];							inform_L[765][6] = l_cell_wire[763];							inform_L[702][6] = l_cell_wire[764];							inform_L[766][6] = l_cell_wire[765];							inform_L[703][6] = l_cell_wire[766];							inform_L[767][6] = l_cell_wire[767];							inform_L[768][6] = l_cell_wire[768];							inform_L[832][6] = l_cell_wire[769];							inform_L[769][6] = l_cell_wire[770];							inform_L[833][6] = l_cell_wire[771];							inform_L[770][6] = l_cell_wire[772];							inform_L[834][6] = l_cell_wire[773];							inform_L[771][6] = l_cell_wire[774];							inform_L[835][6] = l_cell_wire[775];							inform_L[772][6] = l_cell_wire[776];							inform_L[836][6] = l_cell_wire[777];							inform_L[773][6] = l_cell_wire[778];							inform_L[837][6] = l_cell_wire[779];							inform_L[774][6] = l_cell_wire[780];							inform_L[838][6] = l_cell_wire[781];							inform_L[775][6] = l_cell_wire[782];							inform_L[839][6] = l_cell_wire[783];							inform_L[776][6] = l_cell_wire[784];							inform_L[840][6] = l_cell_wire[785];							inform_L[777][6] = l_cell_wire[786];							inform_L[841][6] = l_cell_wire[787];							inform_L[778][6] = l_cell_wire[788];							inform_L[842][6] = l_cell_wire[789];							inform_L[779][6] = l_cell_wire[790];							inform_L[843][6] = l_cell_wire[791];							inform_L[780][6] = l_cell_wire[792];							inform_L[844][6] = l_cell_wire[793];							inform_L[781][6] = l_cell_wire[794];							inform_L[845][6] = l_cell_wire[795];							inform_L[782][6] = l_cell_wire[796];							inform_L[846][6] = l_cell_wire[797];							inform_L[783][6] = l_cell_wire[798];							inform_L[847][6] = l_cell_wire[799];							inform_L[784][6] = l_cell_wire[800];							inform_L[848][6] = l_cell_wire[801];							inform_L[785][6] = l_cell_wire[802];							inform_L[849][6] = l_cell_wire[803];							inform_L[786][6] = l_cell_wire[804];							inform_L[850][6] = l_cell_wire[805];							inform_L[787][6] = l_cell_wire[806];							inform_L[851][6] = l_cell_wire[807];							inform_L[788][6] = l_cell_wire[808];							inform_L[852][6] = l_cell_wire[809];							inform_L[789][6] = l_cell_wire[810];							inform_L[853][6] = l_cell_wire[811];							inform_L[790][6] = l_cell_wire[812];							inform_L[854][6] = l_cell_wire[813];							inform_L[791][6] = l_cell_wire[814];							inform_L[855][6] = l_cell_wire[815];							inform_L[792][6] = l_cell_wire[816];							inform_L[856][6] = l_cell_wire[817];							inform_L[793][6] = l_cell_wire[818];							inform_L[857][6] = l_cell_wire[819];							inform_L[794][6] = l_cell_wire[820];							inform_L[858][6] = l_cell_wire[821];							inform_L[795][6] = l_cell_wire[822];							inform_L[859][6] = l_cell_wire[823];							inform_L[796][6] = l_cell_wire[824];							inform_L[860][6] = l_cell_wire[825];							inform_L[797][6] = l_cell_wire[826];							inform_L[861][6] = l_cell_wire[827];							inform_L[798][6] = l_cell_wire[828];							inform_L[862][6] = l_cell_wire[829];							inform_L[799][6] = l_cell_wire[830];							inform_L[863][6] = l_cell_wire[831];							inform_L[800][6] = l_cell_wire[832];							inform_L[864][6] = l_cell_wire[833];							inform_L[801][6] = l_cell_wire[834];							inform_L[865][6] = l_cell_wire[835];							inform_L[802][6] = l_cell_wire[836];							inform_L[866][6] = l_cell_wire[837];							inform_L[803][6] = l_cell_wire[838];							inform_L[867][6] = l_cell_wire[839];							inform_L[804][6] = l_cell_wire[840];							inform_L[868][6] = l_cell_wire[841];							inform_L[805][6] = l_cell_wire[842];							inform_L[869][6] = l_cell_wire[843];							inform_L[806][6] = l_cell_wire[844];							inform_L[870][6] = l_cell_wire[845];							inform_L[807][6] = l_cell_wire[846];							inform_L[871][6] = l_cell_wire[847];							inform_L[808][6] = l_cell_wire[848];							inform_L[872][6] = l_cell_wire[849];							inform_L[809][6] = l_cell_wire[850];							inform_L[873][6] = l_cell_wire[851];							inform_L[810][6] = l_cell_wire[852];							inform_L[874][6] = l_cell_wire[853];							inform_L[811][6] = l_cell_wire[854];							inform_L[875][6] = l_cell_wire[855];							inform_L[812][6] = l_cell_wire[856];							inform_L[876][6] = l_cell_wire[857];							inform_L[813][6] = l_cell_wire[858];							inform_L[877][6] = l_cell_wire[859];							inform_L[814][6] = l_cell_wire[860];							inform_L[878][6] = l_cell_wire[861];							inform_L[815][6] = l_cell_wire[862];							inform_L[879][6] = l_cell_wire[863];							inform_L[816][6] = l_cell_wire[864];							inform_L[880][6] = l_cell_wire[865];							inform_L[817][6] = l_cell_wire[866];							inform_L[881][6] = l_cell_wire[867];							inform_L[818][6] = l_cell_wire[868];							inform_L[882][6] = l_cell_wire[869];							inform_L[819][6] = l_cell_wire[870];							inform_L[883][6] = l_cell_wire[871];							inform_L[820][6] = l_cell_wire[872];							inform_L[884][6] = l_cell_wire[873];							inform_L[821][6] = l_cell_wire[874];							inform_L[885][6] = l_cell_wire[875];							inform_L[822][6] = l_cell_wire[876];							inform_L[886][6] = l_cell_wire[877];							inform_L[823][6] = l_cell_wire[878];							inform_L[887][6] = l_cell_wire[879];							inform_L[824][6] = l_cell_wire[880];							inform_L[888][6] = l_cell_wire[881];							inform_L[825][6] = l_cell_wire[882];							inform_L[889][6] = l_cell_wire[883];							inform_L[826][6] = l_cell_wire[884];							inform_L[890][6] = l_cell_wire[885];							inform_L[827][6] = l_cell_wire[886];							inform_L[891][6] = l_cell_wire[887];							inform_L[828][6] = l_cell_wire[888];							inform_L[892][6] = l_cell_wire[889];							inform_L[829][6] = l_cell_wire[890];							inform_L[893][6] = l_cell_wire[891];							inform_L[830][6] = l_cell_wire[892];							inform_L[894][6] = l_cell_wire[893];							inform_L[831][6] = l_cell_wire[894];							inform_L[895][6] = l_cell_wire[895];							inform_L[896][6] = l_cell_wire[896];							inform_L[960][6] = l_cell_wire[897];							inform_L[897][6] = l_cell_wire[898];							inform_L[961][6] = l_cell_wire[899];							inform_L[898][6] = l_cell_wire[900];							inform_L[962][6] = l_cell_wire[901];							inform_L[899][6] = l_cell_wire[902];							inform_L[963][6] = l_cell_wire[903];							inform_L[900][6] = l_cell_wire[904];							inform_L[964][6] = l_cell_wire[905];							inform_L[901][6] = l_cell_wire[906];							inform_L[965][6] = l_cell_wire[907];							inform_L[902][6] = l_cell_wire[908];							inform_L[966][6] = l_cell_wire[909];							inform_L[903][6] = l_cell_wire[910];							inform_L[967][6] = l_cell_wire[911];							inform_L[904][6] = l_cell_wire[912];							inform_L[968][6] = l_cell_wire[913];							inform_L[905][6] = l_cell_wire[914];							inform_L[969][6] = l_cell_wire[915];							inform_L[906][6] = l_cell_wire[916];							inform_L[970][6] = l_cell_wire[917];							inform_L[907][6] = l_cell_wire[918];							inform_L[971][6] = l_cell_wire[919];							inform_L[908][6] = l_cell_wire[920];							inform_L[972][6] = l_cell_wire[921];							inform_L[909][6] = l_cell_wire[922];							inform_L[973][6] = l_cell_wire[923];							inform_L[910][6] = l_cell_wire[924];							inform_L[974][6] = l_cell_wire[925];							inform_L[911][6] = l_cell_wire[926];							inform_L[975][6] = l_cell_wire[927];							inform_L[912][6] = l_cell_wire[928];							inform_L[976][6] = l_cell_wire[929];							inform_L[913][6] = l_cell_wire[930];							inform_L[977][6] = l_cell_wire[931];							inform_L[914][6] = l_cell_wire[932];							inform_L[978][6] = l_cell_wire[933];							inform_L[915][6] = l_cell_wire[934];							inform_L[979][6] = l_cell_wire[935];							inform_L[916][6] = l_cell_wire[936];							inform_L[980][6] = l_cell_wire[937];							inform_L[917][6] = l_cell_wire[938];							inform_L[981][6] = l_cell_wire[939];							inform_L[918][6] = l_cell_wire[940];							inform_L[982][6] = l_cell_wire[941];							inform_L[919][6] = l_cell_wire[942];							inform_L[983][6] = l_cell_wire[943];							inform_L[920][6] = l_cell_wire[944];							inform_L[984][6] = l_cell_wire[945];							inform_L[921][6] = l_cell_wire[946];							inform_L[985][6] = l_cell_wire[947];							inform_L[922][6] = l_cell_wire[948];							inform_L[986][6] = l_cell_wire[949];							inform_L[923][6] = l_cell_wire[950];							inform_L[987][6] = l_cell_wire[951];							inform_L[924][6] = l_cell_wire[952];							inform_L[988][6] = l_cell_wire[953];							inform_L[925][6] = l_cell_wire[954];							inform_L[989][6] = l_cell_wire[955];							inform_L[926][6] = l_cell_wire[956];							inform_L[990][6] = l_cell_wire[957];							inform_L[927][6] = l_cell_wire[958];							inform_L[991][6] = l_cell_wire[959];							inform_L[928][6] = l_cell_wire[960];							inform_L[992][6] = l_cell_wire[961];							inform_L[929][6] = l_cell_wire[962];							inform_L[993][6] = l_cell_wire[963];							inform_L[930][6] = l_cell_wire[964];							inform_L[994][6] = l_cell_wire[965];							inform_L[931][6] = l_cell_wire[966];							inform_L[995][6] = l_cell_wire[967];							inform_L[932][6] = l_cell_wire[968];							inform_L[996][6] = l_cell_wire[969];							inform_L[933][6] = l_cell_wire[970];							inform_L[997][6] = l_cell_wire[971];							inform_L[934][6] = l_cell_wire[972];							inform_L[998][6] = l_cell_wire[973];							inform_L[935][6] = l_cell_wire[974];							inform_L[999][6] = l_cell_wire[975];							inform_L[936][6] = l_cell_wire[976];							inform_L[1000][6] = l_cell_wire[977];							inform_L[937][6] = l_cell_wire[978];							inform_L[1001][6] = l_cell_wire[979];							inform_L[938][6] = l_cell_wire[980];							inform_L[1002][6] = l_cell_wire[981];							inform_L[939][6] = l_cell_wire[982];							inform_L[1003][6] = l_cell_wire[983];							inform_L[940][6] = l_cell_wire[984];							inform_L[1004][6] = l_cell_wire[985];							inform_L[941][6] = l_cell_wire[986];							inform_L[1005][6] = l_cell_wire[987];							inform_L[942][6] = l_cell_wire[988];							inform_L[1006][6] = l_cell_wire[989];							inform_L[943][6] = l_cell_wire[990];							inform_L[1007][6] = l_cell_wire[991];							inform_L[944][6] = l_cell_wire[992];							inform_L[1008][6] = l_cell_wire[993];							inform_L[945][6] = l_cell_wire[994];							inform_L[1009][6] = l_cell_wire[995];							inform_L[946][6] = l_cell_wire[996];							inform_L[1010][6] = l_cell_wire[997];							inform_L[947][6] = l_cell_wire[998];							inform_L[1011][6] = l_cell_wire[999];							inform_L[948][6] = l_cell_wire[1000];							inform_L[1012][6] = l_cell_wire[1001];							inform_L[949][6] = l_cell_wire[1002];							inform_L[1013][6] = l_cell_wire[1003];							inform_L[950][6] = l_cell_wire[1004];							inform_L[1014][6] = l_cell_wire[1005];							inform_L[951][6] = l_cell_wire[1006];							inform_L[1015][6] = l_cell_wire[1007];							inform_L[952][6] = l_cell_wire[1008];							inform_L[1016][6] = l_cell_wire[1009];							inform_L[953][6] = l_cell_wire[1010];							inform_L[1017][6] = l_cell_wire[1011];							inform_L[954][6] = l_cell_wire[1012];							inform_L[1018][6] = l_cell_wire[1013];							inform_L[955][6] = l_cell_wire[1014];							inform_L[1019][6] = l_cell_wire[1015];							inform_L[956][6] = l_cell_wire[1016];							inform_L[1020][6] = l_cell_wire[1017];							inform_L[957][6] = l_cell_wire[1018];							inform_L[1021][6] = l_cell_wire[1019];							inform_L[958][6] = l_cell_wire[1020];							inform_L[1022][6] = l_cell_wire[1021];							inform_L[959][6] = l_cell_wire[1022];							inform_L[1023][6] = l_cell_wire[1023];						end
						8:						begin							inform_R[0][8] = r_cell_wire[0];							inform_R[128][8] = r_cell_wire[1];							inform_R[1][8] = r_cell_wire[2];							inform_R[129][8] = r_cell_wire[3];							inform_R[2][8] = r_cell_wire[4];							inform_R[130][8] = r_cell_wire[5];							inform_R[3][8] = r_cell_wire[6];							inform_R[131][8] = r_cell_wire[7];							inform_R[4][8] = r_cell_wire[8];							inform_R[132][8] = r_cell_wire[9];							inform_R[5][8] = r_cell_wire[10];							inform_R[133][8] = r_cell_wire[11];							inform_R[6][8] = r_cell_wire[12];							inform_R[134][8] = r_cell_wire[13];							inform_R[7][8] = r_cell_wire[14];							inform_R[135][8] = r_cell_wire[15];							inform_R[8][8] = r_cell_wire[16];							inform_R[136][8] = r_cell_wire[17];							inform_R[9][8] = r_cell_wire[18];							inform_R[137][8] = r_cell_wire[19];							inform_R[10][8] = r_cell_wire[20];							inform_R[138][8] = r_cell_wire[21];							inform_R[11][8] = r_cell_wire[22];							inform_R[139][8] = r_cell_wire[23];							inform_R[12][8] = r_cell_wire[24];							inform_R[140][8] = r_cell_wire[25];							inform_R[13][8] = r_cell_wire[26];							inform_R[141][8] = r_cell_wire[27];							inform_R[14][8] = r_cell_wire[28];							inform_R[142][8] = r_cell_wire[29];							inform_R[15][8] = r_cell_wire[30];							inform_R[143][8] = r_cell_wire[31];							inform_R[16][8] = r_cell_wire[32];							inform_R[144][8] = r_cell_wire[33];							inform_R[17][8] = r_cell_wire[34];							inform_R[145][8] = r_cell_wire[35];							inform_R[18][8] = r_cell_wire[36];							inform_R[146][8] = r_cell_wire[37];							inform_R[19][8] = r_cell_wire[38];							inform_R[147][8] = r_cell_wire[39];							inform_R[20][8] = r_cell_wire[40];							inform_R[148][8] = r_cell_wire[41];							inform_R[21][8] = r_cell_wire[42];							inform_R[149][8] = r_cell_wire[43];							inform_R[22][8] = r_cell_wire[44];							inform_R[150][8] = r_cell_wire[45];							inform_R[23][8] = r_cell_wire[46];							inform_R[151][8] = r_cell_wire[47];							inform_R[24][8] = r_cell_wire[48];							inform_R[152][8] = r_cell_wire[49];							inform_R[25][8] = r_cell_wire[50];							inform_R[153][8] = r_cell_wire[51];							inform_R[26][8] = r_cell_wire[52];							inform_R[154][8] = r_cell_wire[53];							inform_R[27][8] = r_cell_wire[54];							inform_R[155][8] = r_cell_wire[55];							inform_R[28][8] = r_cell_wire[56];							inform_R[156][8] = r_cell_wire[57];							inform_R[29][8] = r_cell_wire[58];							inform_R[157][8] = r_cell_wire[59];							inform_R[30][8] = r_cell_wire[60];							inform_R[158][8] = r_cell_wire[61];							inform_R[31][8] = r_cell_wire[62];							inform_R[159][8] = r_cell_wire[63];							inform_R[32][8] = r_cell_wire[64];							inform_R[160][8] = r_cell_wire[65];							inform_R[33][8] = r_cell_wire[66];							inform_R[161][8] = r_cell_wire[67];							inform_R[34][8] = r_cell_wire[68];							inform_R[162][8] = r_cell_wire[69];							inform_R[35][8] = r_cell_wire[70];							inform_R[163][8] = r_cell_wire[71];							inform_R[36][8] = r_cell_wire[72];							inform_R[164][8] = r_cell_wire[73];							inform_R[37][8] = r_cell_wire[74];							inform_R[165][8] = r_cell_wire[75];							inform_R[38][8] = r_cell_wire[76];							inform_R[166][8] = r_cell_wire[77];							inform_R[39][8] = r_cell_wire[78];							inform_R[167][8] = r_cell_wire[79];							inform_R[40][8] = r_cell_wire[80];							inform_R[168][8] = r_cell_wire[81];							inform_R[41][8] = r_cell_wire[82];							inform_R[169][8] = r_cell_wire[83];							inform_R[42][8] = r_cell_wire[84];							inform_R[170][8] = r_cell_wire[85];							inform_R[43][8] = r_cell_wire[86];							inform_R[171][8] = r_cell_wire[87];							inform_R[44][8] = r_cell_wire[88];							inform_R[172][8] = r_cell_wire[89];							inform_R[45][8] = r_cell_wire[90];							inform_R[173][8] = r_cell_wire[91];							inform_R[46][8] = r_cell_wire[92];							inform_R[174][8] = r_cell_wire[93];							inform_R[47][8] = r_cell_wire[94];							inform_R[175][8] = r_cell_wire[95];							inform_R[48][8] = r_cell_wire[96];							inform_R[176][8] = r_cell_wire[97];							inform_R[49][8] = r_cell_wire[98];							inform_R[177][8] = r_cell_wire[99];							inform_R[50][8] = r_cell_wire[100];							inform_R[178][8] = r_cell_wire[101];							inform_R[51][8] = r_cell_wire[102];							inform_R[179][8] = r_cell_wire[103];							inform_R[52][8] = r_cell_wire[104];							inform_R[180][8] = r_cell_wire[105];							inform_R[53][8] = r_cell_wire[106];							inform_R[181][8] = r_cell_wire[107];							inform_R[54][8] = r_cell_wire[108];							inform_R[182][8] = r_cell_wire[109];							inform_R[55][8] = r_cell_wire[110];							inform_R[183][8] = r_cell_wire[111];							inform_R[56][8] = r_cell_wire[112];							inform_R[184][8] = r_cell_wire[113];							inform_R[57][8] = r_cell_wire[114];							inform_R[185][8] = r_cell_wire[115];							inform_R[58][8] = r_cell_wire[116];							inform_R[186][8] = r_cell_wire[117];							inform_R[59][8] = r_cell_wire[118];							inform_R[187][8] = r_cell_wire[119];							inform_R[60][8] = r_cell_wire[120];							inform_R[188][8] = r_cell_wire[121];							inform_R[61][8] = r_cell_wire[122];							inform_R[189][8] = r_cell_wire[123];							inform_R[62][8] = r_cell_wire[124];							inform_R[190][8] = r_cell_wire[125];							inform_R[63][8] = r_cell_wire[126];							inform_R[191][8] = r_cell_wire[127];							inform_R[64][8] = r_cell_wire[128];							inform_R[192][8] = r_cell_wire[129];							inform_R[65][8] = r_cell_wire[130];							inform_R[193][8] = r_cell_wire[131];							inform_R[66][8] = r_cell_wire[132];							inform_R[194][8] = r_cell_wire[133];							inform_R[67][8] = r_cell_wire[134];							inform_R[195][8] = r_cell_wire[135];							inform_R[68][8] = r_cell_wire[136];							inform_R[196][8] = r_cell_wire[137];							inform_R[69][8] = r_cell_wire[138];							inform_R[197][8] = r_cell_wire[139];							inform_R[70][8] = r_cell_wire[140];							inform_R[198][8] = r_cell_wire[141];							inform_R[71][8] = r_cell_wire[142];							inform_R[199][8] = r_cell_wire[143];							inform_R[72][8] = r_cell_wire[144];							inform_R[200][8] = r_cell_wire[145];							inform_R[73][8] = r_cell_wire[146];							inform_R[201][8] = r_cell_wire[147];							inform_R[74][8] = r_cell_wire[148];							inform_R[202][8] = r_cell_wire[149];							inform_R[75][8] = r_cell_wire[150];							inform_R[203][8] = r_cell_wire[151];							inform_R[76][8] = r_cell_wire[152];							inform_R[204][8] = r_cell_wire[153];							inform_R[77][8] = r_cell_wire[154];							inform_R[205][8] = r_cell_wire[155];							inform_R[78][8] = r_cell_wire[156];							inform_R[206][8] = r_cell_wire[157];							inform_R[79][8] = r_cell_wire[158];							inform_R[207][8] = r_cell_wire[159];							inform_R[80][8] = r_cell_wire[160];							inform_R[208][8] = r_cell_wire[161];							inform_R[81][8] = r_cell_wire[162];							inform_R[209][8] = r_cell_wire[163];							inform_R[82][8] = r_cell_wire[164];							inform_R[210][8] = r_cell_wire[165];							inform_R[83][8] = r_cell_wire[166];							inform_R[211][8] = r_cell_wire[167];							inform_R[84][8] = r_cell_wire[168];							inform_R[212][8] = r_cell_wire[169];							inform_R[85][8] = r_cell_wire[170];							inform_R[213][8] = r_cell_wire[171];							inform_R[86][8] = r_cell_wire[172];							inform_R[214][8] = r_cell_wire[173];							inform_R[87][8] = r_cell_wire[174];							inform_R[215][8] = r_cell_wire[175];							inform_R[88][8] = r_cell_wire[176];							inform_R[216][8] = r_cell_wire[177];							inform_R[89][8] = r_cell_wire[178];							inform_R[217][8] = r_cell_wire[179];							inform_R[90][8] = r_cell_wire[180];							inform_R[218][8] = r_cell_wire[181];							inform_R[91][8] = r_cell_wire[182];							inform_R[219][8] = r_cell_wire[183];							inform_R[92][8] = r_cell_wire[184];							inform_R[220][8] = r_cell_wire[185];							inform_R[93][8] = r_cell_wire[186];							inform_R[221][8] = r_cell_wire[187];							inform_R[94][8] = r_cell_wire[188];							inform_R[222][8] = r_cell_wire[189];							inform_R[95][8] = r_cell_wire[190];							inform_R[223][8] = r_cell_wire[191];							inform_R[96][8] = r_cell_wire[192];							inform_R[224][8] = r_cell_wire[193];							inform_R[97][8] = r_cell_wire[194];							inform_R[225][8] = r_cell_wire[195];							inform_R[98][8] = r_cell_wire[196];							inform_R[226][8] = r_cell_wire[197];							inform_R[99][8] = r_cell_wire[198];							inform_R[227][8] = r_cell_wire[199];							inform_R[100][8] = r_cell_wire[200];							inform_R[228][8] = r_cell_wire[201];							inform_R[101][8] = r_cell_wire[202];							inform_R[229][8] = r_cell_wire[203];							inform_R[102][8] = r_cell_wire[204];							inform_R[230][8] = r_cell_wire[205];							inform_R[103][8] = r_cell_wire[206];							inform_R[231][8] = r_cell_wire[207];							inform_R[104][8] = r_cell_wire[208];							inform_R[232][8] = r_cell_wire[209];							inform_R[105][8] = r_cell_wire[210];							inform_R[233][8] = r_cell_wire[211];							inform_R[106][8] = r_cell_wire[212];							inform_R[234][8] = r_cell_wire[213];							inform_R[107][8] = r_cell_wire[214];							inform_R[235][8] = r_cell_wire[215];							inform_R[108][8] = r_cell_wire[216];							inform_R[236][8] = r_cell_wire[217];							inform_R[109][8] = r_cell_wire[218];							inform_R[237][8] = r_cell_wire[219];							inform_R[110][8] = r_cell_wire[220];							inform_R[238][8] = r_cell_wire[221];							inform_R[111][8] = r_cell_wire[222];							inform_R[239][8] = r_cell_wire[223];							inform_R[112][8] = r_cell_wire[224];							inform_R[240][8] = r_cell_wire[225];							inform_R[113][8] = r_cell_wire[226];							inform_R[241][8] = r_cell_wire[227];							inform_R[114][8] = r_cell_wire[228];							inform_R[242][8] = r_cell_wire[229];							inform_R[115][8] = r_cell_wire[230];							inform_R[243][8] = r_cell_wire[231];							inform_R[116][8] = r_cell_wire[232];							inform_R[244][8] = r_cell_wire[233];							inform_R[117][8] = r_cell_wire[234];							inform_R[245][8] = r_cell_wire[235];							inform_R[118][8] = r_cell_wire[236];							inform_R[246][8] = r_cell_wire[237];							inform_R[119][8] = r_cell_wire[238];							inform_R[247][8] = r_cell_wire[239];							inform_R[120][8] = r_cell_wire[240];							inform_R[248][8] = r_cell_wire[241];							inform_R[121][8] = r_cell_wire[242];							inform_R[249][8] = r_cell_wire[243];							inform_R[122][8] = r_cell_wire[244];							inform_R[250][8] = r_cell_wire[245];							inform_R[123][8] = r_cell_wire[246];							inform_R[251][8] = r_cell_wire[247];							inform_R[124][8] = r_cell_wire[248];							inform_R[252][8] = r_cell_wire[249];							inform_R[125][8] = r_cell_wire[250];							inform_R[253][8] = r_cell_wire[251];							inform_R[126][8] = r_cell_wire[252];							inform_R[254][8] = r_cell_wire[253];							inform_R[127][8] = r_cell_wire[254];							inform_R[255][8] = r_cell_wire[255];							inform_R[256][8] = r_cell_wire[256];							inform_R[384][8] = r_cell_wire[257];							inform_R[257][8] = r_cell_wire[258];							inform_R[385][8] = r_cell_wire[259];							inform_R[258][8] = r_cell_wire[260];							inform_R[386][8] = r_cell_wire[261];							inform_R[259][8] = r_cell_wire[262];							inform_R[387][8] = r_cell_wire[263];							inform_R[260][8] = r_cell_wire[264];							inform_R[388][8] = r_cell_wire[265];							inform_R[261][8] = r_cell_wire[266];							inform_R[389][8] = r_cell_wire[267];							inform_R[262][8] = r_cell_wire[268];							inform_R[390][8] = r_cell_wire[269];							inform_R[263][8] = r_cell_wire[270];							inform_R[391][8] = r_cell_wire[271];							inform_R[264][8] = r_cell_wire[272];							inform_R[392][8] = r_cell_wire[273];							inform_R[265][8] = r_cell_wire[274];							inform_R[393][8] = r_cell_wire[275];							inform_R[266][8] = r_cell_wire[276];							inform_R[394][8] = r_cell_wire[277];							inform_R[267][8] = r_cell_wire[278];							inform_R[395][8] = r_cell_wire[279];							inform_R[268][8] = r_cell_wire[280];							inform_R[396][8] = r_cell_wire[281];							inform_R[269][8] = r_cell_wire[282];							inform_R[397][8] = r_cell_wire[283];							inform_R[270][8] = r_cell_wire[284];							inform_R[398][8] = r_cell_wire[285];							inform_R[271][8] = r_cell_wire[286];							inform_R[399][8] = r_cell_wire[287];							inform_R[272][8] = r_cell_wire[288];							inform_R[400][8] = r_cell_wire[289];							inform_R[273][8] = r_cell_wire[290];							inform_R[401][8] = r_cell_wire[291];							inform_R[274][8] = r_cell_wire[292];							inform_R[402][8] = r_cell_wire[293];							inform_R[275][8] = r_cell_wire[294];							inform_R[403][8] = r_cell_wire[295];							inform_R[276][8] = r_cell_wire[296];							inform_R[404][8] = r_cell_wire[297];							inform_R[277][8] = r_cell_wire[298];							inform_R[405][8] = r_cell_wire[299];							inform_R[278][8] = r_cell_wire[300];							inform_R[406][8] = r_cell_wire[301];							inform_R[279][8] = r_cell_wire[302];							inform_R[407][8] = r_cell_wire[303];							inform_R[280][8] = r_cell_wire[304];							inform_R[408][8] = r_cell_wire[305];							inform_R[281][8] = r_cell_wire[306];							inform_R[409][8] = r_cell_wire[307];							inform_R[282][8] = r_cell_wire[308];							inform_R[410][8] = r_cell_wire[309];							inform_R[283][8] = r_cell_wire[310];							inform_R[411][8] = r_cell_wire[311];							inform_R[284][8] = r_cell_wire[312];							inform_R[412][8] = r_cell_wire[313];							inform_R[285][8] = r_cell_wire[314];							inform_R[413][8] = r_cell_wire[315];							inform_R[286][8] = r_cell_wire[316];							inform_R[414][8] = r_cell_wire[317];							inform_R[287][8] = r_cell_wire[318];							inform_R[415][8] = r_cell_wire[319];							inform_R[288][8] = r_cell_wire[320];							inform_R[416][8] = r_cell_wire[321];							inform_R[289][8] = r_cell_wire[322];							inform_R[417][8] = r_cell_wire[323];							inform_R[290][8] = r_cell_wire[324];							inform_R[418][8] = r_cell_wire[325];							inform_R[291][8] = r_cell_wire[326];							inform_R[419][8] = r_cell_wire[327];							inform_R[292][8] = r_cell_wire[328];							inform_R[420][8] = r_cell_wire[329];							inform_R[293][8] = r_cell_wire[330];							inform_R[421][8] = r_cell_wire[331];							inform_R[294][8] = r_cell_wire[332];							inform_R[422][8] = r_cell_wire[333];							inform_R[295][8] = r_cell_wire[334];							inform_R[423][8] = r_cell_wire[335];							inform_R[296][8] = r_cell_wire[336];							inform_R[424][8] = r_cell_wire[337];							inform_R[297][8] = r_cell_wire[338];							inform_R[425][8] = r_cell_wire[339];							inform_R[298][8] = r_cell_wire[340];							inform_R[426][8] = r_cell_wire[341];							inform_R[299][8] = r_cell_wire[342];							inform_R[427][8] = r_cell_wire[343];							inform_R[300][8] = r_cell_wire[344];							inform_R[428][8] = r_cell_wire[345];							inform_R[301][8] = r_cell_wire[346];							inform_R[429][8] = r_cell_wire[347];							inform_R[302][8] = r_cell_wire[348];							inform_R[430][8] = r_cell_wire[349];							inform_R[303][8] = r_cell_wire[350];							inform_R[431][8] = r_cell_wire[351];							inform_R[304][8] = r_cell_wire[352];							inform_R[432][8] = r_cell_wire[353];							inform_R[305][8] = r_cell_wire[354];							inform_R[433][8] = r_cell_wire[355];							inform_R[306][8] = r_cell_wire[356];							inform_R[434][8] = r_cell_wire[357];							inform_R[307][8] = r_cell_wire[358];							inform_R[435][8] = r_cell_wire[359];							inform_R[308][8] = r_cell_wire[360];							inform_R[436][8] = r_cell_wire[361];							inform_R[309][8] = r_cell_wire[362];							inform_R[437][8] = r_cell_wire[363];							inform_R[310][8] = r_cell_wire[364];							inform_R[438][8] = r_cell_wire[365];							inform_R[311][8] = r_cell_wire[366];							inform_R[439][8] = r_cell_wire[367];							inform_R[312][8] = r_cell_wire[368];							inform_R[440][8] = r_cell_wire[369];							inform_R[313][8] = r_cell_wire[370];							inform_R[441][8] = r_cell_wire[371];							inform_R[314][8] = r_cell_wire[372];							inform_R[442][8] = r_cell_wire[373];							inform_R[315][8] = r_cell_wire[374];							inform_R[443][8] = r_cell_wire[375];							inform_R[316][8] = r_cell_wire[376];							inform_R[444][8] = r_cell_wire[377];							inform_R[317][8] = r_cell_wire[378];							inform_R[445][8] = r_cell_wire[379];							inform_R[318][8] = r_cell_wire[380];							inform_R[446][8] = r_cell_wire[381];							inform_R[319][8] = r_cell_wire[382];							inform_R[447][8] = r_cell_wire[383];							inform_R[320][8] = r_cell_wire[384];							inform_R[448][8] = r_cell_wire[385];							inform_R[321][8] = r_cell_wire[386];							inform_R[449][8] = r_cell_wire[387];							inform_R[322][8] = r_cell_wire[388];							inform_R[450][8] = r_cell_wire[389];							inform_R[323][8] = r_cell_wire[390];							inform_R[451][8] = r_cell_wire[391];							inform_R[324][8] = r_cell_wire[392];							inform_R[452][8] = r_cell_wire[393];							inform_R[325][8] = r_cell_wire[394];							inform_R[453][8] = r_cell_wire[395];							inform_R[326][8] = r_cell_wire[396];							inform_R[454][8] = r_cell_wire[397];							inform_R[327][8] = r_cell_wire[398];							inform_R[455][8] = r_cell_wire[399];							inform_R[328][8] = r_cell_wire[400];							inform_R[456][8] = r_cell_wire[401];							inform_R[329][8] = r_cell_wire[402];							inform_R[457][8] = r_cell_wire[403];							inform_R[330][8] = r_cell_wire[404];							inform_R[458][8] = r_cell_wire[405];							inform_R[331][8] = r_cell_wire[406];							inform_R[459][8] = r_cell_wire[407];							inform_R[332][8] = r_cell_wire[408];							inform_R[460][8] = r_cell_wire[409];							inform_R[333][8] = r_cell_wire[410];							inform_R[461][8] = r_cell_wire[411];							inform_R[334][8] = r_cell_wire[412];							inform_R[462][8] = r_cell_wire[413];							inform_R[335][8] = r_cell_wire[414];							inform_R[463][8] = r_cell_wire[415];							inform_R[336][8] = r_cell_wire[416];							inform_R[464][8] = r_cell_wire[417];							inform_R[337][8] = r_cell_wire[418];							inform_R[465][8] = r_cell_wire[419];							inform_R[338][8] = r_cell_wire[420];							inform_R[466][8] = r_cell_wire[421];							inform_R[339][8] = r_cell_wire[422];							inform_R[467][8] = r_cell_wire[423];							inform_R[340][8] = r_cell_wire[424];							inform_R[468][8] = r_cell_wire[425];							inform_R[341][8] = r_cell_wire[426];							inform_R[469][8] = r_cell_wire[427];							inform_R[342][8] = r_cell_wire[428];							inform_R[470][8] = r_cell_wire[429];							inform_R[343][8] = r_cell_wire[430];							inform_R[471][8] = r_cell_wire[431];							inform_R[344][8] = r_cell_wire[432];							inform_R[472][8] = r_cell_wire[433];							inform_R[345][8] = r_cell_wire[434];							inform_R[473][8] = r_cell_wire[435];							inform_R[346][8] = r_cell_wire[436];							inform_R[474][8] = r_cell_wire[437];							inform_R[347][8] = r_cell_wire[438];							inform_R[475][8] = r_cell_wire[439];							inform_R[348][8] = r_cell_wire[440];							inform_R[476][8] = r_cell_wire[441];							inform_R[349][8] = r_cell_wire[442];							inform_R[477][8] = r_cell_wire[443];							inform_R[350][8] = r_cell_wire[444];							inform_R[478][8] = r_cell_wire[445];							inform_R[351][8] = r_cell_wire[446];							inform_R[479][8] = r_cell_wire[447];							inform_R[352][8] = r_cell_wire[448];							inform_R[480][8] = r_cell_wire[449];							inform_R[353][8] = r_cell_wire[450];							inform_R[481][8] = r_cell_wire[451];							inform_R[354][8] = r_cell_wire[452];							inform_R[482][8] = r_cell_wire[453];							inform_R[355][8] = r_cell_wire[454];							inform_R[483][8] = r_cell_wire[455];							inform_R[356][8] = r_cell_wire[456];							inform_R[484][8] = r_cell_wire[457];							inform_R[357][8] = r_cell_wire[458];							inform_R[485][8] = r_cell_wire[459];							inform_R[358][8] = r_cell_wire[460];							inform_R[486][8] = r_cell_wire[461];							inform_R[359][8] = r_cell_wire[462];							inform_R[487][8] = r_cell_wire[463];							inform_R[360][8] = r_cell_wire[464];							inform_R[488][8] = r_cell_wire[465];							inform_R[361][8] = r_cell_wire[466];							inform_R[489][8] = r_cell_wire[467];							inform_R[362][8] = r_cell_wire[468];							inform_R[490][8] = r_cell_wire[469];							inform_R[363][8] = r_cell_wire[470];							inform_R[491][8] = r_cell_wire[471];							inform_R[364][8] = r_cell_wire[472];							inform_R[492][8] = r_cell_wire[473];							inform_R[365][8] = r_cell_wire[474];							inform_R[493][8] = r_cell_wire[475];							inform_R[366][8] = r_cell_wire[476];							inform_R[494][8] = r_cell_wire[477];							inform_R[367][8] = r_cell_wire[478];							inform_R[495][8] = r_cell_wire[479];							inform_R[368][8] = r_cell_wire[480];							inform_R[496][8] = r_cell_wire[481];							inform_R[369][8] = r_cell_wire[482];							inform_R[497][8] = r_cell_wire[483];							inform_R[370][8] = r_cell_wire[484];							inform_R[498][8] = r_cell_wire[485];							inform_R[371][8] = r_cell_wire[486];							inform_R[499][8] = r_cell_wire[487];							inform_R[372][8] = r_cell_wire[488];							inform_R[500][8] = r_cell_wire[489];							inform_R[373][8] = r_cell_wire[490];							inform_R[501][8] = r_cell_wire[491];							inform_R[374][8] = r_cell_wire[492];							inform_R[502][8] = r_cell_wire[493];							inform_R[375][8] = r_cell_wire[494];							inform_R[503][8] = r_cell_wire[495];							inform_R[376][8] = r_cell_wire[496];							inform_R[504][8] = r_cell_wire[497];							inform_R[377][8] = r_cell_wire[498];							inform_R[505][8] = r_cell_wire[499];							inform_R[378][8] = r_cell_wire[500];							inform_R[506][8] = r_cell_wire[501];							inform_R[379][8] = r_cell_wire[502];							inform_R[507][8] = r_cell_wire[503];							inform_R[380][8] = r_cell_wire[504];							inform_R[508][8] = r_cell_wire[505];							inform_R[381][8] = r_cell_wire[506];							inform_R[509][8] = r_cell_wire[507];							inform_R[382][8] = r_cell_wire[508];							inform_R[510][8] = r_cell_wire[509];							inform_R[383][8] = r_cell_wire[510];							inform_R[511][8] = r_cell_wire[511];							inform_R[512][8] = r_cell_wire[512];							inform_R[640][8] = r_cell_wire[513];							inform_R[513][8] = r_cell_wire[514];							inform_R[641][8] = r_cell_wire[515];							inform_R[514][8] = r_cell_wire[516];							inform_R[642][8] = r_cell_wire[517];							inform_R[515][8] = r_cell_wire[518];							inform_R[643][8] = r_cell_wire[519];							inform_R[516][8] = r_cell_wire[520];							inform_R[644][8] = r_cell_wire[521];							inform_R[517][8] = r_cell_wire[522];							inform_R[645][8] = r_cell_wire[523];							inform_R[518][8] = r_cell_wire[524];							inform_R[646][8] = r_cell_wire[525];							inform_R[519][8] = r_cell_wire[526];							inform_R[647][8] = r_cell_wire[527];							inform_R[520][8] = r_cell_wire[528];							inform_R[648][8] = r_cell_wire[529];							inform_R[521][8] = r_cell_wire[530];							inform_R[649][8] = r_cell_wire[531];							inform_R[522][8] = r_cell_wire[532];							inform_R[650][8] = r_cell_wire[533];							inform_R[523][8] = r_cell_wire[534];							inform_R[651][8] = r_cell_wire[535];							inform_R[524][8] = r_cell_wire[536];							inform_R[652][8] = r_cell_wire[537];							inform_R[525][8] = r_cell_wire[538];							inform_R[653][8] = r_cell_wire[539];							inform_R[526][8] = r_cell_wire[540];							inform_R[654][8] = r_cell_wire[541];							inform_R[527][8] = r_cell_wire[542];							inform_R[655][8] = r_cell_wire[543];							inform_R[528][8] = r_cell_wire[544];							inform_R[656][8] = r_cell_wire[545];							inform_R[529][8] = r_cell_wire[546];							inform_R[657][8] = r_cell_wire[547];							inform_R[530][8] = r_cell_wire[548];							inform_R[658][8] = r_cell_wire[549];							inform_R[531][8] = r_cell_wire[550];							inform_R[659][8] = r_cell_wire[551];							inform_R[532][8] = r_cell_wire[552];							inform_R[660][8] = r_cell_wire[553];							inform_R[533][8] = r_cell_wire[554];							inform_R[661][8] = r_cell_wire[555];							inform_R[534][8] = r_cell_wire[556];							inform_R[662][8] = r_cell_wire[557];							inform_R[535][8] = r_cell_wire[558];							inform_R[663][8] = r_cell_wire[559];							inform_R[536][8] = r_cell_wire[560];							inform_R[664][8] = r_cell_wire[561];							inform_R[537][8] = r_cell_wire[562];							inform_R[665][8] = r_cell_wire[563];							inform_R[538][8] = r_cell_wire[564];							inform_R[666][8] = r_cell_wire[565];							inform_R[539][8] = r_cell_wire[566];							inform_R[667][8] = r_cell_wire[567];							inform_R[540][8] = r_cell_wire[568];							inform_R[668][8] = r_cell_wire[569];							inform_R[541][8] = r_cell_wire[570];							inform_R[669][8] = r_cell_wire[571];							inform_R[542][8] = r_cell_wire[572];							inform_R[670][8] = r_cell_wire[573];							inform_R[543][8] = r_cell_wire[574];							inform_R[671][8] = r_cell_wire[575];							inform_R[544][8] = r_cell_wire[576];							inform_R[672][8] = r_cell_wire[577];							inform_R[545][8] = r_cell_wire[578];							inform_R[673][8] = r_cell_wire[579];							inform_R[546][8] = r_cell_wire[580];							inform_R[674][8] = r_cell_wire[581];							inform_R[547][8] = r_cell_wire[582];							inform_R[675][8] = r_cell_wire[583];							inform_R[548][8] = r_cell_wire[584];							inform_R[676][8] = r_cell_wire[585];							inform_R[549][8] = r_cell_wire[586];							inform_R[677][8] = r_cell_wire[587];							inform_R[550][8] = r_cell_wire[588];							inform_R[678][8] = r_cell_wire[589];							inform_R[551][8] = r_cell_wire[590];							inform_R[679][8] = r_cell_wire[591];							inform_R[552][8] = r_cell_wire[592];							inform_R[680][8] = r_cell_wire[593];							inform_R[553][8] = r_cell_wire[594];							inform_R[681][8] = r_cell_wire[595];							inform_R[554][8] = r_cell_wire[596];							inform_R[682][8] = r_cell_wire[597];							inform_R[555][8] = r_cell_wire[598];							inform_R[683][8] = r_cell_wire[599];							inform_R[556][8] = r_cell_wire[600];							inform_R[684][8] = r_cell_wire[601];							inform_R[557][8] = r_cell_wire[602];							inform_R[685][8] = r_cell_wire[603];							inform_R[558][8] = r_cell_wire[604];							inform_R[686][8] = r_cell_wire[605];							inform_R[559][8] = r_cell_wire[606];							inform_R[687][8] = r_cell_wire[607];							inform_R[560][8] = r_cell_wire[608];							inform_R[688][8] = r_cell_wire[609];							inform_R[561][8] = r_cell_wire[610];							inform_R[689][8] = r_cell_wire[611];							inform_R[562][8] = r_cell_wire[612];							inform_R[690][8] = r_cell_wire[613];							inform_R[563][8] = r_cell_wire[614];							inform_R[691][8] = r_cell_wire[615];							inform_R[564][8] = r_cell_wire[616];							inform_R[692][8] = r_cell_wire[617];							inform_R[565][8] = r_cell_wire[618];							inform_R[693][8] = r_cell_wire[619];							inform_R[566][8] = r_cell_wire[620];							inform_R[694][8] = r_cell_wire[621];							inform_R[567][8] = r_cell_wire[622];							inform_R[695][8] = r_cell_wire[623];							inform_R[568][8] = r_cell_wire[624];							inform_R[696][8] = r_cell_wire[625];							inform_R[569][8] = r_cell_wire[626];							inform_R[697][8] = r_cell_wire[627];							inform_R[570][8] = r_cell_wire[628];							inform_R[698][8] = r_cell_wire[629];							inform_R[571][8] = r_cell_wire[630];							inform_R[699][8] = r_cell_wire[631];							inform_R[572][8] = r_cell_wire[632];							inform_R[700][8] = r_cell_wire[633];							inform_R[573][8] = r_cell_wire[634];							inform_R[701][8] = r_cell_wire[635];							inform_R[574][8] = r_cell_wire[636];							inform_R[702][8] = r_cell_wire[637];							inform_R[575][8] = r_cell_wire[638];							inform_R[703][8] = r_cell_wire[639];							inform_R[576][8] = r_cell_wire[640];							inform_R[704][8] = r_cell_wire[641];							inform_R[577][8] = r_cell_wire[642];							inform_R[705][8] = r_cell_wire[643];							inform_R[578][8] = r_cell_wire[644];							inform_R[706][8] = r_cell_wire[645];							inform_R[579][8] = r_cell_wire[646];							inform_R[707][8] = r_cell_wire[647];							inform_R[580][8] = r_cell_wire[648];							inform_R[708][8] = r_cell_wire[649];							inform_R[581][8] = r_cell_wire[650];							inform_R[709][8] = r_cell_wire[651];							inform_R[582][8] = r_cell_wire[652];							inform_R[710][8] = r_cell_wire[653];							inform_R[583][8] = r_cell_wire[654];							inform_R[711][8] = r_cell_wire[655];							inform_R[584][8] = r_cell_wire[656];							inform_R[712][8] = r_cell_wire[657];							inform_R[585][8] = r_cell_wire[658];							inform_R[713][8] = r_cell_wire[659];							inform_R[586][8] = r_cell_wire[660];							inform_R[714][8] = r_cell_wire[661];							inform_R[587][8] = r_cell_wire[662];							inform_R[715][8] = r_cell_wire[663];							inform_R[588][8] = r_cell_wire[664];							inform_R[716][8] = r_cell_wire[665];							inform_R[589][8] = r_cell_wire[666];							inform_R[717][8] = r_cell_wire[667];							inform_R[590][8] = r_cell_wire[668];							inform_R[718][8] = r_cell_wire[669];							inform_R[591][8] = r_cell_wire[670];							inform_R[719][8] = r_cell_wire[671];							inform_R[592][8] = r_cell_wire[672];							inform_R[720][8] = r_cell_wire[673];							inform_R[593][8] = r_cell_wire[674];							inform_R[721][8] = r_cell_wire[675];							inform_R[594][8] = r_cell_wire[676];							inform_R[722][8] = r_cell_wire[677];							inform_R[595][8] = r_cell_wire[678];							inform_R[723][8] = r_cell_wire[679];							inform_R[596][8] = r_cell_wire[680];							inform_R[724][8] = r_cell_wire[681];							inform_R[597][8] = r_cell_wire[682];							inform_R[725][8] = r_cell_wire[683];							inform_R[598][8] = r_cell_wire[684];							inform_R[726][8] = r_cell_wire[685];							inform_R[599][8] = r_cell_wire[686];							inform_R[727][8] = r_cell_wire[687];							inform_R[600][8] = r_cell_wire[688];							inform_R[728][8] = r_cell_wire[689];							inform_R[601][8] = r_cell_wire[690];							inform_R[729][8] = r_cell_wire[691];							inform_R[602][8] = r_cell_wire[692];							inform_R[730][8] = r_cell_wire[693];							inform_R[603][8] = r_cell_wire[694];							inform_R[731][8] = r_cell_wire[695];							inform_R[604][8] = r_cell_wire[696];							inform_R[732][8] = r_cell_wire[697];							inform_R[605][8] = r_cell_wire[698];							inform_R[733][8] = r_cell_wire[699];							inform_R[606][8] = r_cell_wire[700];							inform_R[734][8] = r_cell_wire[701];							inform_R[607][8] = r_cell_wire[702];							inform_R[735][8] = r_cell_wire[703];							inform_R[608][8] = r_cell_wire[704];							inform_R[736][8] = r_cell_wire[705];							inform_R[609][8] = r_cell_wire[706];							inform_R[737][8] = r_cell_wire[707];							inform_R[610][8] = r_cell_wire[708];							inform_R[738][8] = r_cell_wire[709];							inform_R[611][8] = r_cell_wire[710];							inform_R[739][8] = r_cell_wire[711];							inform_R[612][8] = r_cell_wire[712];							inform_R[740][8] = r_cell_wire[713];							inform_R[613][8] = r_cell_wire[714];							inform_R[741][8] = r_cell_wire[715];							inform_R[614][8] = r_cell_wire[716];							inform_R[742][8] = r_cell_wire[717];							inform_R[615][8] = r_cell_wire[718];							inform_R[743][8] = r_cell_wire[719];							inform_R[616][8] = r_cell_wire[720];							inform_R[744][8] = r_cell_wire[721];							inform_R[617][8] = r_cell_wire[722];							inform_R[745][8] = r_cell_wire[723];							inform_R[618][8] = r_cell_wire[724];							inform_R[746][8] = r_cell_wire[725];							inform_R[619][8] = r_cell_wire[726];							inform_R[747][8] = r_cell_wire[727];							inform_R[620][8] = r_cell_wire[728];							inform_R[748][8] = r_cell_wire[729];							inform_R[621][8] = r_cell_wire[730];							inform_R[749][8] = r_cell_wire[731];							inform_R[622][8] = r_cell_wire[732];							inform_R[750][8] = r_cell_wire[733];							inform_R[623][8] = r_cell_wire[734];							inform_R[751][8] = r_cell_wire[735];							inform_R[624][8] = r_cell_wire[736];							inform_R[752][8] = r_cell_wire[737];							inform_R[625][8] = r_cell_wire[738];							inform_R[753][8] = r_cell_wire[739];							inform_R[626][8] = r_cell_wire[740];							inform_R[754][8] = r_cell_wire[741];							inform_R[627][8] = r_cell_wire[742];							inform_R[755][8] = r_cell_wire[743];							inform_R[628][8] = r_cell_wire[744];							inform_R[756][8] = r_cell_wire[745];							inform_R[629][8] = r_cell_wire[746];							inform_R[757][8] = r_cell_wire[747];							inform_R[630][8] = r_cell_wire[748];							inform_R[758][8] = r_cell_wire[749];							inform_R[631][8] = r_cell_wire[750];							inform_R[759][8] = r_cell_wire[751];							inform_R[632][8] = r_cell_wire[752];							inform_R[760][8] = r_cell_wire[753];							inform_R[633][8] = r_cell_wire[754];							inform_R[761][8] = r_cell_wire[755];							inform_R[634][8] = r_cell_wire[756];							inform_R[762][8] = r_cell_wire[757];							inform_R[635][8] = r_cell_wire[758];							inform_R[763][8] = r_cell_wire[759];							inform_R[636][8] = r_cell_wire[760];							inform_R[764][8] = r_cell_wire[761];							inform_R[637][8] = r_cell_wire[762];							inform_R[765][8] = r_cell_wire[763];							inform_R[638][8] = r_cell_wire[764];							inform_R[766][8] = r_cell_wire[765];							inform_R[639][8] = r_cell_wire[766];							inform_R[767][8] = r_cell_wire[767];							inform_R[768][8] = r_cell_wire[768];							inform_R[896][8] = r_cell_wire[769];							inform_R[769][8] = r_cell_wire[770];							inform_R[897][8] = r_cell_wire[771];							inform_R[770][8] = r_cell_wire[772];							inform_R[898][8] = r_cell_wire[773];							inform_R[771][8] = r_cell_wire[774];							inform_R[899][8] = r_cell_wire[775];							inform_R[772][8] = r_cell_wire[776];							inform_R[900][8] = r_cell_wire[777];							inform_R[773][8] = r_cell_wire[778];							inform_R[901][8] = r_cell_wire[779];							inform_R[774][8] = r_cell_wire[780];							inform_R[902][8] = r_cell_wire[781];							inform_R[775][8] = r_cell_wire[782];							inform_R[903][8] = r_cell_wire[783];							inform_R[776][8] = r_cell_wire[784];							inform_R[904][8] = r_cell_wire[785];							inform_R[777][8] = r_cell_wire[786];							inform_R[905][8] = r_cell_wire[787];							inform_R[778][8] = r_cell_wire[788];							inform_R[906][8] = r_cell_wire[789];							inform_R[779][8] = r_cell_wire[790];							inform_R[907][8] = r_cell_wire[791];							inform_R[780][8] = r_cell_wire[792];							inform_R[908][8] = r_cell_wire[793];							inform_R[781][8] = r_cell_wire[794];							inform_R[909][8] = r_cell_wire[795];							inform_R[782][8] = r_cell_wire[796];							inform_R[910][8] = r_cell_wire[797];							inform_R[783][8] = r_cell_wire[798];							inform_R[911][8] = r_cell_wire[799];							inform_R[784][8] = r_cell_wire[800];							inform_R[912][8] = r_cell_wire[801];							inform_R[785][8] = r_cell_wire[802];							inform_R[913][8] = r_cell_wire[803];							inform_R[786][8] = r_cell_wire[804];							inform_R[914][8] = r_cell_wire[805];							inform_R[787][8] = r_cell_wire[806];							inform_R[915][8] = r_cell_wire[807];							inform_R[788][8] = r_cell_wire[808];							inform_R[916][8] = r_cell_wire[809];							inform_R[789][8] = r_cell_wire[810];							inform_R[917][8] = r_cell_wire[811];							inform_R[790][8] = r_cell_wire[812];							inform_R[918][8] = r_cell_wire[813];							inform_R[791][8] = r_cell_wire[814];							inform_R[919][8] = r_cell_wire[815];							inform_R[792][8] = r_cell_wire[816];							inform_R[920][8] = r_cell_wire[817];							inform_R[793][8] = r_cell_wire[818];							inform_R[921][8] = r_cell_wire[819];							inform_R[794][8] = r_cell_wire[820];							inform_R[922][8] = r_cell_wire[821];							inform_R[795][8] = r_cell_wire[822];							inform_R[923][8] = r_cell_wire[823];							inform_R[796][8] = r_cell_wire[824];							inform_R[924][8] = r_cell_wire[825];							inform_R[797][8] = r_cell_wire[826];							inform_R[925][8] = r_cell_wire[827];							inform_R[798][8] = r_cell_wire[828];							inform_R[926][8] = r_cell_wire[829];							inform_R[799][8] = r_cell_wire[830];							inform_R[927][8] = r_cell_wire[831];							inform_R[800][8] = r_cell_wire[832];							inform_R[928][8] = r_cell_wire[833];							inform_R[801][8] = r_cell_wire[834];							inform_R[929][8] = r_cell_wire[835];							inform_R[802][8] = r_cell_wire[836];							inform_R[930][8] = r_cell_wire[837];							inform_R[803][8] = r_cell_wire[838];							inform_R[931][8] = r_cell_wire[839];							inform_R[804][8] = r_cell_wire[840];							inform_R[932][8] = r_cell_wire[841];							inform_R[805][8] = r_cell_wire[842];							inform_R[933][8] = r_cell_wire[843];							inform_R[806][8] = r_cell_wire[844];							inform_R[934][8] = r_cell_wire[845];							inform_R[807][8] = r_cell_wire[846];							inform_R[935][8] = r_cell_wire[847];							inform_R[808][8] = r_cell_wire[848];							inform_R[936][8] = r_cell_wire[849];							inform_R[809][8] = r_cell_wire[850];							inform_R[937][8] = r_cell_wire[851];							inform_R[810][8] = r_cell_wire[852];							inform_R[938][8] = r_cell_wire[853];							inform_R[811][8] = r_cell_wire[854];							inform_R[939][8] = r_cell_wire[855];							inform_R[812][8] = r_cell_wire[856];							inform_R[940][8] = r_cell_wire[857];							inform_R[813][8] = r_cell_wire[858];							inform_R[941][8] = r_cell_wire[859];							inform_R[814][8] = r_cell_wire[860];							inform_R[942][8] = r_cell_wire[861];							inform_R[815][8] = r_cell_wire[862];							inform_R[943][8] = r_cell_wire[863];							inform_R[816][8] = r_cell_wire[864];							inform_R[944][8] = r_cell_wire[865];							inform_R[817][8] = r_cell_wire[866];							inform_R[945][8] = r_cell_wire[867];							inform_R[818][8] = r_cell_wire[868];							inform_R[946][8] = r_cell_wire[869];							inform_R[819][8] = r_cell_wire[870];							inform_R[947][8] = r_cell_wire[871];							inform_R[820][8] = r_cell_wire[872];							inform_R[948][8] = r_cell_wire[873];							inform_R[821][8] = r_cell_wire[874];							inform_R[949][8] = r_cell_wire[875];							inform_R[822][8] = r_cell_wire[876];							inform_R[950][8] = r_cell_wire[877];							inform_R[823][8] = r_cell_wire[878];							inform_R[951][8] = r_cell_wire[879];							inform_R[824][8] = r_cell_wire[880];							inform_R[952][8] = r_cell_wire[881];							inform_R[825][8] = r_cell_wire[882];							inform_R[953][8] = r_cell_wire[883];							inform_R[826][8] = r_cell_wire[884];							inform_R[954][8] = r_cell_wire[885];							inform_R[827][8] = r_cell_wire[886];							inform_R[955][8] = r_cell_wire[887];							inform_R[828][8] = r_cell_wire[888];							inform_R[956][8] = r_cell_wire[889];							inform_R[829][8] = r_cell_wire[890];							inform_R[957][8] = r_cell_wire[891];							inform_R[830][8] = r_cell_wire[892];							inform_R[958][8] = r_cell_wire[893];							inform_R[831][8] = r_cell_wire[894];							inform_R[959][8] = r_cell_wire[895];							inform_R[832][8] = r_cell_wire[896];							inform_R[960][8] = r_cell_wire[897];							inform_R[833][8] = r_cell_wire[898];							inform_R[961][8] = r_cell_wire[899];							inform_R[834][8] = r_cell_wire[900];							inform_R[962][8] = r_cell_wire[901];							inform_R[835][8] = r_cell_wire[902];							inform_R[963][8] = r_cell_wire[903];							inform_R[836][8] = r_cell_wire[904];							inform_R[964][8] = r_cell_wire[905];							inform_R[837][8] = r_cell_wire[906];							inform_R[965][8] = r_cell_wire[907];							inform_R[838][8] = r_cell_wire[908];							inform_R[966][8] = r_cell_wire[909];							inform_R[839][8] = r_cell_wire[910];							inform_R[967][8] = r_cell_wire[911];							inform_R[840][8] = r_cell_wire[912];							inform_R[968][8] = r_cell_wire[913];							inform_R[841][8] = r_cell_wire[914];							inform_R[969][8] = r_cell_wire[915];							inform_R[842][8] = r_cell_wire[916];							inform_R[970][8] = r_cell_wire[917];							inform_R[843][8] = r_cell_wire[918];							inform_R[971][8] = r_cell_wire[919];							inform_R[844][8] = r_cell_wire[920];							inform_R[972][8] = r_cell_wire[921];							inform_R[845][8] = r_cell_wire[922];							inform_R[973][8] = r_cell_wire[923];							inform_R[846][8] = r_cell_wire[924];							inform_R[974][8] = r_cell_wire[925];							inform_R[847][8] = r_cell_wire[926];							inform_R[975][8] = r_cell_wire[927];							inform_R[848][8] = r_cell_wire[928];							inform_R[976][8] = r_cell_wire[929];							inform_R[849][8] = r_cell_wire[930];							inform_R[977][8] = r_cell_wire[931];							inform_R[850][8] = r_cell_wire[932];							inform_R[978][8] = r_cell_wire[933];							inform_R[851][8] = r_cell_wire[934];							inform_R[979][8] = r_cell_wire[935];							inform_R[852][8] = r_cell_wire[936];							inform_R[980][8] = r_cell_wire[937];							inform_R[853][8] = r_cell_wire[938];							inform_R[981][8] = r_cell_wire[939];							inform_R[854][8] = r_cell_wire[940];							inform_R[982][8] = r_cell_wire[941];							inform_R[855][8] = r_cell_wire[942];							inform_R[983][8] = r_cell_wire[943];							inform_R[856][8] = r_cell_wire[944];							inform_R[984][8] = r_cell_wire[945];							inform_R[857][8] = r_cell_wire[946];							inform_R[985][8] = r_cell_wire[947];							inform_R[858][8] = r_cell_wire[948];							inform_R[986][8] = r_cell_wire[949];							inform_R[859][8] = r_cell_wire[950];							inform_R[987][8] = r_cell_wire[951];							inform_R[860][8] = r_cell_wire[952];							inform_R[988][8] = r_cell_wire[953];							inform_R[861][8] = r_cell_wire[954];							inform_R[989][8] = r_cell_wire[955];							inform_R[862][8] = r_cell_wire[956];							inform_R[990][8] = r_cell_wire[957];							inform_R[863][8] = r_cell_wire[958];							inform_R[991][8] = r_cell_wire[959];							inform_R[864][8] = r_cell_wire[960];							inform_R[992][8] = r_cell_wire[961];							inform_R[865][8] = r_cell_wire[962];							inform_R[993][8] = r_cell_wire[963];							inform_R[866][8] = r_cell_wire[964];							inform_R[994][8] = r_cell_wire[965];							inform_R[867][8] = r_cell_wire[966];							inform_R[995][8] = r_cell_wire[967];							inform_R[868][8] = r_cell_wire[968];							inform_R[996][8] = r_cell_wire[969];							inform_R[869][8] = r_cell_wire[970];							inform_R[997][8] = r_cell_wire[971];							inform_R[870][8] = r_cell_wire[972];							inform_R[998][8] = r_cell_wire[973];							inform_R[871][8] = r_cell_wire[974];							inform_R[999][8] = r_cell_wire[975];							inform_R[872][8] = r_cell_wire[976];							inform_R[1000][8] = r_cell_wire[977];							inform_R[873][8] = r_cell_wire[978];							inform_R[1001][8] = r_cell_wire[979];							inform_R[874][8] = r_cell_wire[980];							inform_R[1002][8] = r_cell_wire[981];							inform_R[875][8] = r_cell_wire[982];							inform_R[1003][8] = r_cell_wire[983];							inform_R[876][8] = r_cell_wire[984];							inform_R[1004][8] = r_cell_wire[985];							inform_R[877][8] = r_cell_wire[986];							inform_R[1005][8] = r_cell_wire[987];							inform_R[878][8] = r_cell_wire[988];							inform_R[1006][8] = r_cell_wire[989];							inform_R[879][8] = r_cell_wire[990];							inform_R[1007][8] = r_cell_wire[991];							inform_R[880][8] = r_cell_wire[992];							inform_R[1008][8] = r_cell_wire[993];							inform_R[881][8] = r_cell_wire[994];							inform_R[1009][8] = r_cell_wire[995];							inform_R[882][8] = r_cell_wire[996];							inform_R[1010][8] = r_cell_wire[997];							inform_R[883][8] = r_cell_wire[998];							inform_R[1011][8] = r_cell_wire[999];							inform_R[884][8] = r_cell_wire[1000];							inform_R[1012][8] = r_cell_wire[1001];							inform_R[885][8] = r_cell_wire[1002];							inform_R[1013][8] = r_cell_wire[1003];							inform_R[886][8] = r_cell_wire[1004];							inform_R[1014][8] = r_cell_wire[1005];							inform_R[887][8] = r_cell_wire[1006];							inform_R[1015][8] = r_cell_wire[1007];							inform_R[888][8] = r_cell_wire[1008];							inform_R[1016][8] = r_cell_wire[1009];							inform_R[889][8] = r_cell_wire[1010];							inform_R[1017][8] = r_cell_wire[1011];							inform_R[890][8] = r_cell_wire[1012];							inform_R[1018][8] = r_cell_wire[1013];							inform_R[891][8] = r_cell_wire[1014];							inform_R[1019][8] = r_cell_wire[1015];							inform_R[892][8] = r_cell_wire[1016];							inform_R[1020][8] = r_cell_wire[1017];							inform_R[893][8] = r_cell_wire[1018];							inform_R[1021][8] = r_cell_wire[1019];							inform_R[894][8] = r_cell_wire[1020];							inform_R[1022][8] = r_cell_wire[1021];							inform_R[895][8] = r_cell_wire[1022];							inform_R[1023][8] = r_cell_wire[1023];							inform_L[0][7] = l_cell_wire[0];							inform_L[128][7] = l_cell_wire[1];							inform_L[1][7] = l_cell_wire[2];							inform_L[129][7] = l_cell_wire[3];							inform_L[2][7] = l_cell_wire[4];							inform_L[130][7] = l_cell_wire[5];							inform_L[3][7] = l_cell_wire[6];							inform_L[131][7] = l_cell_wire[7];							inform_L[4][7] = l_cell_wire[8];							inform_L[132][7] = l_cell_wire[9];							inform_L[5][7] = l_cell_wire[10];							inform_L[133][7] = l_cell_wire[11];							inform_L[6][7] = l_cell_wire[12];							inform_L[134][7] = l_cell_wire[13];							inform_L[7][7] = l_cell_wire[14];							inform_L[135][7] = l_cell_wire[15];							inform_L[8][7] = l_cell_wire[16];							inform_L[136][7] = l_cell_wire[17];							inform_L[9][7] = l_cell_wire[18];							inform_L[137][7] = l_cell_wire[19];							inform_L[10][7] = l_cell_wire[20];							inform_L[138][7] = l_cell_wire[21];							inform_L[11][7] = l_cell_wire[22];							inform_L[139][7] = l_cell_wire[23];							inform_L[12][7] = l_cell_wire[24];							inform_L[140][7] = l_cell_wire[25];							inform_L[13][7] = l_cell_wire[26];							inform_L[141][7] = l_cell_wire[27];							inform_L[14][7] = l_cell_wire[28];							inform_L[142][7] = l_cell_wire[29];							inform_L[15][7] = l_cell_wire[30];							inform_L[143][7] = l_cell_wire[31];							inform_L[16][7] = l_cell_wire[32];							inform_L[144][7] = l_cell_wire[33];							inform_L[17][7] = l_cell_wire[34];							inform_L[145][7] = l_cell_wire[35];							inform_L[18][7] = l_cell_wire[36];							inform_L[146][7] = l_cell_wire[37];							inform_L[19][7] = l_cell_wire[38];							inform_L[147][7] = l_cell_wire[39];							inform_L[20][7] = l_cell_wire[40];							inform_L[148][7] = l_cell_wire[41];							inform_L[21][7] = l_cell_wire[42];							inform_L[149][7] = l_cell_wire[43];							inform_L[22][7] = l_cell_wire[44];							inform_L[150][7] = l_cell_wire[45];							inform_L[23][7] = l_cell_wire[46];							inform_L[151][7] = l_cell_wire[47];							inform_L[24][7] = l_cell_wire[48];							inform_L[152][7] = l_cell_wire[49];							inform_L[25][7] = l_cell_wire[50];							inform_L[153][7] = l_cell_wire[51];							inform_L[26][7] = l_cell_wire[52];							inform_L[154][7] = l_cell_wire[53];							inform_L[27][7] = l_cell_wire[54];							inform_L[155][7] = l_cell_wire[55];							inform_L[28][7] = l_cell_wire[56];							inform_L[156][7] = l_cell_wire[57];							inform_L[29][7] = l_cell_wire[58];							inform_L[157][7] = l_cell_wire[59];							inform_L[30][7] = l_cell_wire[60];							inform_L[158][7] = l_cell_wire[61];							inform_L[31][7] = l_cell_wire[62];							inform_L[159][7] = l_cell_wire[63];							inform_L[32][7] = l_cell_wire[64];							inform_L[160][7] = l_cell_wire[65];							inform_L[33][7] = l_cell_wire[66];							inform_L[161][7] = l_cell_wire[67];							inform_L[34][7] = l_cell_wire[68];							inform_L[162][7] = l_cell_wire[69];							inform_L[35][7] = l_cell_wire[70];							inform_L[163][7] = l_cell_wire[71];							inform_L[36][7] = l_cell_wire[72];							inform_L[164][7] = l_cell_wire[73];							inform_L[37][7] = l_cell_wire[74];							inform_L[165][7] = l_cell_wire[75];							inform_L[38][7] = l_cell_wire[76];							inform_L[166][7] = l_cell_wire[77];							inform_L[39][7] = l_cell_wire[78];							inform_L[167][7] = l_cell_wire[79];							inform_L[40][7] = l_cell_wire[80];							inform_L[168][7] = l_cell_wire[81];							inform_L[41][7] = l_cell_wire[82];							inform_L[169][7] = l_cell_wire[83];							inform_L[42][7] = l_cell_wire[84];							inform_L[170][7] = l_cell_wire[85];							inform_L[43][7] = l_cell_wire[86];							inform_L[171][7] = l_cell_wire[87];							inform_L[44][7] = l_cell_wire[88];							inform_L[172][7] = l_cell_wire[89];							inform_L[45][7] = l_cell_wire[90];							inform_L[173][7] = l_cell_wire[91];							inform_L[46][7] = l_cell_wire[92];							inform_L[174][7] = l_cell_wire[93];							inform_L[47][7] = l_cell_wire[94];							inform_L[175][7] = l_cell_wire[95];							inform_L[48][7] = l_cell_wire[96];							inform_L[176][7] = l_cell_wire[97];							inform_L[49][7] = l_cell_wire[98];							inform_L[177][7] = l_cell_wire[99];							inform_L[50][7] = l_cell_wire[100];							inform_L[178][7] = l_cell_wire[101];							inform_L[51][7] = l_cell_wire[102];							inform_L[179][7] = l_cell_wire[103];							inform_L[52][7] = l_cell_wire[104];							inform_L[180][7] = l_cell_wire[105];							inform_L[53][7] = l_cell_wire[106];							inform_L[181][7] = l_cell_wire[107];							inform_L[54][7] = l_cell_wire[108];							inform_L[182][7] = l_cell_wire[109];							inform_L[55][7] = l_cell_wire[110];							inform_L[183][7] = l_cell_wire[111];							inform_L[56][7] = l_cell_wire[112];							inform_L[184][7] = l_cell_wire[113];							inform_L[57][7] = l_cell_wire[114];							inform_L[185][7] = l_cell_wire[115];							inform_L[58][7] = l_cell_wire[116];							inform_L[186][7] = l_cell_wire[117];							inform_L[59][7] = l_cell_wire[118];							inform_L[187][7] = l_cell_wire[119];							inform_L[60][7] = l_cell_wire[120];							inform_L[188][7] = l_cell_wire[121];							inform_L[61][7] = l_cell_wire[122];							inform_L[189][7] = l_cell_wire[123];							inform_L[62][7] = l_cell_wire[124];							inform_L[190][7] = l_cell_wire[125];							inform_L[63][7] = l_cell_wire[126];							inform_L[191][7] = l_cell_wire[127];							inform_L[64][7] = l_cell_wire[128];							inform_L[192][7] = l_cell_wire[129];							inform_L[65][7] = l_cell_wire[130];							inform_L[193][7] = l_cell_wire[131];							inform_L[66][7] = l_cell_wire[132];							inform_L[194][7] = l_cell_wire[133];							inform_L[67][7] = l_cell_wire[134];							inform_L[195][7] = l_cell_wire[135];							inform_L[68][7] = l_cell_wire[136];							inform_L[196][7] = l_cell_wire[137];							inform_L[69][7] = l_cell_wire[138];							inform_L[197][7] = l_cell_wire[139];							inform_L[70][7] = l_cell_wire[140];							inform_L[198][7] = l_cell_wire[141];							inform_L[71][7] = l_cell_wire[142];							inform_L[199][7] = l_cell_wire[143];							inform_L[72][7] = l_cell_wire[144];							inform_L[200][7] = l_cell_wire[145];							inform_L[73][7] = l_cell_wire[146];							inform_L[201][7] = l_cell_wire[147];							inform_L[74][7] = l_cell_wire[148];							inform_L[202][7] = l_cell_wire[149];							inform_L[75][7] = l_cell_wire[150];							inform_L[203][7] = l_cell_wire[151];							inform_L[76][7] = l_cell_wire[152];							inform_L[204][7] = l_cell_wire[153];							inform_L[77][7] = l_cell_wire[154];							inform_L[205][7] = l_cell_wire[155];							inform_L[78][7] = l_cell_wire[156];							inform_L[206][7] = l_cell_wire[157];							inform_L[79][7] = l_cell_wire[158];							inform_L[207][7] = l_cell_wire[159];							inform_L[80][7] = l_cell_wire[160];							inform_L[208][7] = l_cell_wire[161];							inform_L[81][7] = l_cell_wire[162];							inform_L[209][7] = l_cell_wire[163];							inform_L[82][7] = l_cell_wire[164];							inform_L[210][7] = l_cell_wire[165];							inform_L[83][7] = l_cell_wire[166];							inform_L[211][7] = l_cell_wire[167];							inform_L[84][7] = l_cell_wire[168];							inform_L[212][7] = l_cell_wire[169];							inform_L[85][7] = l_cell_wire[170];							inform_L[213][7] = l_cell_wire[171];							inform_L[86][7] = l_cell_wire[172];							inform_L[214][7] = l_cell_wire[173];							inform_L[87][7] = l_cell_wire[174];							inform_L[215][7] = l_cell_wire[175];							inform_L[88][7] = l_cell_wire[176];							inform_L[216][7] = l_cell_wire[177];							inform_L[89][7] = l_cell_wire[178];							inform_L[217][7] = l_cell_wire[179];							inform_L[90][7] = l_cell_wire[180];							inform_L[218][7] = l_cell_wire[181];							inform_L[91][7] = l_cell_wire[182];							inform_L[219][7] = l_cell_wire[183];							inform_L[92][7] = l_cell_wire[184];							inform_L[220][7] = l_cell_wire[185];							inform_L[93][7] = l_cell_wire[186];							inform_L[221][7] = l_cell_wire[187];							inform_L[94][7] = l_cell_wire[188];							inform_L[222][7] = l_cell_wire[189];							inform_L[95][7] = l_cell_wire[190];							inform_L[223][7] = l_cell_wire[191];							inform_L[96][7] = l_cell_wire[192];							inform_L[224][7] = l_cell_wire[193];							inform_L[97][7] = l_cell_wire[194];							inform_L[225][7] = l_cell_wire[195];							inform_L[98][7] = l_cell_wire[196];							inform_L[226][7] = l_cell_wire[197];							inform_L[99][7] = l_cell_wire[198];							inform_L[227][7] = l_cell_wire[199];							inform_L[100][7] = l_cell_wire[200];							inform_L[228][7] = l_cell_wire[201];							inform_L[101][7] = l_cell_wire[202];							inform_L[229][7] = l_cell_wire[203];							inform_L[102][7] = l_cell_wire[204];							inform_L[230][7] = l_cell_wire[205];							inform_L[103][7] = l_cell_wire[206];							inform_L[231][7] = l_cell_wire[207];							inform_L[104][7] = l_cell_wire[208];							inform_L[232][7] = l_cell_wire[209];							inform_L[105][7] = l_cell_wire[210];							inform_L[233][7] = l_cell_wire[211];							inform_L[106][7] = l_cell_wire[212];							inform_L[234][7] = l_cell_wire[213];							inform_L[107][7] = l_cell_wire[214];							inform_L[235][7] = l_cell_wire[215];							inform_L[108][7] = l_cell_wire[216];							inform_L[236][7] = l_cell_wire[217];							inform_L[109][7] = l_cell_wire[218];							inform_L[237][7] = l_cell_wire[219];							inform_L[110][7] = l_cell_wire[220];							inform_L[238][7] = l_cell_wire[221];							inform_L[111][7] = l_cell_wire[222];							inform_L[239][7] = l_cell_wire[223];							inform_L[112][7] = l_cell_wire[224];							inform_L[240][7] = l_cell_wire[225];							inform_L[113][7] = l_cell_wire[226];							inform_L[241][7] = l_cell_wire[227];							inform_L[114][7] = l_cell_wire[228];							inform_L[242][7] = l_cell_wire[229];							inform_L[115][7] = l_cell_wire[230];							inform_L[243][7] = l_cell_wire[231];							inform_L[116][7] = l_cell_wire[232];							inform_L[244][7] = l_cell_wire[233];							inform_L[117][7] = l_cell_wire[234];							inform_L[245][7] = l_cell_wire[235];							inform_L[118][7] = l_cell_wire[236];							inform_L[246][7] = l_cell_wire[237];							inform_L[119][7] = l_cell_wire[238];							inform_L[247][7] = l_cell_wire[239];							inform_L[120][7] = l_cell_wire[240];							inform_L[248][7] = l_cell_wire[241];							inform_L[121][7] = l_cell_wire[242];							inform_L[249][7] = l_cell_wire[243];							inform_L[122][7] = l_cell_wire[244];							inform_L[250][7] = l_cell_wire[245];							inform_L[123][7] = l_cell_wire[246];							inform_L[251][7] = l_cell_wire[247];							inform_L[124][7] = l_cell_wire[248];							inform_L[252][7] = l_cell_wire[249];							inform_L[125][7] = l_cell_wire[250];							inform_L[253][7] = l_cell_wire[251];							inform_L[126][7] = l_cell_wire[252];							inform_L[254][7] = l_cell_wire[253];							inform_L[127][7] = l_cell_wire[254];							inform_L[255][7] = l_cell_wire[255];							inform_L[256][7] = l_cell_wire[256];							inform_L[384][7] = l_cell_wire[257];							inform_L[257][7] = l_cell_wire[258];							inform_L[385][7] = l_cell_wire[259];							inform_L[258][7] = l_cell_wire[260];							inform_L[386][7] = l_cell_wire[261];							inform_L[259][7] = l_cell_wire[262];							inform_L[387][7] = l_cell_wire[263];							inform_L[260][7] = l_cell_wire[264];							inform_L[388][7] = l_cell_wire[265];							inform_L[261][7] = l_cell_wire[266];							inform_L[389][7] = l_cell_wire[267];							inform_L[262][7] = l_cell_wire[268];							inform_L[390][7] = l_cell_wire[269];							inform_L[263][7] = l_cell_wire[270];							inform_L[391][7] = l_cell_wire[271];							inform_L[264][7] = l_cell_wire[272];							inform_L[392][7] = l_cell_wire[273];							inform_L[265][7] = l_cell_wire[274];							inform_L[393][7] = l_cell_wire[275];							inform_L[266][7] = l_cell_wire[276];							inform_L[394][7] = l_cell_wire[277];							inform_L[267][7] = l_cell_wire[278];							inform_L[395][7] = l_cell_wire[279];							inform_L[268][7] = l_cell_wire[280];							inform_L[396][7] = l_cell_wire[281];							inform_L[269][7] = l_cell_wire[282];							inform_L[397][7] = l_cell_wire[283];							inform_L[270][7] = l_cell_wire[284];							inform_L[398][7] = l_cell_wire[285];							inform_L[271][7] = l_cell_wire[286];							inform_L[399][7] = l_cell_wire[287];							inform_L[272][7] = l_cell_wire[288];							inform_L[400][7] = l_cell_wire[289];							inform_L[273][7] = l_cell_wire[290];							inform_L[401][7] = l_cell_wire[291];							inform_L[274][7] = l_cell_wire[292];							inform_L[402][7] = l_cell_wire[293];							inform_L[275][7] = l_cell_wire[294];							inform_L[403][7] = l_cell_wire[295];							inform_L[276][7] = l_cell_wire[296];							inform_L[404][7] = l_cell_wire[297];							inform_L[277][7] = l_cell_wire[298];							inform_L[405][7] = l_cell_wire[299];							inform_L[278][7] = l_cell_wire[300];							inform_L[406][7] = l_cell_wire[301];							inform_L[279][7] = l_cell_wire[302];							inform_L[407][7] = l_cell_wire[303];							inform_L[280][7] = l_cell_wire[304];							inform_L[408][7] = l_cell_wire[305];							inform_L[281][7] = l_cell_wire[306];							inform_L[409][7] = l_cell_wire[307];							inform_L[282][7] = l_cell_wire[308];							inform_L[410][7] = l_cell_wire[309];							inform_L[283][7] = l_cell_wire[310];							inform_L[411][7] = l_cell_wire[311];							inform_L[284][7] = l_cell_wire[312];							inform_L[412][7] = l_cell_wire[313];							inform_L[285][7] = l_cell_wire[314];							inform_L[413][7] = l_cell_wire[315];							inform_L[286][7] = l_cell_wire[316];							inform_L[414][7] = l_cell_wire[317];							inform_L[287][7] = l_cell_wire[318];							inform_L[415][7] = l_cell_wire[319];							inform_L[288][7] = l_cell_wire[320];							inform_L[416][7] = l_cell_wire[321];							inform_L[289][7] = l_cell_wire[322];							inform_L[417][7] = l_cell_wire[323];							inform_L[290][7] = l_cell_wire[324];							inform_L[418][7] = l_cell_wire[325];							inform_L[291][7] = l_cell_wire[326];							inform_L[419][7] = l_cell_wire[327];							inform_L[292][7] = l_cell_wire[328];							inform_L[420][7] = l_cell_wire[329];							inform_L[293][7] = l_cell_wire[330];							inform_L[421][7] = l_cell_wire[331];							inform_L[294][7] = l_cell_wire[332];							inform_L[422][7] = l_cell_wire[333];							inform_L[295][7] = l_cell_wire[334];							inform_L[423][7] = l_cell_wire[335];							inform_L[296][7] = l_cell_wire[336];							inform_L[424][7] = l_cell_wire[337];							inform_L[297][7] = l_cell_wire[338];							inform_L[425][7] = l_cell_wire[339];							inform_L[298][7] = l_cell_wire[340];							inform_L[426][7] = l_cell_wire[341];							inform_L[299][7] = l_cell_wire[342];							inform_L[427][7] = l_cell_wire[343];							inform_L[300][7] = l_cell_wire[344];							inform_L[428][7] = l_cell_wire[345];							inform_L[301][7] = l_cell_wire[346];							inform_L[429][7] = l_cell_wire[347];							inform_L[302][7] = l_cell_wire[348];							inform_L[430][7] = l_cell_wire[349];							inform_L[303][7] = l_cell_wire[350];							inform_L[431][7] = l_cell_wire[351];							inform_L[304][7] = l_cell_wire[352];							inform_L[432][7] = l_cell_wire[353];							inform_L[305][7] = l_cell_wire[354];							inform_L[433][7] = l_cell_wire[355];							inform_L[306][7] = l_cell_wire[356];							inform_L[434][7] = l_cell_wire[357];							inform_L[307][7] = l_cell_wire[358];							inform_L[435][7] = l_cell_wire[359];							inform_L[308][7] = l_cell_wire[360];							inform_L[436][7] = l_cell_wire[361];							inform_L[309][7] = l_cell_wire[362];							inform_L[437][7] = l_cell_wire[363];							inform_L[310][7] = l_cell_wire[364];							inform_L[438][7] = l_cell_wire[365];							inform_L[311][7] = l_cell_wire[366];							inform_L[439][7] = l_cell_wire[367];							inform_L[312][7] = l_cell_wire[368];							inform_L[440][7] = l_cell_wire[369];							inform_L[313][7] = l_cell_wire[370];							inform_L[441][7] = l_cell_wire[371];							inform_L[314][7] = l_cell_wire[372];							inform_L[442][7] = l_cell_wire[373];							inform_L[315][7] = l_cell_wire[374];							inform_L[443][7] = l_cell_wire[375];							inform_L[316][7] = l_cell_wire[376];							inform_L[444][7] = l_cell_wire[377];							inform_L[317][7] = l_cell_wire[378];							inform_L[445][7] = l_cell_wire[379];							inform_L[318][7] = l_cell_wire[380];							inform_L[446][7] = l_cell_wire[381];							inform_L[319][7] = l_cell_wire[382];							inform_L[447][7] = l_cell_wire[383];							inform_L[320][7] = l_cell_wire[384];							inform_L[448][7] = l_cell_wire[385];							inform_L[321][7] = l_cell_wire[386];							inform_L[449][7] = l_cell_wire[387];							inform_L[322][7] = l_cell_wire[388];							inform_L[450][7] = l_cell_wire[389];							inform_L[323][7] = l_cell_wire[390];							inform_L[451][7] = l_cell_wire[391];							inform_L[324][7] = l_cell_wire[392];							inform_L[452][7] = l_cell_wire[393];							inform_L[325][7] = l_cell_wire[394];							inform_L[453][7] = l_cell_wire[395];							inform_L[326][7] = l_cell_wire[396];							inform_L[454][7] = l_cell_wire[397];							inform_L[327][7] = l_cell_wire[398];							inform_L[455][7] = l_cell_wire[399];							inform_L[328][7] = l_cell_wire[400];							inform_L[456][7] = l_cell_wire[401];							inform_L[329][7] = l_cell_wire[402];							inform_L[457][7] = l_cell_wire[403];							inform_L[330][7] = l_cell_wire[404];							inform_L[458][7] = l_cell_wire[405];							inform_L[331][7] = l_cell_wire[406];							inform_L[459][7] = l_cell_wire[407];							inform_L[332][7] = l_cell_wire[408];							inform_L[460][7] = l_cell_wire[409];							inform_L[333][7] = l_cell_wire[410];							inform_L[461][7] = l_cell_wire[411];							inform_L[334][7] = l_cell_wire[412];							inform_L[462][7] = l_cell_wire[413];							inform_L[335][7] = l_cell_wire[414];							inform_L[463][7] = l_cell_wire[415];							inform_L[336][7] = l_cell_wire[416];							inform_L[464][7] = l_cell_wire[417];							inform_L[337][7] = l_cell_wire[418];							inform_L[465][7] = l_cell_wire[419];							inform_L[338][7] = l_cell_wire[420];							inform_L[466][7] = l_cell_wire[421];							inform_L[339][7] = l_cell_wire[422];							inform_L[467][7] = l_cell_wire[423];							inform_L[340][7] = l_cell_wire[424];							inform_L[468][7] = l_cell_wire[425];							inform_L[341][7] = l_cell_wire[426];							inform_L[469][7] = l_cell_wire[427];							inform_L[342][7] = l_cell_wire[428];							inform_L[470][7] = l_cell_wire[429];							inform_L[343][7] = l_cell_wire[430];							inform_L[471][7] = l_cell_wire[431];							inform_L[344][7] = l_cell_wire[432];							inform_L[472][7] = l_cell_wire[433];							inform_L[345][7] = l_cell_wire[434];							inform_L[473][7] = l_cell_wire[435];							inform_L[346][7] = l_cell_wire[436];							inform_L[474][7] = l_cell_wire[437];							inform_L[347][7] = l_cell_wire[438];							inform_L[475][7] = l_cell_wire[439];							inform_L[348][7] = l_cell_wire[440];							inform_L[476][7] = l_cell_wire[441];							inform_L[349][7] = l_cell_wire[442];							inform_L[477][7] = l_cell_wire[443];							inform_L[350][7] = l_cell_wire[444];							inform_L[478][7] = l_cell_wire[445];							inform_L[351][7] = l_cell_wire[446];							inform_L[479][7] = l_cell_wire[447];							inform_L[352][7] = l_cell_wire[448];							inform_L[480][7] = l_cell_wire[449];							inform_L[353][7] = l_cell_wire[450];							inform_L[481][7] = l_cell_wire[451];							inform_L[354][7] = l_cell_wire[452];							inform_L[482][7] = l_cell_wire[453];							inform_L[355][7] = l_cell_wire[454];							inform_L[483][7] = l_cell_wire[455];							inform_L[356][7] = l_cell_wire[456];							inform_L[484][7] = l_cell_wire[457];							inform_L[357][7] = l_cell_wire[458];							inform_L[485][7] = l_cell_wire[459];							inform_L[358][7] = l_cell_wire[460];							inform_L[486][7] = l_cell_wire[461];							inform_L[359][7] = l_cell_wire[462];							inform_L[487][7] = l_cell_wire[463];							inform_L[360][7] = l_cell_wire[464];							inform_L[488][7] = l_cell_wire[465];							inform_L[361][7] = l_cell_wire[466];							inform_L[489][7] = l_cell_wire[467];							inform_L[362][7] = l_cell_wire[468];							inform_L[490][7] = l_cell_wire[469];							inform_L[363][7] = l_cell_wire[470];							inform_L[491][7] = l_cell_wire[471];							inform_L[364][7] = l_cell_wire[472];							inform_L[492][7] = l_cell_wire[473];							inform_L[365][7] = l_cell_wire[474];							inform_L[493][7] = l_cell_wire[475];							inform_L[366][7] = l_cell_wire[476];							inform_L[494][7] = l_cell_wire[477];							inform_L[367][7] = l_cell_wire[478];							inform_L[495][7] = l_cell_wire[479];							inform_L[368][7] = l_cell_wire[480];							inform_L[496][7] = l_cell_wire[481];							inform_L[369][7] = l_cell_wire[482];							inform_L[497][7] = l_cell_wire[483];							inform_L[370][7] = l_cell_wire[484];							inform_L[498][7] = l_cell_wire[485];							inform_L[371][7] = l_cell_wire[486];							inform_L[499][7] = l_cell_wire[487];							inform_L[372][7] = l_cell_wire[488];							inform_L[500][7] = l_cell_wire[489];							inform_L[373][7] = l_cell_wire[490];							inform_L[501][7] = l_cell_wire[491];							inform_L[374][7] = l_cell_wire[492];							inform_L[502][7] = l_cell_wire[493];							inform_L[375][7] = l_cell_wire[494];							inform_L[503][7] = l_cell_wire[495];							inform_L[376][7] = l_cell_wire[496];							inform_L[504][7] = l_cell_wire[497];							inform_L[377][7] = l_cell_wire[498];							inform_L[505][7] = l_cell_wire[499];							inform_L[378][7] = l_cell_wire[500];							inform_L[506][7] = l_cell_wire[501];							inform_L[379][7] = l_cell_wire[502];							inform_L[507][7] = l_cell_wire[503];							inform_L[380][7] = l_cell_wire[504];							inform_L[508][7] = l_cell_wire[505];							inform_L[381][7] = l_cell_wire[506];							inform_L[509][7] = l_cell_wire[507];							inform_L[382][7] = l_cell_wire[508];							inform_L[510][7] = l_cell_wire[509];							inform_L[383][7] = l_cell_wire[510];							inform_L[511][7] = l_cell_wire[511];							inform_L[512][7] = l_cell_wire[512];							inform_L[640][7] = l_cell_wire[513];							inform_L[513][7] = l_cell_wire[514];							inform_L[641][7] = l_cell_wire[515];							inform_L[514][7] = l_cell_wire[516];							inform_L[642][7] = l_cell_wire[517];							inform_L[515][7] = l_cell_wire[518];							inform_L[643][7] = l_cell_wire[519];							inform_L[516][7] = l_cell_wire[520];							inform_L[644][7] = l_cell_wire[521];							inform_L[517][7] = l_cell_wire[522];							inform_L[645][7] = l_cell_wire[523];							inform_L[518][7] = l_cell_wire[524];							inform_L[646][7] = l_cell_wire[525];							inform_L[519][7] = l_cell_wire[526];							inform_L[647][7] = l_cell_wire[527];							inform_L[520][7] = l_cell_wire[528];							inform_L[648][7] = l_cell_wire[529];							inform_L[521][7] = l_cell_wire[530];							inform_L[649][7] = l_cell_wire[531];							inform_L[522][7] = l_cell_wire[532];							inform_L[650][7] = l_cell_wire[533];							inform_L[523][7] = l_cell_wire[534];							inform_L[651][7] = l_cell_wire[535];							inform_L[524][7] = l_cell_wire[536];							inform_L[652][7] = l_cell_wire[537];							inform_L[525][7] = l_cell_wire[538];							inform_L[653][7] = l_cell_wire[539];							inform_L[526][7] = l_cell_wire[540];							inform_L[654][7] = l_cell_wire[541];							inform_L[527][7] = l_cell_wire[542];							inform_L[655][7] = l_cell_wire[543];							inform_L[528][7] = l_cell_wire[544];							inform_L[656][7] = l_cell_wire[545];							inform_L[529][7] = l_cell_wire[546];							inform_L[657][7] = l_cell_wire[547];							inform_L[530][7] = l_cell_wire[548];							inform_L[658][7] = l_cell_wire[549];							inform_L[531][7] = l_cell_wire[550];							inform_L[659][7] = l_cell_wire[551];							inform_L[532][7] = l_cell_wire[552];							inform_L[660][7] = l_cell_wire[553];							inform_L[533][7] = l_cell_wire[554];							inform_L[661][7] = l_cell_wire[555];							inform_L[534][7] = l_cell_wire[556];							inform_L[662][7] = l_cell_wire[557];							inform_L[535][7] = l_cell_wire[558];							inform_L[663][7] = l_cell_wire[559];							inform_L[536][7] = l_cell_wire[560];							inform_L[664][7] = l_cell_wire[561];							inform_L[537][7] = l_cell_wire[562];							inform_L[665][7] = l_cell_wire[563];							inform_L[538][7] = l_cell_wire[564];							inform_L[666][7] = l_cell_wire[565];							inform_L[539][7] = l_cell_wire[566];							inform_L[667][7] = l_cell_wire[567];							inform_L[540][7] = l_cell_wire[568];							inform_L[668][7] = l_cell_wire[569];							inform_L[541][7] = l_cell_wire[570];							inform_L[669][7] = l_cell_wire[571];							inform_L[542][7] = l_cell_wire[572];							inform_L[670][7] = l_cell_wire[573];							inform_L[543][7] = l_cell_wire[574];							inform_L[671][7] = l_cell_wire[575];							inform_L[544][7] = l_cell_wire[576];							inform_L[672][7] = l_cell_wire[577];							inform_L[545][7] = l_cell_wire[578];							inform_L[673][7] = l_cell_wire[579];							inform_L[546][7] = l_cell_wire[580];							inform_L[674][7] = l_cell_wire[581];							inform_L[547][7] = l_cell_wire[582];							inform_L[675][7] = l_cell_wire[583];							inform_L[548][7] = l_cell_wire[584];							inform_L[676][7] = l_cell_wire[585];							inform_L[549][7] = l_cell_wire[586];							inform_L[677][7] = l_cell_wire[587];							inform_L[550][7] = l_cell_wire[588];							inform_L[678][7] = l_cell_wire[589];							inform_L[551][7] = l_cell_wire[590];							inform_L[679][7] = l_cell_wire[591];							inform_L[552][7] = l_cell_wire[592];							inform_L[680][7] = l_cell_wire[593];							inform_L[553][7] = l_cell_wire[594];							inform_L[681][7] = l_cell_wire[595];							inform_L[554][7] = l_cell_wire[596];							inform_L[682][7] = l_cell_wire[597];							inform_L[555][7] = l_cell_wire[598];							inform_L[683][7] = l_cell_wire[599];							inform_L[556][7] = l_cell_wire[600];							inform_L[684][7] = l_cell_wire[601];							inform_L[557][7] = l_cell_wire[602];							inform_L[685][7] = l_cell_wire[603];							inform_L[558][7] = l_cell_wire[604];							inform_L[686][7] = l_cell_wire[605];							inform_L[559][7] = l_cell_wire[606];							inform_L[687][7] = l_cell_wire[607];							inform_L[560][7] = l_cell_wire[608];							inform_L[688][7] = l_cell_wire[609];							inform_L[561][7] = l_cell_wire[610];							inform_L[689][7] = l_cell_wire[611];							inform_L[562][7] = l_cell_wire[612];							inform_L[690][7] = l_cell_wire[613];							inform_L[563][7] = l_cell_wire[614];							inform_L[691][7] = l_cell_wire[615];							inform_L[564][7] = l_cell_wire[616];							inform_L[692][7] = l_cell_wire[617];							inform_L[565][7] = l_cell_wire[618];							inform_L[693][7] = l_cell_wire[619];							inform_L[566][7] = l_cell_wire[620];							inform_L[694][7] = l_cell_wire[621];							inform_L[567][7] = l_cell_wire[622];							inform_L[695][7] = l_cell_wire[623];							inform_L[568][7] = l_cell_wire[624];							inform_L[696][7] = l_cell_wire[625];							inform_L[569][7] = l_cell_wire[626];							inform_L[697][7] = l_cell_wire[627];							inform_L[570][7] = l_cell_wire[628];							inform_L[698][7] = l_cell_wire[629];							inform_L[571][7] = l_cell_wire[630];							inform_L[699][7] = l_cell_wire[631];							inform_L[572][7] = l_cell_wire[632];							inform_L[700][7] = l_cell_wire[633];							inform_L[573][7] = l_cell_wire[634];							inform_L[701][7] = l_cell_wire[635];							inform_L[574][7] = l_cell_wire[636];							inform_L[702][7] = l_cell_wire[637];							inform_L[575][7] = l_cell_wire[638];							inform_L[703][7] = l_cell_wire[639];							inform_L[576][7] = l_cell_wire[640];							inform_L[704][7] = l_cell_wire[641];							inform_L[577][7] = l_cell_wire[642];							inform_L[705][7] = l_cell_wire[643];							inform_L[578][7] = l_cell_wire[644];							inform_L[706][7] = l_cell_wire[645];							inform_L[579][7] = l_cell_wire[646];							inform_L[707][7] = l_cell_wire[647];							inform_L[580][7] = l_cell_wire[648];							inform_L[708][7] = l_cell_wire[649];							inform_L[581][7] = l_cell_wire[650];							inform_L[709][7] = l_cell_wire[651];							inform_L[582][7] = l_cell_wire[652];							inform_L[710][7] = l_cell_wire[653];							inform_L[583][7] = l_cell_wire[654];							inform_L[711][7] = l_cell_wire[655];							inform_L[584][7] = l_cell_wire[656];							inform_L[712][7] = l_cell_wire[657];							inform_L[585][7] = l_cell_wire[658];							inform_L[713][7] = l_cell_wire[659];							inform_L[586][7] = l_cell_wire[660];							inform_L[714][7] = l_cell_wire[661];							inform_L[587][7] = l_cell_wire[662];							inform_L[715][7] = l_cell_wire[663];							inform_L[588][7] = l_cell_wire[664];							inform_L[716][7] = l_cell_wire[665];							inform_L[589][7] = l_cell_wire[666];							inform_L[717][7] = l_cell_wire[667];							inform_L[590][7] = l_cell_wire[668];							inform_L[718][7] = l_cell_wire[669];							inform_L[591][7] = l_cell_wire[670];							inform_L[719][7] = l_cell_wire[671];							inform_L[592][7] = l_cell_wire[672];							inform_L[720][7] = l_cell_wire[673];							inform_L[593][7] = l_cell_wire[674];							inform_L[721][7] = l_cell_wire[675];							inform_L[594][7] = l_cell_wire[676];							inform_L[722][7] = l_cell_wire[677];							inform_L[595][7] = l_cell_wire[678];							inform_L[723][7] = l_cell_wire[679];							inform_L[596][7] = l_cell_wire[680];							inform_L[724][7] = l_cell_wire[681];							inform_L[597][7] = l_cell_wire[682];							inform_L[725][7] = l_cell_wire[683];							inform_L[598][7] = l_cell_wire[684];							inform_L[726][7] = l_cell_wire[685];							inform_L[599][7] = l_cell_wire[686];							inform_L[727][7] = l_cell_wire[687];							inform_L[600][7] = l_cell_wire[688];							inform_L[728][7] = l_cell_wire[689];							inform_L[601][7] = l_cell_wire[690];							inform_L[729][7] = l_cell_wire[691];							inform_L[602][7] = l_cell_wire[692];							inform_L[730][7] = l_cell_wire[693];							inform_L[603][7] = l_cell_wire[694];							inform_L[731][7] = l_cell_wire[695];							inform_L[604][7] = l_cell_wire[696];							inform_L[732][7] = l_cell_wire[697];							inform_L[605][7] = l_cell_wire[698];							inform_L[733][7] = l_cell_wire[699];							inform_L[606][7] = l_cell_wire[700];							inform_L[734][7] = l_cell_wire[701];							inform_L[607][7] = l_cell_wire[702];							inform_L[735][7] = l_cell_wire[703];							inform_L[608][7] = l_cell_wire[704];							inform_L[736][7] = l_cell_wire[705];							inform_L[609][7] = l_cell_wire[706];							inform_L[737][7] = l_cell_wire[707];							inform_L[610][7] = l_cell_wire[708];							inform_L[738][7] = l_cell_wire[709];							inform_L[611][7] = l_cell_wire[710];							inform_L[739][7] = l_cell_wire[711];							inform_L[612][7] = l_cell_wire[712];							inform_L[740][7] = l_cell_wire[713];							inform_L[613][7] = l_cell_wire[714];							inform_L[741][7] = l_cell_wire[715];							inform_L[614][7] = l_cell_wire[716];							inform_L[742][7] = l_cell_wire[717];							inform_L[615][7] = l_cell_wire[718];							inform_L[743][7] = l_cell_wire[719];							inform_L[616][7] = l_cell_wire[720];							inform_L[744][7] = l_cell_wire[721];							inform_L[617][7] = l_cell_wire[722];							inform_L[745][7] = l_cell_wire[723];							inform_L[618][7] = l_cell_wire[724];							inform_L[746][7] = l_cell_wire[725];							inform_L[619][7] = l_cell_wire[726];							inform_L[747][7] = l_cell_wire[727];							inform_L[620][7] = l_cell_wire[728];							inform_L[748][7] = l_cell_wire[729];							inform_L[621][7] = l_cell_wire[730];							inform_L[749][7] = l_cell_wire[731];							inform_L[622][7] = l_cell_wire[732];							inform_L[750][7] = l_cell_wire[733];							inform_L[623][7] = l_cell_wire[734];							inform_L[751][7] = l_cell_wire[735];							inform_L[624][7] = l_cell_wire[736];							inform_L[752][7] = l_cell_wire[737];							inform_L[625][7] = l_cell_wire[738];							inform_L[753][7] = l_cell_wire[739];							inform_L[626][7] = l_cell_wire[740];							inform_L[754][7] = l_cell_wire[741];							inform_L[627][7] = l_cell_wire[742];							inform_L[755][7] = l_cell_wire[743];							inform_L[628][7] = l_cell_wire[744];							inform_L[756][7] = l_cell_wire[745];							inform_L[629][7] = l_cell_wire[746];							inform_L[757][7] = l_cell_wire[747];							inform_L[630][7] = l_cell_wire[748];							inform_L[758][7] = l_cell_wire[749];							inform_L[631][7] = l_cell_wire[750];							inform_L[759][7] = l_cell_wire[751];							inform_L[632][7] = l_cell_wire[752];							inform_L[760][7] = l_cell_wire[753];							inform_L[633][7] = l_cell_wire[754];							inform_L[761][7] = l_cell_wire[755];							inform_L[634][7] = l_cell_wire[756];							inform_L[762][7] = l_cell_wire[757];							inform_L[635][7] = l_cell_wire[758];							inform_L[763][7] = l_cell_wire[759];							inform_L[636][7] = l_cell_wire[760];							inform_L[764][7] = l_cell_wire[761];							inform_L[637][7] = l_cell_wire[762];							inform_L[765][7] = l_cell_wire[763];							inform_L[638][7] = l_cell_wire[764];							inform_L[766][7] = l_cell_wire[765];							inform_L[639][7] = l_cell_wire[766];							inform_L[767][7] = l_cell_wire[767];							inform_L[768][7] = l_cell_wire[768];							inform_L[896][7] = l_cell_wire[769];							inform_L[769][7] = l_cell_wire[770];							inform_L[897][7] = l_cell_wire[771];							inform_L[770][7] = l_cell_wire[772];							inform_L[898][7] = l_cell_wire[773];							inform_L[771][7] = l_cell_wire[774];							inform_L[899][7] = l_cell_wire[775];							inform_L[772][7] = l_cell_wire[776];							inform_L[900][7] = l_cell_wire[777];							inform_L[773][7] = l_cell_wire[778];							inform_L[901][7] = l_cell_wire[779];							inform_L[774][7] = l_cell_wire[780];							inform_L[902][7] = l_cell_wire[781];							inform_L[775][7] = l_cell_wire[782];							inform_L[903][7] = l_cell_wire[783];							inform_L[776][7] = l_cell_wire[784];							inform_L[904][7] = l_cell_wire[785];							inform_L[777][7] = l_cell_wire[786];							inform_L[905][7] = l_cell_wire[787];							inform_L[778][7] = l_cell_wire[788];							inform_L[906][7] = l_cell_wire[789];							inform_L[779][7] = l_cell_wire[790];							inform_L[907][7] = l_cell_wire[791];							inform_L[780][7] = l_cell_wire[792];							inform_L[908][7] = l_cell_wire[793];							inform_L[781][7] = l_cell_wire[794];							inform_L[909][7] = l_cell_wire[795];							inform_L[782][7] = l_cell_wire[796];							inform_L[910][7] = l_cell_wire[797];							inform_L[783][7] = l_cell_wire[798];							inform_L[911][7] = l_cell_wire[799];							inform_L[784][7] = l_cell_wire[800];							inform_L[912][7] = l_cell_wire[801];							inform_L[785][7] = l_cell_wire[802];							inform_L[913][7] = l_cell_wire[803];							inform_L[786][7] = l_cell_wire[804];							inform_L[914][7] = l_cell_wire[805];							inform_L[787][7] = l_cell_wire[806];							inform_L[915][7] = l_cell_wire[807];							inform_L[788][7] = l_cell_wire[808];							inform_L[916][7] = l_cell_wire[809];							inform_L[789][7] = l_cell_wire[810];							inform_L[917][7] = l_cell_wire[811];							inform_L[790][7] = l_cell_wire[812];							inform_L[918][7] = l_cell_wire[813];							inform_L[791][7] = l_cell_wire[814];							inform_L[919][7] = l_cell_wire[815];							inform_L[792][7] = l_cell_wire[816];							inform_L[920][7] = l_cell_wire[817];							inform_L[793][7] = l_cell_wire[818];							inform_L[921][7] = l_cell_wire[819];							inform_L[794][7] = l_cell_wire[820];							inform_L[922][7] = l_cell_wire[821];							inform_L[795][7] = l_cell_wire[822];							inform_L[923][7] = l_cell_wire[823];							inform_L[796][7] = l_cell_wire[824];							inform_L[924][7] = l_cell_wire[825];							inform_L[797][7] = l_cell_wire[826];							inform_L[925][7] = l_cell_wire[827];							inform_L[798][7] = l_cell_wire[828];							inform_L[926][7] = l_cell_wire[829];							inform_L[799][7] = l_cell_wire[830];							inform_L[927][7] = l_cell_wire[831];							inform_L[800][7] = l_cell_wire[832];							inform_L[928][7] = l_cell_wire[833];							inform_L[801][7] = l_cell_wire[834];							inform_L[929][7] = l_cell_wire[835];							inform_L[802][7] = l_cell_wire[836];							inform_L[930][7] = l_cell_wire[837];							inform_L[803][7] = l_cell_wire[838];							inform_L[931][7] = l_cell_wire[839];							inform_L[804][7] = l_cell_wire[840];							inform_L[932][7] = l_cell_wire[841];							inform_L[805][7] = l_cell_wire[842];							inform_L[933][7] = l_cell_wire[843];							inform_L[806][7] = l_cell_wire[844];							inform_L[934][7] = l_cell_wire[845];							inform_L[807][7] = l_cell_wire[846];							inform_L[935][7] = l_cell_wire[847];							inform_L[808][7] = l_cell_wire[848];							inform_L[936][7] = l_cell_wire[849];							inform_L[809][7] = l_cell_wire[850];							inform_L[937][7] = l_cell_wire[851];							inform_L[810][7] = l_cell_wire[852];							inform_L[938][7] = l_cell_wire[853];							inform_L[811][7] = l_cell_wire[854];							inform_L[939][7] = l_cell_wire[855];							inform_L[812][7] = l_cell_wire[856];							inform_L[940][7] = l_cell_wire[857];							inform_L[813][7] = l_cell_wire[858];							inform_L[941][7] = l_cell_wire[859];							inform_L[814][7] = l_cell_wire[860];							inform_L[942][7] = l_cell_wire[861];							inform_L[815][7] = l_cell_wire[862];							inform_L[943][7] = l_cell_wire[863];							inform_L[816][7] = l_cell_wire[864];							inform_L[944][7] = l_cell_wire[865];							inform_L[817][7] = l_cell_wire[866];							inform_L[945][7] = l_cell_wire[867];							inform_L[818][7] = l_cell_wire[868];							inform_L[946][7] = l_cell_wire[869];							inform_L[819][7] = l_cell_wire[870];							inform_L[947][7] = l_cell_wire[871];							inform_L[820][7] = l_cell_wire[872];							inform_L[948][7] = l_cell_wire[873];							inform_L[821][7] = l_cell_wire[874];							inform_L[949][7] = l_cell_wire[875];							inform_L[822][7] = l_cell_wire[876];							inform_L[950][7] = l_cell_wire[877];							inform_L[823][7] = l_cell_wire[878];							inform_L[951][7] = l_cell_wire[879];							inform_L[824][7] = l_cell_wire[880];							inform_L[952][7] = l_cell_wire[881];							inform_L[825][7] = l_cell_wire[882];							inform_L[953][7] = l_cell_wire[883];							inform_L[826][7] = l_cell_wire[884];							inform_L[954][7] = l_cell_wire[885];							inform_L[827][7] = l_cell_wire[886];							inform_L[955][7] = l_cell_wire[887];							inform_L[828][7] = l_cell_wire[888];							inform_L[956][7] = l_cell_wire[889];							inform_L[829][7] = l_cell_wire[890];							inform_L[957][7] = l_cell_wire[891];							inform_L[830][7] = l_cell_wire[892];							inform_L[958][7] = l_cell_wire[893];							inform_L[831][7] = l_cell_wire[894];							inform_L[959][7] = l_cell_wire[895];							inform_L[832][7] = l_cell_wire[896];							inform_L[960][7] = l_cell_wire[897];							inform_L[833][7] = l_cell_wire[898];							inform_L[961][7] = l_cell_wire[899];							inform_L[834][7] = l_cell_wire[900];							inform_L[962][7] = l_cell_wire[901];							inform_L[835][7] = l_cell_wire[902];							inform_L[963][7] = l_cell_wire[903];							inform_L[836][7] = l_cell_wire[904];							inform_L[964][7] = l_cell_wire[905];							inform_L[837][7] = l_cell_wire[906];							inform_L[965][7] = l_cell_wire[907];							inform_L[838][7] = l_cell_wire[908];							inform_L[966][7] = l_cell_wire[909];							inform_L[839][7] = l_cell_wire[910];							inform_L[967][7] = l_cell_wire[911];							inform_L[840][7] = l_cell_wire[912];							inform_L[968][7] = l_cell_wire[913];							inform_L[841][7] = l_cell_wire[914];							inform_L[969][7] = l_cell_wire[915];							inform_L[842][7] = l_cell_wire[916];							inform_L[970][7] = l_cell_wire[917];							inform_L[843][7] = l_cell_wire[918];							inform_L[971][7] = l_cell_wire[919];							inform_L[844][7] = l_cell_wire[920];							inform_L[972][7] = l_cell_wire[921];							inform_L[845][7] = l_cell_wire[922];							inform_L[973][7] = l_cell_wire[923];							inform_L[846][7] = l_cell_wire[924];							inform_L[974][7] = l_cell_wire[925];							inform_L[847][7] = l_cell_wire[926];							inform_L[975][7] = l_cell_wire[927];							inform_L[848][7] = l_cell_wire[928];							inform_L[976][7] = l_cell_wire[929];							inform_L[849][7] = l_cell_wire[930];							inform_L[977][7] = l_cell_wire[931];							inform_L[850][7] = l_cell_wire[932];							inform_L[978][7] = l_cell_wire[933];							inform_L[851][7] = l_cell_wire[934];							inform_L[979][7] = l_cell_wire[935];							inform_L[852][7] = l_cell_wire[936];							inform_L[980][7] = l_cell_wire[937];							inform_L[853][7] = l_cell_wire[938];							inform_L[981][7] = l_cell_wire[939];							inform_L[854][7] = l_cell_wire[940];							inform_L[982][7] = l_cell_wire[941];							inform_L[855][7] = l_cell_wire[942];							inform_L[983][7] = l_cell_wire[943];							inform_L[856][7] = l_cell_wire[944];							inform_L[984][7] = l_cell_wire[945];							inform_L[857][7] = l_cell_wire[946];							inform_L[985][7] = l_cell_wire[947];							inform_L[858][7] = l_cell_wire[948];							inform_L[986][7] = l_cell_wire[949];							inform_L[859][7] = l_cell_wire[950];							inform_L[987][7] = l_cell_wire[951];							inform_L[860][7] = l_cell_wire[952];							inform_L[988][7] = l_cell_wire[953];							inform_L[861][7] = l_cell_wire[954];							inform_L[989][7] = l_cell_wire[955];							inform_L[862][7] = l_cell_wire[956];							inform_L[990][7] = l_cell_wire[957];							inform_L[863][7] = l_cell_wire[958];							inform_L[991][7] = l_cell_wire[959];							inform_L[864][7] = l_cell_wire[960];							inform_L[992][7] = l_cell_wire[961];							inform_L[865][7] = l_cell_wire[962];							inform_L[993][7] = l_cell_wire[963];							inform_L[866][7] = l_cell_wire[964];							inform_L[994][7] = l_cell_wire[965];							inform_L[867][7] = l_cell_wire[966];							inform_L[995][7] = l_cell_wire[967];							inform_L[868][7] = l_cell_wire[968];							inform_L[996][7] = l_cell_wire[969];							inform_L[869][7] = l_cell_wire[970];							inform_L[997][7] = l_cell_wire[971];							inform_L[870][7] = l_cell_wire[972];							inform_L[998][7] = l_cell_wire[973];							inform_L[871][7] = l_cell_wire[974];							inform_L[999][7] = l_cell_wire[975];							inform_L[872][7] = l_cell_wire[976];							inform_L[1000][7] = l_cell_wire[977];							inform_L[873][7] = l_cell_wire[978];							inform_L[1001][7] = l_cell_wire[979];							inform_L[874][7] = l_cell_wire[980];							inform_L[1002][7] = l_cell_wire[981];							inform_L[875][7] = l_cell_wire[982];							inform_L[1003][7] = l_cell_wire[983];							inform_L[876][7] = l_cell_wire[984];							inform_L[1004][7] = l_cell_wire[985];							inform_L[877][7] = l_cell_wire[986];							inform_L[1005][7] = l_cell_wire[987];							inform_L[878][7] = l_cell_wire[988];							inform_L[1006][7] = l_cell_wire[989];							inform_L[879][7] = l_cell_wire[990];							inform_L[1007][7] = l_cell_wire[991];							inform_L[880][7] = l_cell_wire[992];							inform_L[1008][7] = l_cell_wire[993];							inform_L[881][7] = l_cell_wire[994];							inform_L[1009][7] = l_cell_wire[995];							inform_L[882][7] = l_cell_wire[996];							inform_L[1010][7] = l_cell_wire[997];							inform_L[883][7] = l_cell_wire[998];							inform_L[1011][7] = l_cell_wire[999];							inform_L[884][7] = l_cell_wire[1000];							inform_L[1012][7] = l_cell_wire[1001];							inform_L[885][7] = l_cell_wire[1002];							inform_L[1013][7] = l_cell_wire[1003];							inform_L[886][7] = l_cell_wire[1004];							inform_L[1014][7] = l_cell_wire[1005];							inform_L[887][7] = l_cell_wire[1006];							inform_L[1015][7] = l_cell_wire[1007];							inform_L[888][7] = l_cell_wire[1008];							inform_L[1016][7] = l_cell_wire[1009];							inform_L[889][7] = l_cell_wire[1010];							inform_L[1017][7] = l_cell_wire[1011];							inform_L[890][7] = l_cell_wire[1012];							inform_L[1018][7] = l_cell_wire[1013];							inform_L[891][7] = l_cell_wire[1014];							inform_L[1019][7] = l_cell_wire[1015];							inform_L[892][7] = l_cell_wire[1016];							inform_L[1020][7] = l_cell_wire[1017];							inform_L[893][7] = l_cell_wire[1018];							inform_L[1021][7] = l_cell_wire[1019];							inform_L[894][7] = l_cell_wire[1020];							inform_L[1022][7] = l_cell_wire[1021];							inform_L[895][7] = l_cell_wire[1022];							inform_L[1023][7] = l_cell_wire[1023];						end
						9:						begin							inform_R[0][9] = r_cell_wire[0];							inform_R[256][9] = r_cell_wire[1];							inform_R[1][9] = r_cell_wire[2];							inform_R[257][9] = r_cell_wire[3];							inform_R[2][9] = r_cell_wire[4];							inform_R[258][9] = r_cell_wire[5];							inform_R[3][9] = r_cell_wire[6];							inform_R[259][9] = r_cell_wire[7];							inform_R[4][9] = r_cell_wire[8];							inform_R[260][9] = r_cell_wire[9];							inform_R[5][9] = r_cell_wire[10];							inform_R[261][9] = r_cell_wire[11];							inform_R[6][9] = r_cell_wire[12];							inform_R[262][9] = r_cell_wire[13];							inform_R[7][9] = r_cell_wire[14];							inform_R[263][9] = r_cell_wire[15];							inform_R[8][9] = r_cell_wire[16];							inform_R[264][9] = r_cell_wire[17];							inform_R[9][9] = r_cell_wire[18];							inform_R[265][9] = r_cell_wire[19];							inform_R[10][9] = r_cell_wire[20];							inform_R[266][9] = r_cell_wire[21];							inform_R[11][9] = r_cell_wire[22];							inform_R[267][9] = r_cell_wire[23];							inform_R[12][9] = r_cell_wire[24];							inform_R[268][9] = r_cell_wire[25];							inform_R[13][9] = r_cell_wire[26];							inform_R[269][9] = r_cell_wire[27];							inform_R[14][9] = r_cell_wire[28];							inform_R[270][9] = r_cell_wire[29];							inform_R[15][9] = r_cell_wire[30];							inform_R[271][9] = r_cell_wire[31];							inform_R[16][9] = r_cell_wire[32];							inform_R[272][9] = r_cell_wire[33];							inform_R[17][9] = r_cell_wire[34];							inform_R[273][9] = r_cell_wire[35];							inform_R[18][9] = r_cell_wire[36];							inform_R[274][9] = r_cell_wire[37];							inform_R[19][9] = r_cell_wire[38];							inform_R[275][9] = r_cell_wire[39];							inform_R[20][9] = r_cell_wire[40];							inform_R[276][9] = r_cell_wire[41];							inform_R[21][9] = r_cell_wire[42];							inform_R[277][9] = r_cell_wire[43];							inform_R[22][9] = r_cell_wire[44];							inform_R[278][9] = r_cell_wire[45];							inform_R[23][9] = r_cell_wire[46];							inform_R[279][9] = r_cell_wire[47];							inform_R[24][9] = r_cell_wire[48];							inform_R[280][9] = r_cell_wire[49];							inform_R[25][9] = r_cell_wire[50];							inform_R[281][9] = r_cell_wire[51];							inform_R[26][9] = r_cell_wire[52];							inform_R[282][9] = r_cell_wire[53];							inform_R[27][9] = r_cell_wire[54];							inform_R[283][9] = r_cell_wire[55];							inform_R[28][9] = r_cell_wire[56];							inform_R[284][9] = r_cell_wire[57];							inform_R[29][9] = r_cell_wire[58];							inform_R[285][9] = r_cell_wire[59];							inform_R[30][9] = r_cell_wire[60];							inform_R[286][9] = r_cell_wire[61];							inform_R[31][9] = r_cell_wire[62];							inform_R[287][9] = r_cell_wire[63];							inform_R[32][9] = r_cell_wire[64];							inform_R[288][9] = r_cell_wire[65];							inform_R[33][9] = r_cell_wire[66];							inform_R[289][9] = r_cell_wire[67];							inform_R[34][9] = r_cell_wire[68];							inform_R[290][9] = r_cell_wire[69];							inform_R[35][9] = r_cell_wire[70];							inform_R[291][9] = r_cell_wire[71];							inform_R[36][9] = r_cell_wire[72];							inform_R[292][9] = r_cell_wire[73];							inform_R[37][9] = r_cell_wire[74];							inform_R[293][9] = r_cell_wire[75];							inform_R[38][9] = r_cell_wire[76];							inform_R[294][9] = r_cell_wire[77];							inform_R[39][9] = r_cell_wire[78];							inform_R[295][9] = r_cell_wire[79];							inform_R[40][9] = r_cell_wire[80];							inform_R[296][9] = r_cell_wire[81];							inform_R[41][9] = r_cell_wire[82];							inform_R[297][9] = r_cell_wire[83];							inform_R[42][9] = r_cell_wire[84];							inform_R[298][9] = r_cell_wire[85];							inform_R[43][9] = r_cell_wire[86];							inform_R[299][9] = r_cell_wire[87];							inform_R[44][9] = r_cell_wire[88];							inform_R[300][9] = r_cell_wire[89];							inform_R[45][9] = r_cell_wire[90];							inform_R[301][9] = r_cell_wire[91];							inform_R[46][9] = r_cell_wire[92];							inform_R[302][9] = r_cell_wire[93];							inform_R[47][9] = r_cell_wire[94];							inform_R[303][9] = r_cell_wire[95];							inform_R[48][9] = r_cell_wire[96];							inform_R[304][9] = r_cell_wire[97];							inform_R[49][9] = r_cell_wire[98];							inform_R[305][9] = r_cell_wire[99];							inform_R[50][9] = r_cell_wire[100];							inform_R[306][9] = r_cell_wire[101];							inform_R[51][9] = r_cell_wire[102];							inform_R[307][9] = r_cell_wire[103];							inform_R[52][9] = r_cell_wire[104];							inform_R[308][9] = r_cell_wire[105];							inform_R[53][9] = r_cell_wire[106];							inform_R[309][9] = r_cell_wire[107];							inform_R[54][9] = r_cell_wire[108];							inform_R[310][9] = r_cell_wire[109];							inform_R[55][9] = r_cell_wire[110];							inform_R[311][9] = r_cell_wire[111];							inform_R[56][9] = r_cell_wire[112];							inform_R[312][9] = r_cell_wire[113];							inform_R[57][9] = r_cell_wire[114];							inform_R[313][9] = r_cell_wire[115];							inform_R[58][9] = r_cell_wire[116];							inform_R[314][9] = r_cell_wire[117];							inform_R[59][9] = r_cell_wire[118];							inform_R[315][9] = r_cell_wire[119];							inform_R[60][9] = r_cell_wire[120];							inform_R[316][9] = r_cell_wire[121];							inform_R[61][9] = r_cell_wire[122];							inform_R[317][9] = r_cell_wire[123];							inform_R[62][9] = r_cell_wire[124];							inform_R[318][9] = r_cell_wire[125];							inform_R[63][9] = r_cell_wire[126];							inform_R[319][9] = r_cell_wire[127];							inform_R[64][9] = r_cell_wire[128];							inform_R[320][9] = r_cell_wire[129];							inform_R[65][9] = r_cell_wire[130];							inform_R[321][9] = r_cell_wire[131];							inform_R[66][9] = r_cell_wire[132];							inform_R[322][9] = r_cell_wire[133];							inform_R[67][9] = r_cell_wire[134];							inform_R[323][9] = r_cell_wire[135];							inform_R[68][9] = r_cell_wire[136];							inform_R[324][9] = r_cell_wire[137];							inform_R[69][9] = r_cell_wire[138];							inform_R[325][9] = r_cell_wire[139];							inform_R[70][9] = r_cell_wire[140];							inform_R[326][9] = r_cell_wire[141];							inform_R[71][9] = r_cell_wire[142];							inform_R[327][9] = r_cell_wire[143];							inform_R[72][9] = r_cell_wire[144];							inform_R[328][9] = r_cell_wire[145];							inform_R[73][9] = r_cell_wire[146];							inform_R[329][9] = r_cell_wire[147];							inform_R[74][9] = r_cell_wire[148];							inform_R[330][9] = r_cell_wire[149];							inform_R[75][9] = r_cell_wire[150];							inform_R[331][9] = r_cell_wire[151];							inform_R[76][9] = r_cell_wire[152];							inform_R[332][9] = r_cell_wire[153];							inform_R[77][9] = r_cell_wire[154];							inform_R[333][9] = r_cell_wire[155];							inform_R[78][9] = r_cell_wire[156];							inform_R[334][9] = r_cell_wire[157];							inform_R[79][9] = r_cell_wire[158];							inform_R[335][9] = r_cell_wire[159];							inform_R[80][9] = r_cell_wire[160];							inform_R[336][9] = r_cell_wire[161];							inform_R[81][9] = r_cell_wire[162];							inform_R[337][9] = r_cell_wire[163];							inform_R[82][9] = r_cell_wire[164];							inform_R[338][9] = r_cell_wire[165];							inform_R[83][9] = r_cell_wire[166];							inform_R[339][9] = r_cell_wire[167];							inform_R[84][9] = r_cell_wire[168];							inform_R[340][9] = r_cell_wire[169];							inform_R[85][9] = r_cell_wire[170];							inform_R[341][9] = r_cell_wire[171];							inform_R[86][9] = r_cell_wire[172];							inform_R[342][9] = r_cell_wire[173];							inform_R[87][9] = r_cell_wire[174];							inform_R[343][9] = r_cell_wire[175];							inform_R[88][9] = r_cell_wire[176];							inform_R[344][9] = r_cell_wire[177];							inform_R[89][9] = r_cell_wire[178];							inform_R[345][9] = r_cell_wire[179];							inform_R[90][9] = r_cell_wire[180];							inform_R[346][9] = r_cell_wire[181];							inform_R[91][9] = r_cell_wire[182];							inform_R[347][9] = r_cell_wire[183];							inform_R[92][9] = r_cell_wire[184];							inform_R[348][9] = r_cell_wire[185];							inform_R[93][9] = r_cell_wire[186];							inform_R[349][9] = r_cell_wire[187];							inform_R[94][9] = r_cell_wire[188];							inform_R[350][9] = r_cell_wire[189];							inform_R[95][9] = r_cell_wire[190];							inform_R[351][9] = r_cell_wire[191];							inform_R[96][9] = r_cell_wire[192];							inform_R[352][9] = r_cell_wire[193];							inform_R[97][9] = r_cell_wire[194];							inform_R[353][9] = r_cell_wire[195];							inform_R[98][9] = r_cell_wire[196];							inform_R[354][9] = r_cell_wire[197];							inform_R[99][9] = r_cell_wire[198];							inform_R[355][9] = r_cell_wire[199];							inform_R[100][9] = r_cell_wire[200];							inform_R[356][9] = r_cell_wire[201];							inform_R[101][9] = r_cell_wire[202];							inform_R[357][9] = r_cell_wire[203];							inform_R[102][9] = r_cell_wire[204];							inform_R[358][9] = r_cell_wire[205];							inform_R[103][9] = r_cell_wire[206];							inform_R[359][9] = r_cell_wire[207];							inform_R[104][9] = r_cell_wire[208];							inform_R[360][9] = r_cell_wire[209];							inform_R[105][9] = r_cell_wire[210];							inform_R[361][9] = r_cell_wire[211];							inform_R[106][9] = r_cell_wire[212];							inform_R[362][9] = r_cell_wire[213];							inform_R[107][9] = r_cell_wire[214];							inform_R[363][9] = r_cell_wire[215];							inform_R[108][9] = r_cell_wire[216];							inform_R[364][9] = r_cell_wire[217];							inform_R[109][9] = r_cell_wire[218];							inform_R[365][9] = r_cell_wire[219];							inform_R[110][9] = r_cell_wire[220];							inform_R[366][9] = r_cell_wire[221];							inform_R[111][9] = r_cell_wire[222];							inform_R[367][9] = r_cell_wire[223];							inform_R[112][9] = r_cell_wire[224];							inform_R[368][9] = r_cell_wire[225];							inform_R[113][9] = r_cell_wire[226];							inform_R[369][9] = r_cell_wire[227];							inform_R[114][9] = r_cell_wire[228];							inform_R[370][9] = r_cell_wire[229];							inform_R[115][9] = r_cell_wire[230];							inform_R[371][9] = r_cell_wire[231];							inform_R[116][9] = r_cell_wire[232];							inform_R[372][9] = r_cell_wire[233];							inform_R[117][9] = r_cell_wire[234];							inform_R[373][9] = r_cell_wire[235];							inform_R[118][9] = r_cell_wire[236];							inform_R[374][9] = r_cell_wire[237];							inform_R[119][9] = r_cell_wire[238];							inform_R[375][9] = r_cell_wire[239];							inform_R[120][9] = r_cell_wire[240];							inform_R[376][9] = r_cell_wire[241];							inform_R[121][9] = r_cell_wire[242];							inform_R[377][9] = r_cell_wire[243];							inform_R[122][9] = r_cell_wire[244];							inform_R[378][9] = r_cell_wire[245];							inform_R[123][9] = r_cell_wire[246];							inform_R[379][9] = r_cell_wire[247];							inform_R[124][9] = r_cell_wire[248];							inform_R[380][9] = r_cell_wire[249];							inform_R[125][9] = r_cell_wire[250];							inform_R[381][9] = r_cell_wire[251];							inform_R[126][9] = r_cell_wire[252];							inform_R[382][9] = r_cell_wire[253];							inform_R[127][9] = r_cell_wire[254];							inform_R[383][9] = r_cell_wire[255];							inform_R[128][9] = r_cell_wire[256];							inform_R[384][9] = r_cell_wire[257];							inform_R[129][9] = r_cell_wire[258];							inform_R[385][9] = r_cell_wire[259];							inform_R[130][9] = r_cell_wire[260];							inform_R[386][9] = r_cell_wire[261];							inform_R[131][9] = r_cell_wire[262];							inform_R[387][9] = r_cell_wire[263];							inform_R[132][9] = r_cell_wire[264];							inform_R[388][9] = r_cell_wire[265];							inform_R[133][9] = r_cell_wire[266];							inform_R[389][9] = r_cell_wire[267];							inform_R[134][9] = r_cell_wire[268];							inform_R[390][9] = r_cell_wire[269];							inform_R[135][9] = r_cell_wire[270];							inform_R[391][9] = r_cell_wire[271];							inform_R[136][9] = r_cell_wire[272];							inform_R[392][9] = r_cell_wire[273];							inform_R[137][9] = r_cell_wire[274];							inform_R[393][9] = r_cell_wire[275];							inform_R[138][9] = r_cell_wire[276];							inform_R[394][9] = r_cell_wire[277];							inform_R[139][9] = r_cell_wire[278];							inform_R[395][9] = r_cell_wire[279];							inform_R[140][9] = r_cell_wire[280];							inform_R[396][9] = r_cell_wire[281];							inform_R[141][9] = r_cell_wire[282];							inform_R[397][9] = r_cell_wire[283];							inform_R[142][9] = r_cell_wire[284];							inform_R[398][9] = r_cell_wire[285];							inform_R[143][9] = r_cell_wire[286];							inform_R[399][9] = r_cell_wire[287];							inform_R[144][9] = r_cell_wire[288];							inform_R[400][9] = r_cell_wire[289];							inform_R[145][9] = r_cell_wire[290];							inform_R[401][9] = r_cell_wire[291];							inform_R[146][9] = r_cell_wire[292];							inform_R[402][9] = r_cell_wire[293];							inform_R[147][9] = r_cell_wire[294];							inform_R[403][9] = r_cell_wire[295];							inform_R[148][9] = r_cell_wire[296];							inform_R[404][9] = r_cell_wire[297];							inform_R[149][9] = r_cell_wire[298];							inform_R[405][9] = r_cell_wire[299];							inform_R[150][9] = r_cell_wire[300];							inform_R[406][9] = r_cell_wire[301];							inform_R[151][9] = r_cell_wire[302];							inform_R[407][9] = r_cell_wire[303];							inform_R[152][9] = r_cell_wire[304];							inform_R[408][9] = r_cell_wire[305];							inform_R[153][9] = r_cell_wire[306];							inform_R[409][9] = r_cell_wire[307];							inform_R[154][9] = r_cell_wire[308];							inform_R[410][9] = r_cell_wire[309];							inform_R[155][9] = r_cell_wire[310];							inform_R[411][9] = r_cell_wire[311];							inform_R[156][9] = r_cell_wire[312];							inform_R[412][9] = r_cell_wire[313];							inform_R[157][9] = r_cell_wire[314];							inform_R[413][9] = r_cell_wire[315];							inform_R[158][9] = r_cell_wire[316];							inform_R[414][9] = r_cell_wire[317];							inform_R[159][9] = r_cell_wire[318];							inform_R[415][9] = r_cell_wire[319];							inform_R[160][9] = r_cell_wire[320];							inform_R[416][9] = r_cell_wire[321];							inform_R[161][9] = r_cell_wire[322];							inform_R[417][9] = r_cell_wire[323];							inform_R[162][9] = r_cell_wire[324];							inform_R[418][9] = r_cell_wire[325];							inform_R[163][9] = r_cell_wire[326];							inform_R[419][9] = r_cell_wire[327];							inform_R[164][9] = r_cell_wire[328];							inform_R[420][9] = r_cell_wire[329];							inform_R[165][9] = r_cell_wire[330];							inform_R[421][9] = r_cell_wire[331];							inform_R[166][9] = r_cell_wire[332];							inform_R[422][9] = r_cell_wire[333];							inform_R[167][9] = r_cell_wire[334];							inform_R[423][9] = r_cell_wire[335];							inform_R[168][9] = r_cell_wire[336];							inform_R[424][9] = r_cell_wire[337];							inform_R[169][9] = r_cell_wire[338];							inform_R[425][9] = r_cell_wire[339];							inform_R[170][9] = r_cell_wire[340];							inform_R[426][9] = r_cell_wire[341];							inform_R[171][9] = r_cell_wire[342];							inform_R[427][9] = r_cell_wire[343];							inform_R[172][9] = r_cell_wire[344];							inform_R[428][9] = r_cell_wire[345];							inform_R[173][9] = r_cell_wire[346];							inform_R[429][9] = r_cell_wire[347];							inform_R[174][9] = r_cell_wire[348];							inform_R[430][9] = r_cell_wire[349];							inform_R[175][9] = r_cell_wire[350];							inform_R[431][9] = r_cell_wire[351];							inform_R[176][9] = r_cell_wire[352];							inform_R[432][9] = r_cell_wire[353];							inform_R[177][9] = r_cell_wire[354];							inform_R[433][9] = r_cell_wire[355];							inform_R[178][9] = r_cell_wire[356];							inform_R[434][9] = r_cell_wire[357];							inform_R[179][9] = r_cell_wire[358];							inform_R[435][9] = r_cell_wire[359];							inform_R[180][9] = r_cell_wire[360];							inform_R[436][9] = r_cell_wire[361];							inform_R[181][9] = r_cell_wire[362];							inform_R[437][9] = r_cell_wire[363];							inform_R[182][9] = r_cell_wire[364];							inform_R[438][9] = r_cell_wire[365];							inform_R[183][9] = r_cell_wire[366];							inform_R[439][9] = r_cell_wire[367];							inform_R[184][9] = r_cell_wire[368];							inform_R[440][9] = r_cell_wire[369];							inform_R[185][9] = r_cell_wire[370];							inform_R[441][9] = r_cell_wire[371];							inform_R[186][9] = r_cell_wire[372];							inform_R[442][9] = r_cell_wire[373];							inform_R[187][9] = r_cell_wire[374];							inform_R[443][9] = r_cell_wire[375];							inform_R[188][9] = r_cell_wire[376];							inform_R[444][9] = r_cell_wire[377];							inform_R[189][9] = r_cell_wire[378];							inform_R[445][9] = r_cell_wire[379];							inform_R[190][9] = r_cell_wire[380];							inform_R[446][9] = r_cell_wire[381];							inform_R[191][9] = r_cell_wire[382];							inform_R[447][9] = r_cell_wire[383];							inform_R[192][9] = r_cell_wire[384];							inform_R[448][9] = r_cell_wire[385];							inform_R[193][9] = r_cell_wire[386];							inform_R[449][9] = r_cell_wire[387];							inform_R[194][9] = r_cell_wire[388];							inform_R[450][9] = r_cell_wire[389];							inform_R[195][9] = r_cell_wire[390];							inform_R[451][9] = r_cell_wire[391];							inform_R[196][9] = r_cell_wire[392];							inform_R[452][9] = r_cell_wire[393];							inform_R[197][9] = r_cell_wire[394];							inform_R[453][9] = r_cell_wire[395];							inform_R[198][9] = r_cell_wire[396];							inform_R[454][9] = r_cell_wire[397];							inform_R[199][9] = r_cell_wire[398];							inform_R[455][9] = r_cell_wire[399];							inform_R[200][9] = r_cell_wire[400];							inform_R[456][9] = r_cell_wire[401];							inform_R[201][9] = r_cell_wire[402];							inform_R[457][9] = r_cell_wire[403];							inform_R[202][9] = r_cell_wire[404];							inform_R[458][9] = r_cell_wire[405];							inform_R[203][9] = r_cell_wire[406];							inform_R[459][9] = r_cell_wire[407];							inform_R[204][9] = r_cell_wire[408];							inform_R[460][9] = r_cell_wire[409];							inform_R[205][9] = r_cell_wire[410];							inform_R[461][9] = r_cell_wire[411];							inform_R[206][9] = r_cell_wire[412];							inform_R[462][9] = r_cell_wire[413];							inform_R[207][9] = r_cell_wire[414];							inform_R[463][9] = r_cell_wire[415];							inform_R[208][9] = r_cell_wire[416];							inform_R[464][9] = r_cell_wire[417];							inform_R[209][9] = r_cell_wire[418];							inform_R[465][9] = r_cell_wire[419];							inform_R[210][9] = r_cell_wire[420];							inform_R[466][9] = r_cell_wire[421];							inform_R[211][9] = r_cell_wire[422];							inform_R[467][9] = r_cell_wire[423];							inform_R[212][9] = r_cell_wire[424];							inform_R[468][9] = r_cell_wire[425];							inform_R[213][9] = r_cell_wire[426];							inform_R[469][9] = r_cell_wire[427];							inform_R[214][9] = r_cell_wire[428];							inform_R[470][9] = r_cell_wire[429];							inform_R[215][9] = r_cell_wire[430];							inform_R[471][9] = r_cell_wire[431];							inform_R[216][9] = r_cell_wire[432];							inform_R[472][9] = r_cell_wire[433];							inform_R[217][9] = r_cell_wire[434];							inform_R[473][9] = r_cell_wire[435];							inform_R[218][9] = r_cell_wire[436];							inform_R[474][9] = r_cell_wire[437];							inform_R[219][9] = r_cell_wire[438];							inform_R[475][9] = r_cell_wire[439];							inform_R[220][9] = r_cell_wire[440];							inform_R[476][9] = r_cell_wire[441];							inform_R[221][9] = r_cell_wire[442];							inform_R[477][9] = r_cell_wire[443];							inform_R[222][9] = r_cell_wire[444];							inform_R[478][9] = r_cell_wire[445];							inform_R[223][9] = r_cell_wire[446];							inform_R[479][9] = r_cell_wire[447];							inform_R[224][9] = r_cell_wire[448];							inform_R[480][9] = r_cell_wire[449];							inform_R[225][9] = r_cell_wire[450];							inform_R[481][9] = r_cell_wire[451];							inform_R[226][9] = r_cell_wire[452];							inform_R[482][9] = r_cell_wire[453];							inform_R[227][9] = r_cell_wire[454];							inform_R[483][9] = r_cell_wire[455];							inform_R[228][9] = r_cell_wire[456];							inform_R[484][9] = r_cell_wire[457];							inform_R[229][9] = r_cell_wire[458];							inform_R[485][9] = r_cell_wire[459];							inform_R[230][9] = r_cell_wire[460];							inform_R[486][9] = r_cell_wire[461];							inform_R[231][9] = r_cell_wire[462];							inform_R[487][9] = r_cell_wire[463];							inform_R[232][9] = r_cell_wire[464];							inform_R[488][9] = r_cell_wire[465];							inform_R[233][9] = r_cell_wire[466];							inform_R[489][9] = r_cell_wire[467];							inform_R[234][9] = r_cell_wire[468];							inform_R[490][9] = r_cell_wire[469];							inform_R[235][9] = r_cell_wire[470];							inform_R[491][9] = r_cell_wire[471];							inform_R[236][9] = r_cell_wire[472];							inform_R[492][9] = r_cell_wire[473];							inform_R[237][9] = r_cell_wire[474];							inform_R[493][9] = r_cell_wire[475];							inform_R[238][9] = r_cell_wire[476];							inform_R[494][9] = r_cell_wire[477];							inform_R[239][9] = r_cell_wire[478];							inform_R[495][9] = r_cell_wire[479];							inform_R[240][9] = r_cell_wire[480];							inform_R[496][9] = r_cell_wire[481];							inform_R[241][9] = r_cell_wire[482];							inform_R[497][9] = r_cell_wire[483];							inform_R[242][9] = r_cell_wire[484];							inform_R[498][9] = r_cell_wire[485];							inform_R[243][9] = r_cell_wire[486];							inform_R[499][9] = r_cell_wire[487];							inform_R[244][9] = r_cell_wire[488];							inform_R[500][9] = r_cell_wire[489];							inform_R[245][9] = r_cell_wire[490];							inform_R[501][9] = r_cell_wire[491];							inform_R[246][9] = r_cell_wire[492];							inform_R[502][9] = r_cell_wire[493];							inform_R[247][9] = r_cell_wire[494];							inform_R[503][9] = r_cell_wire[495];							inform_R[248][9] = r_cell_wire[496];							inform_R[504][9] = r_cell_wire[497];							inform_R[249][9] = r_cell_wire[498];							inform_R[505][9] = r_cell_wire[499];							inform_R[250][9] = r_cell_wire[500];							inform_R[506][9] = r_cell_wire[501];							inform_R[251][9] = r_cell_wire[502];							inform_R[507][9] = r_cell_wire[503];							inform_R[252][9] = r_cell_wire[504];							inform_R[508][9] = r_cell_wire[505];							inform_R[253][9] = r_cell_wire[506];							inform_R[509][9] = r_cell_wire[507];							inform_R[254][9] = r_cell_wire[508];							inform_R[510][9] = r_cell_wire[509];							inform_R[255][9] = r_cell_wire[510];							inform_R[511][9] = r_cell_wire[511];							inform_R[512][9] = r_cell_wire[512];							inform_R[768][9] = r_cell_wire[513];							inform_R[513][9] = r_cell_wire[514];							inform_R[769][9] = r_cell_wire[515];							inform_R[514][9] = r_cell_wire[516];							inform_R[770][9] = r_cell_wire[517];							inform_R[515][9] = r_cell_wire[518];							inform_R[771][9] = r_cell_wire[519];							inform_R[516][9] = r_cell_wire[520];							inform_R[772][9] = r_cell_wire[521];							inform_R[517][9] = r_cell_wire[522];							inform_R[773][9] = r_cell_wire[523];							inform_R[518][9] = r_cell_wire[524];							inform_R[774][9] = r_cell_wire[525];							inform_R[519][9] = r_cell_wire[526];							inform_R[775][9] = r_cell_wire[527];							inform_R[520][9] = r_cell_wire[528];							inform_R[776][9] = r_cell_wire[529];							inform_R[521][9] = r_cell_wire[530];							inform_R[777][9] = r_cell_wire[531];							inform_R[522][9] = r_cell_wire[532];							inform_R[778][9] = r_cell_wire[533];							inform_R[523][9] = r_cell_wire[534];							inform_R[779][9] = r_cell_wire[535];							inform_R[524][9] = r_cell_wire[536];							inform_R[780][9] = r_cell_wire[537];							inform_R[525][9] = r_cell_wire[538];							inform_R[781][9] = r_cell_wire[539];							inform_R[526][9] = r_cell_wire[540];							inform_R[782][9] = r_cell_wire[541];							inform_R[527][9] = r_cell_wire[542];							inform_R[783][9] = r_cell_wire[543];							inform_R[528][9] = r_cell_wire[544];							inform_R[784][9] = r_cell_wire[545];							inform_R[529][9] = r_cell_wire[546];							inform_R[785][9] = r_cell_wire[547];							inform_R[530][9] = r_cell_wire[548];							inform_R[786][9] = r_cell_wire[549];							inform_R[531][9] = r_cell_wire[550];							inform_R[787][9] = r_cell_wire[551];							inform_R[532][9] = r_cell_wire[552];							inform_R[788][9] = r_cell_wire[553];							inform_R[533][9] = r_cell_wire[554];							inform_R[789][9] = r_cell_wire[555];							inform_R[534][9] = r_cell_wire[556];							inform_R[790][9] = r_cell_wire[557];							inform_R[535][9] = r_cell_wire[558];							inform_R[791][9] = r_cell_wire[559];							inform_R[536][9] = r_cell_wire[560];							inform_R[792][9] = r_cell_wire[561];							inform_R[537][9] = r_cell_wire[562];							inform_R[793][9] = r_cell_wire[563];							inform_R[538][9] = r_cell_wire[564];							inform_R[794][9] = r_cell_wire[565];							inform_R[539][9] = r_cell_wire[566];							inform_R[795][9] = r_cell_wire[567];							inform_R[540][9] = r_cell_wire[568];							inform_R[796][9] = r_cell_wire[569];							inform_R[541][9] = r_cell_wire[570];							inform_R[797][9] = r_cell_wire[571];							inform_R[542][9] = r_cell_wire[572];							inform_R[798][9] = r_cell_wire[573];							inform_R[543][9] = r_cell_wire[574];							inform_R[799][9] = r_cell_wire[575];							inform_R[544][9] = r_cell_wire[576];							inform_R[800][9] = r_cell_wire[577];							inform_R[545][9] = r_cell_wire[578];							inform_R[801][9] = r_cell_wire[579];							inform_R[546][9] = r_cell_wire[580];							inform_R[802][9] = r_cell_wire[581];							inform_R[547][9] = r_cell_wire[582];							inform_R[803][9] = r_cell_wire[583];							inform_R[548][9] = r_cell_wire[584];							inform_R[804][9] = r_cell_wire[585];							inform_R[549][9] = r_cell_wire[586];							inform_R[805][9] = r_cell_wire[587];							inform_R[550][9] = r_cell_wire[588];							inform_R[806][9] = r_cell_wire[589];							inform_R[551][9] = r_cell_wire[590];							inform_R[807][9] = r_cell_wire[591];							inform_R[552][9] = r_cell_wire[592];							inform_R[808][9] = r_cell_wire[593];							inform_R[553][9] = r_cell_wire[594];							inform_R[809][9] = r_cell_wire[595];							inform_R[554][9] = r_cell_wire[596];							inform_R[810][9] = r_cell_wire[597];							inform_R[555][9] = r_cell_wire[598];							inform_R[811][9] = r_cell_wire[599];							inform_R[556][9] = r_cell_wire[600];							inform_R[812][9] = r_cell_wire[601];							inform_R[557][9] = r_cell_wire[602];							inform_R[813][9] = r_cell_wire[603];							inform_R[558][9] = r_cell_wire[604];							inform_R[814][9] = r_cell_wire[605];							inform_R[559][9] = r_cell_wire[606];							inform_R[815][9] = r_cell_wire[607];							inform_R[560][9] = r_cell_wire[608];							inform_R[816][9] = r_cell_wire[609];							inform_R[561][9] = r_cell_wire[610];							inform_R[817][9] = r_cell_wire[611];							inform_R[562][9] = r_cell_wire[612];							inform_R[818][9] = r_cell_wire[613];							inform_R[563][9] = r_cell_wire[614];							inform_R[819][9] = r_cell_wire[615];							inform_R[564][9] = r_cell_wire[616];							inform_R[820][9] = r_cell_wire[617];							inform_R[565][9] = r_cell_wire[618];							inform_R[821][9] = r_cell_wire[619];							inform_R[566][9] = r_cell_wire[620];							inform_R[822][9] = r_cell_wire[621];							inform_R[567][9] = r_cell_wire[622];							inform_R[823][9] = r_cell_wire[623];							inform_R[568][9] = r_cell_wire[624];							inform_R[824][9] = r_cell_wire[625];							inform_R[569][9] = r_cell_wire[626];							inform_R[825][9] = r_cell_wire[627];							inform_R[570][9] = r_cell_wire[628];							inform_R[826][9] = r_cell_wire[629];							inform_R[571][9] = r_cell_wire[630];							inform_R[827][9] = r_cell_wire[631];							inform_R[572][9] = r_cell_wire[632];							inform_R[828][9] = r_cell_wire[633];							inform_R[573][9] = r_cell_wire[634];							inform_R[829][9] = r_cell_wire[635];							inform_R[574][9] = r_cell_wire[636];							inform_R[830][9] = r_cell_wire[637];							inform_R[575][9] = r_cell_wire[638];							inform_R[831][9] = r_cell_wire[639];							inform_R[576][9] = r_cell_wire[640];							inform_R[832][9] = r_cell_wire[641];							inform_R[577][9] = r_cell_wire[642];							inform_R[833][9] = r_cell_wire[643];							inform_R[578][9] = r_cell_wire[644];							inform_R[834][9] = r_cell_wire[645];							inform_R[579][9] = r_cell_wire[646];							inform_R[835][9] = r_cell_wire[647];							inform_R[580][9] = r_cell_wire[648];							inform_R[836][9] = r_cell_wire[649];							inform_R[581][9] = r_cell_wire[650];							inform_R[837][9] = r_cell_wire[651];							inform_R[582][9] = r_cell_wire[652];							inform_R[838][9] = r_cell_wire[653];							inform_R[583][9] = r_cell_wire[654];							inform_R[839][9] = r_cell_wire[655];							inform_R[584][9] = r_cell_wire[656];							inform_R[840][9] = r_cell_wire[657];							inform_R[585][9] = r_cell_wire[658];							inform_R[841][9] = r_cell_wire[659];							inform_R[586][9] = r_cell_wire[660];							inform_R[842][9] = r_cell_wire[661];							inform_R[587][9] = r_cell_wire[662];							inform_R[843][9] = r_cell_wire[663];							inform_R[588][9] = r_cell_wire[664];							inform_R[844][9] = r_cell_wire[665];							inform_R[589][9] = r_cell_wire[666];							inform_R[845][9] = r_cell_wire[667];							inform_R[590][9] = r_cell_wire[668];							inform_R[846][9] = r_cell_wire[669];							inform_R[591][9] = r_cell_wire[670];							inform_R[847][9] = r_cell_wire[671];							inform_R[592][9] = r_cell_wire[672];							inform_R[848][9] = r_cell_wire[673];							inform_R[593][9] = r_cell_wire[674];							inform_R[849][9] = r_cell_wire[675];							inform_R[594][9] = r_cell_wire[676];							inform_R[850][9] = r_cell_wire[677];							inform_R[595][9] = r_cell_wire[678];							inform_R[851][9] = r_cell_wire[679];							inform_R[596][9] = r_cell_wire[680];							inform_R[852][9] = r_cell_wire[681];							inform_R[597][9] = r_cell_wire[682];							inform_R[853][9] = r_cell_wire[683];							inform_R[598][9] = r_cell_wire[684];							inform_R[854][9] = r_cell_wire[685];							inform_R[599][9] = r_cell_wire[686];							inform_R[855][9] = r_cell_wire[687];							inform_R[600][9] = r_cell_wire[688];							inform_R[856][9] = r_cell_wire[689];							inform_R[601][9] = r_cell_wire[690];							inform_R[857][9] = r_cell_wire[691];							inform_R[602][9] = r_cell_wire[692];							inform_R[858][9] = r_cell_wire[693];							inform_R[603][9] = r_cell_wire[694];							inform_R[859][9] = r_cell_wire[695];							inform_R[604][9] = r_cell_wire[696];							inform_R[860][9] = r_cell_wire[697];							inform_R[605][9] = r_cell_wire[698];							inform_R[861][9] = r_cell_wire[699];							inform_R[606][9] = r_cell_wire[700];							inform_R[862][9] = r_cell_wire[701];							inform_R[607][9] = r_cell_wire[702];							inform_R[863][9] = r_cell_wire[703];							inform_R[608][9] = r_cell_wire[704];							inform_R[864][9] = r_cell_wire[705];							inform_R[609][9] = r_cell_wire[706];							inform_R[865][9] = r_cell_wire[707];							inform_R[610][9] = r_cell_wire[708];							inform_R[866][9] = r_cell_wire[709];							inform_R[611][9] = r_cell_wire[710];							inform_R[867][9] = r_cell_wire[711];							inform_R[612][9] = r_cell_wire[712];							inform_R[868][9] = r_cell_wire[713];							inform_R[613][9] = r_cell_wire[714];							inform_R[869][9] = r_cell_wire[715];							inform_R[614][9] = r_cell_wire[716];							inform_R[870][9] = r_cell_wire[717];							inform_R[615][9] = r_cell_wire[718];							inform_R[871][9] = r_cell_wire[719];							inform_R[616][9] = r_cell_wire[720];							inform_R[872][9] = r_cell_wire[721];							inform_R[617][9] = r_cell_wire[722];							inform_R[873][9] = r_cell_wire[723];							inform_R[618][9] = r_cell_wire[724];							inform_R[874][9] = r_cell_wire[725];							inform_R[619][9] = r_cell_wire[726];							inform_R[875][9] = r_cell_wire[727];							inform_R[620][9] = r_cell_wire[728];							inform_R[876][9] = r_cell_wire[729];							inform_R[621][9] = r_cell_wire[730];							inform_R[877][9] = r_cell_wire[731];							inform_R[622][9] = r_cell_wire[732];							inform_R[878][9] = r_cell_wire[733];							inform_R[623][9] = r_cell_wire[734];							inform_R[879][9] = r_cell_wire[735];							inform_R[624][9] = r_cell_wire[736];							inform_R[880][9] = r_cell_wire[737];							inform_R[625][9] = r_cell_wire[738];							inform_R[881][9] = r_cell_wire[739];							inform_R[626][9] = r_cell_wire[740];							inform_R[882][9] = r_cell_wire[741];							inform_R[627][9] = r_cell_wire[742];							inform_R[883][9] = r_cell_wire[743];							inform_R[628][9] = r_cell_wire[744];							inform_R[884][9] = r_cell_wire[745];							inform_R[629][9] = r_cell_wire[746];							inform_R[885][9] = r_cell_wire[747];							inform_R[630][9] = r_cell_wire[748];							inform_R[886][9] = r_cell_wire[749];							inform_R[631][9] = r_cell_wire[750];							inform_R[887][9] = r_cell_wire[751];							inform_R[632][9] = r_cell_wire[752];							inform_R[888][9] = r_cell_wire[753];							inform_R[633][9] = r_cell_wire[754];							inform_R[889][9] = r_cell_wire[755];							inform_R[634][9] = r_cell_wire[756];							inform_R[890][9] = r_cell_wire[757];							inform_R[635][9] = r_cell_wire[758];							inform_R[891][9] = r_cell_wire[759];							inform_R[636][9] = r_cell_wire[760];							inform_R[892][9] = r_cell_wire[761];							inform_R[637][9] = r_cell_wire[762];							inform_R[893][9] = r_cell_wire[763];							inform_R[638][9] = r_cell_wire[764];							inform_R[894][9] = r_cell_wire[765];							inform_R[639][9] = r_cell_wire[766];							inform_R[895][9] = r_cell_wire[767];							inform_R[640][9] = r_cell_wire[768];							inform_R[896][9] = r_cell_wire[769];							inform_R[641][9] = r_cell_wire[770];							inform_R[897][9] = r_cell_wire[771];							inform_R[642][9] = r_cell_wire[772];							inform_R[898][9] = r_cell_wire[773];							inform_R[643][9] = r_cell_wire[774];							inform_R[899][9] = r_cell_wire[775];							inform_R[644][9] = r_cell_wire[776];							inform_R[900][9] = r_cell_wire[777];							inform_R[645][9] = r_cell_wire[778];							inform_R[901][9] = r_cell_wire[779];							inform_R[646][9] = r_cell_wire[780];							inform_R[902][9] = r_cell_wire[781];							inform_R[647][9] = r_cell_wire[782];							inform_R[903][9] = r_cell_wire[783];							inform_R[648][9] = r_cell_wire[784];							inform_R[904][9] = r_cell_wire[785];							inform_R[649][9] = r_cell_wire[786];							inform_R[905][9] = r_cell_wire[787];							inform_R[650][9] = r_cell_wire[788];							inform_R[906][9] = r_cell_wire[789];							inform_R[651][9] = r_cell_wire[790];							inform_R[907][9] = r_cell_wire[791];							inform_R[652][9] = r_cell_wire[792];							inform_R[908][9] = r_cell_wire[793];							inform_R[653][9] = r_cell_wire[794];							inform_R[909][9] = r_cell_wire[795];							inform_R[654][9] = r_cell_wire[796];							inform_R[910][9] = r_cell_wire[797];							inform_R[655][9] = r_cell_wire[798];							inform_R[911][9] = r_cell_wire[799];							inform_R[656][9] = r_cell_wire[800];							inform_R[912][9] = r_cell_wire[801];							inform_R[657][9] = r_cell_wire[802];							inform_R[913][9] = r_cell_wire[803];							inform_R[658][9] = r_cell_wire[804];							inform_R[914][9] = r_cell_wire[805];							inform_R[659][9] = r_cell_wire[806];							inform_R[915][9] = r_cell_wire[807];							inform_R[660][9] = r_cell_wire[808];							inform_R[916][9] = r_cell_wire[809];							inform_R[661][9] = r_cell_wire[810];							inform_R[917][9] = r_cell_wire[811];							inform_R[662][9] = r_cell_wire[812];							inform_R[918][9] = r_cell_wire[813];							inform_R[663][9] = r_cell_wire[814];							inform_R[919][9] = r_cell_wire[815];							inform_R[664][9] = r_cell_wire[816];							inform_R[920][9] = r_cell_wire[817];							inform_R[665][9] = r_cell_wire[818];							inform_R[921][9] = r_cell_wire[819];							inform_R[666][9] = r_cell_wire[820];							inform_R[922][9] = r_cell_wire[821];							inform_R[667][9] = r_cell_wire[822];							inform_R[923][9] = r_cell_wire[823];							inform_R[668][9] = r_cell_wire[824];							inform_R[924][9] = r_cell_wire[825];							inform_R[669][9] = r_cell_wire[826];							inform_R[925][9] = r_cell_wire[827];							inform_R[670][9] = r_cell_wire[828];							inform_R[926][9] = r_cell_wire[829];							inform_R[671][9] = r_cell_wire[830];							inform_R[927][9] = r_cell_wire[831];							inform_R[672][9] = r_cell_wire[832];							inform_R[928][9] = r_cell_wire[833];							inform_R[673][9] = r_cell_wire[834];							inform_R[929][9] = r_cell_wire[835];							inform_R[674][9] = r_cell_wire[836];							inform_R[930][9] = r_cell_wire[837];							inform_R[675][9] = r_cell_wire[838];							inform_R[931][9] = r_cell_wire[839];							inform_R[676][9] = r_cell_wire[840];							inform_R[932][9] = r_cell_wire[841];							inform_R[677][9] = r_cell_wire[842];							inform_R[933][9] = r_cell_wire[843];							inform_R[678][9] = r_cell_wire[844];							inform_R[934][9] = r_cell_wire[845];							inform_R[679][9] = r_cell_wire[846];							inform_R[935][9] = r_cell_wire[847];							inform_R[680][9] = r_cell_wire[848];							inform_R[936][9] = r_cell_wire[849];							inform_R[681][9] = r_cell_wire[850];							inform_R[937][9] = r_cell_wire[851];							inform_R[682][9] = r_cell_wire[852];							inform_R[938][9] = r_cell_wire[853];							inform_R[683][9] = r_cell_wire[854];							inform_R[939][9] = r_cell_wire[855];							inform_R[684][9] = r_cell_wire[856];							inform_R[940][9] = r_cell_wire[857];							inform_R[685][9] = r_cell_wire[858];							inform_R[941][9] = r_cell_wire[859];							inform_R[686][9] = r_cell_wire[860];							inform_R[942][9] = r_cell_wire[861];							inform_R[687][9] = r_cell_wire[862];							inform_R[943][9] = r_cell_wire[863];							inform_R[688][9] = r_cell_wire[864];							inform_R[944][9] = r_cell_wire[865];							inform_R[689][9] = r_cell_wire[866];							inform_R[945][9] = r_cell_wire[867];							inform_R[690][9] = r_cell_wire[868];							inform_R[946][9] = r_cell_wire[869];							inform_R[691][9] = r_cell_wire[870];							inform_R[947][9] = r_cell_wire[871];							inform_R[692][9] = r_cell_wire[872];							inform_R[948][9] = r_cell_wire[873];							inform_R[693][9] = r_cell_wire[874];							inform_R[949][9] = r_cell_wire[875];							inform_R[694][9] = r_cell_wire[876];							inform_R[950][9] = r_cell_wire[877];							inform_R[695][9] = r_cell_wire[878];							inform_R[951][9] = r_cell_wire[879];							inform_R[696][9] = r_cell_wire[880];							inform_R[952][9] = r_cell_wire[881];							inform_R[697][9] = r_cell_wire[882];							inform_R[953][9] = r_cell_wire[883];							inform_R[698][9] = r_cell_wire[884];							inform_R[954][9] = r_cell_wire[885];							inform_R[699][9] = r_cell_wire[886];							inform_R[955][9] = r_cell_wire[887];							inform_R[700][9] = r_cell_wire[888];							inform_R[956][9] = r_cell_wire[889];							inform_R[701][9] = r_cell_wire[890];							inform_R[957][9] = r_cell_wire[891];							inform_R[702][9] = r_cell_wire[892];							inform_R[958][9] = r_cell_wire[893];							inform_R[703][9] = r_cell_wire[894];							inform_R[959][9] = r_cell_wire[895];							inform_R[704][9] = r_cell_wire[896];							inform_R[960][9] = r_cell_wire[897];							inform_R[705][9] = r_cell_wire[898];							inform_R[961][9] = r_cell_wire[899];							inform_R[706][9] = r_cell_wire[900];							inform_R[962][9] = r_cell_wire[901];							inform_R[707][9] = r_cell_wire[902];							inform_R[963][9] = r_cell_wire[903];							inform_R[708][9] = r_cell_wire[904];							inform_R[964][9] = r_cell_wire[905];							inform_R[709][9] = r_cell_wire[906];							inform_R[965][9] = r_cell_wire[907];							inform_R[710][9] = r_cell_wire[908];							inform_R[966][9] = r_cell_wire[909];							inform_R[711][9] = r_cell_wire[910];							inform_R[967][9] = r_cell_wire[911];							inform_R[712][9] = r_cell_wire[912];							inform_R[968][9] = r_cell_wire[913];							inform_R[713][9] = r_cell_wire[914];							inform_R[969][9] = r_cell_wire[915];							inform_R[714][9] = r_cell_wire[916];							inform_R[970][9] = r_cell_wire[917];							inform_R[715][9] = r_cell_wire[918];							inform_R[971][9] = r_cell_wire[919];							inform_R[716][9] = r_cell_wire[920];							inform_R[972][9] = r_cell_wire[921];							inform_R[717][9] = r_cell_wire[922];							inform_R[973][9] = r_cell_wire[923];							inform_R[718][9] = r_cell_wire[924];							inform_R[974][9] = r_cell_wire[925];							inform_R[719][9] = r_cell_wire[926];							inform_R[975][9] = r_cell_wire[927];							inform_R[720][9] = r_cell_wire[928];							inform_R[976][9] = r_cell_wire[929];							inform_R[721][9] = r_cell_wire[930];							inform_R[977][9] = r_cell_wire[931];							inform_R[722][9] = r_cell_wire[932];							inform_R[978][9] = r_cell_wire[933];							inform_R[723][9] = r_cell_wire[934];							inform_R[979][9] = r_cell_wire[935];							inform_R[724][9] = r_cell_wire[936];							inform_R[980][9] = r_cell_wire[937];							inform_R[725][9] = r_cell_wire[938];							inform_R[981][9] = r_cell_wire[939];							inform_R[726][9] = r_cell_wire[940];							inform_R[982][9] = r_cell_wire[941];							inform_R[727][9] = r_cell_wire[942];							inform_R[983][9] = r_cell_wire[943];							inform_R[728][9] = r_cell_wire[944];							inform_R[984][9] = r_cell_wire[945];							inform_R[729][9] = r_cell_wire[946];							inform_R[985][9] = r_cell_wire[947];							inform_R[730][9] = r_cell_wire[948];							inform_R[986][9] = r_cell_wire[949];							inform_R[731][9] = r_cell_wire[950];							inform_R[987][9] = r_cell_wire[951];							inform_R[732][9] = r_cell_wire[952];							inform_R[988][9] = r_cell_wire[953];							inform_R[733][9] = r_cell_wire[954];							inform_R[989][9] = r_cell_wire[955];							inform_R[734][9] = r_cell_wire[956];							inform_R[990][9] = r_cell_wire[957];							inform_R[735][9] = r_cell_wire[958];							inform_R[991][9] = r_cell_wire[959];							inform_R[736][9] = r_cell_wire[960];							inform_R[992][9] = r_cell_wire[961];							inform_R[737][9] = r_cell_wire[962];							inform_R[993][9] = r_cell_wire[963];							inform_R[738][9] = r_cell_wire[964];							inform_R[994][9] = r_cell_wire[965];							inform_R[739][9] = r_cell_wire[966];							inform_R[995][9] = r_cell_wire[967];							inform_R[740][9] = r_cell_wire[968];							inform_R[996][9] = r_cell_wire[969];							inform_R[741][9] = r_cell_wire[970];							inform_R[997][9] = r_cell_wire[971];							inform_R[742][9] = r_cell_wire[972];							inform_R[998][9] = r_cell_wire[973];							inform_R[743][9] = r_cell_wire[974];							inform_R[999][9] = r_cell_wire[975];							inform_R[744][9] = r_cell_wire[976];							inform_R[1000][9] = r_cell_wire[977];							inform_R[745][9] = r_cell_wire[978];							inform_R[1001][9] = r_cell_wire[979];							inform_R[746][9] = r_cell_wire[980];							inform_R[1002][9] = r_cell_wire[981];							inform_R[747][9] = r_cell_wire[982];							inform_R[1003][9] = r_cell_wire[983];							inform_R[748][9] = r_cell_wire[984];							inform_R[1004][9] = r_cell_wire[985];							inform_R[749][9] = r_cell_wire[986];							inform_R[1005][9] = r_cell_wire[987];							inform_R[750][9] = r_cell_wire[988];							inform_R[1006][9] = r_cell_wire[989];							inform_R[751][9] = r_cell_wire[990];							inform_R[1007][9] = r_cell_wire[991];							inform_R[752][9] = r_cell_wire[992];							inform_R[1008][9] = r_cell_wire[993];							inform_R[753][9] = r_cell_wire[994];							inform_R[1009][9] = r_cell_wire[995];							inform_R[754][9] = r_cell_wire[996];							inform_R[1010][9] = r_cell_wire[997];							inform_R[755][9] = r_cell_wire[998];							inform_R[1011][9] = r_cell_wire[999];							inform_R[756][9] = r_cell_wire[1000];							inform_R[1012][9] = r_cell_wire[1001];							inform_R[757][9] = r_cell_wire[1002];							inform_R[1013][9] = r_cell_wire[1003];							inform_R[758][9] = r_cell_wire[1004];							inform_R[1014][9] = r_cell_wire[1005];							inform_R[759][9] = r_cell_wire[1006];							inform_R[1015][9] = r_cell_wire[1007];							inform_R[760][9] = r_cell_wire[1008];							inform_R[1016][9] = r_cell_wire[1009];							inform_R[761][9] = r_cell_wire[1010];							inform_R[1017][9] = r_cell_wire[1011];							inform_R[762][9] = r_cell_wire[1012];							inform_R[1018][9] = r_cell_wire[1013];							inform_R[763][9] = r_cell_wire[1014];							inform_R[1019][9] = r_cell_wire[1015];							inform_R[764][9] = r_cell_wire[1016];							inform_R[1020][9] = r_cell_wire[1017];							inform_R[765][9] = r_cell_wire[1018];							inform_R[1021][9] = r_cell_wire[1019];							inform_R[766][9] = r_cell_wire[1020];							inform_R[1022][9] = r_cell_wire[1021];							inform_R[767][9] = r_cell_wire[1022];							inform_R[1023][9] = r_cell_wire[1023];							inform_L[0][8] = l_cell_wire[0];							inform_L[256][8] = l_cell_wire[1];							inform_L[1][8] = l_cell_wire[2];							inform_L[257][8] = l_cell_wire[3];							inform_L[2][8] = l_cell_wire[4];							inform_L[258][8] = l_cell_wire[5];							inform_L[3][8] = l_cell_wire[6];							inform_L[259][8] = l_cell_wire[7];							inform_L[4][8] = l_cell_wire[8];							inform_L[260][8] = l_cell_wire[9];							inform_L[5][8] = l_cell_wire[10];							inform_L[261][8] = l_cell_wire[11];							inform_L[6][8] = l_cell_wire[12];							inform_L[262][8] = l_cell_wire[13];							inform_L[7][8] = l_cell_wire[14];							inform_L[263][8] = l_cell_wire[15];							inform_L[8][8] = l_cell_wire[16];							inform_L[264][8] = l_cell_wire[17];							inform_L[9][8] = l_cell_wire[18];							inform_L[265][8] = l_cell_wire[19];							inform_L[10][8] = l_cell_wire[20];							inform_L[266][8] = l_cell_wire[21];							inform_L[11][8] = l_cell_wire[22];							inform_L[267][8] = l_cell_wire[23];							inform_L[12][8] = l_cell_wire[24];							inform_L[268][8] = l_cell_wire[25];							inform_L[13][8] = l_cell_wire[26];							inform_L[269][8] = l_cell_wire[27];							inform_L[14][8] = l_cell_wire[28];							inform_L[270][8] = l_cell_wire[29];							inform_L[15][8] = l_cell_wire[30];							inform_L[271][8] = l_cell_wire[31];							inform_L[16][8] = l_cell_wire[32];							inform_L[272][8] = l_cell_wire[33];							inform_L[17][8] = l_cell_wire[34];							inform_L[273][8] = l_cell_wire[35];							inform_L[18][8] = l_cell_wire[36];							inform_L[274][8] = l_cell_wire[37];							inform_L[19][8] = l_cell_wire[38];							inform_L[275][8] = l_cell_wire[39];							inform_L[20][8] = l_cell_wire[40];							inform_L[276][8] = l_cell_wire[41];							inform_L[21][8] = l_cell_wire[42];							inform_L[277][8] = l_cell_wire[43];							inform_L[22][8] = l_cell_wire[44];							inform_L[278][8] = l_cell_wire[45];							inform_L[23][8] = l_cell_wire[46];							inform_L[279][8] = l_cell_wire[47];							inform_L[24][8] = l_cell_wire[48];							inform_L[280][8] = l_cell_wire[49];							inform_L[25][8] = l_cell_wire[50];							inform_L[281][8] = l_cell_wire[51];							inform_L[26][8] = l_cell_wire[52];							inform_L[282][8] = l_cell_wire[53];							inform_L[27][8] = l_cell_wire[54];							inform_L[283][8] = l_cell_wire[55];							inform_L[28][8] = l_cell_wire[56];							inform_L[284][8] = l_cell_wire[57];							inform_L[29][8] = l_cell_wire[58];							inform_L[285][8] = l_cell_wire[59];							inform_L[30][8] = l_cell_wire[60];							inform_L[286][8] = l_cell_wire[61];							inform_L[31][8] = l_cell_wire[62];							inform_L[287][8] = l_cell_wire[63];							inform_L[32][8] = l_cell_wire[64];							inform_L[288][8] = l_cell_wire[65];							inform_L[33][8] = l_cell_wire[66];							inform_L[289][8] = l_cell_wire[67];							inform_L[34][8] = l_cell_wire[68];							inform_L[290][8] = l_cell_wire[69];							inform_L[35][8] = l_cell_wire[70];							inform_L[291][8] = l_cell_wire[71];							inform_L[36][8] = l_cell_wire[72];							inform_L[292][8] = l_cell_wire[73];							inform_L[37][8] = l_cell_wire[74];							inform_L[293][8] = l_cell_wire[75];							inform_L[38][8] = l_cell_wire[76];							inform_L[294][8] = l_cell_wire[77];							inform_L[39][8] = l_cell_wire[78];							inform_L[295][8] = l_cell_wire[79];							inform_L[40][8] = l_cell_wire[80];							inform_L[296][8] = l_cell_wire[81];							inform_L[41][8] = l_cell_wire[82];							inform_L[297][8] = l_cell_wire[83];							inform_L[42][8] = l_cell_wire[84];							inform_L[298][8] = l_cell_wire[85];							inform_L[43][8] = l_cell_wire[86];							inform_L[299][8] = l_cell_wire[87];							inform_L[44][8] = l_cell_wire[88];							inform_L[300][8] = l_cell_wire[89];							inform_L[45][8] = l_cell_wire[90];							inform_L[301][8] = l_cell_wire[91];							inform_L[46][8] = l_cell_wire[92];							inform_L[302][8] = l_cell_wire[93];							inform_L[47][8] = l_cell_wire[94];							inform_L[303][8] = l_cell_wire[95];							inform_L[48][8] = l_cell_wire[96];							inform_L[304][8] = l_cell_wire[97];							inform_L[49][8] = l_cell_wire[98];							inform_L[305][8] = l_cell_wire[99];							inform_L[50][8] = l_cell_wire[100];							inform_L[306][8] = l_cell_wire[101];							inform_L[51][8] = l_cell_wire[102];							inform_L[307][8] = l_cell_wire[103];							inform_L[52][8] = l_cell_wire[104];							inform_L[308][8] = l_cell_wire[105];							inform_L[53][8] = l_cell_wire[106];							inform_L[309][8] = l_cell_wire[107];							inform_L[54][8] = l_cell_wire[108];							inform_L[310][8] = l_cell_wire[109];							inform_L[55][8] = l_cell_wire[110];							inform_L[311][8] = l_cell_wire[111];							inform_L[56][8] = l_cell_wire[112];							inform_L[312][8] = l_cell_wire[113];							inform_L[57][8] = l_cell_wire[114];							inform_L[313][8] = l_cell_wire[115];							inform_L[58][8] = l_cell_wire[116];							inform_L[314][8] = l_cell_wire[117];							inform_L[59][8] = l_cell_wire[118];							inform_L[315][8] = l_cell_wire[119];							inform_L[60][8] = l_cell_wire[120];							inform_L[316][8] = l_cell_wire[121];							inform_L[61][8] = l_cell_wire[122];							inform_L[317][8] = l_cell_wire[123];							inform_L[62][8] = l_cell_wire[124];							inform_L[318][8] = l_cell_wire[125];							inform_L[63][8] = l_cell_wire[126];							inform_L[319][8] = l_cell_wire[127];							inform_L[64][8] = l_cell_wire[128];							inform_L[320][8] = l_cell_wire[129];							inform_L[65][8] = l_cell_wire[130];							inform_L[321][8] = l_cell_wire[131];							inform_L[66][8] = l_cell_wire[132];							inform_L[322][8] = l_cell_wire[133];							inform_L[67][8] = l_cell_wire[134];							inform_L[323][8] = l_cell_wire[135];							inform_L[68][8] = l_cell_wire[136];							inform_L[324][8] = l_cell_wire[137];							inform_L[69][8] = l_cell_wire[138];							inform_L[325][8] = l_cell_wire[139];							inform_L[70][8] = l_cell_wire[140];							inform_L[326][8] = l_cell_wire[141];							inform_L[71][8] = l_cell_wire[142];							inform_L[327][8] = l_cell_wire[143];							inform_L[72][8] = l_cell_wire[144];							inform_L[328][8] = l_cell_wire[145];							inform_L[73][8] = l_cell_wire[146];							inform_L[329][8] = l_cell_wire[147];							inform_L[74][8] = l_cell_wire[148];							inform_L[330][8] = l_cell_wire[149];							inform_L[75][8] = l_cell_wire[150];							inform_L[331][8] = l_cell_wire[151];							inform_L[76][8] = l_cell_wire[152];							inform_L[332][8] = l_cell_wire[153];							inform_L[77][8] = l_cell_wire[154];							inform_L[333][8] = l_cell_wire[155];							inform_L[78][8] = l_cell_wire[156];							inform_L[334][8] = l_cell_wire[157];							inform_L[79][8] = l_cell_wire[158];							inform_L[335][8] = l_cell_wire[159];							inform_L[80][8] = l_cell_wire[160];							inform_L[336][8] = l_cell_wire[161];							inform_L[81][8] = l_cell_wire[162];							inform_L[337][8] = l_cell_wire[163];							inform_L[82][8] = l_cell_wire[164];							inform_L[338][8] = l_cell_wire[165];							inform_L[83][8] = l_cell_wire[166];							inform_L[339][8] = l_cell_wire[167];							inform_L[84][8] = l_cell_wire[168];							inform_L[340][8] = l_cell_wire[169];							inform_L[85][8] = l_cell_wire[170];							inform_L[341][8] = l_cell_wire[171];							inform_L[86][8] = l_cell_wire[172];							inform_L[342][8] = l_cell_wire[173];							inform_L[87][8] = l_cell_wire[174];							inform_L[343][8] = l_cell_wire[175];							inform_L[88][8] = l_cell_wire[176];							inform_L[344][8] = l_cell_wire[177];							inform_L[89][8] = l_cell_wire[178];							inform_L[345][8] = l_cell_wire[179];							inform_L[90][8] = l_cell_wire[180];							inform_L[346][8] = l_cell_wire[181];							inform_L[91][8] = l_cell_wire[182];							inform_L[347][8] = l_cell_wire[183];							inform_L[92][8] = l_cell_wire[184];							inform_L[348][8] = l_cell_wire[185];							inform_L[93][8] = l_cell_wire[186];							inform_L[349][8] = l_cell_wire[187];							inform_L[94][8] = l_cell_wire[188];							inform_L[350][8] = l_cell_wire[189];							inform_L[95][8] = l_cell_wire[190];							inform_L[351][8] = l_cell_wire[191];							inform_L[96][8] = l_cell_wire[192];							inform_L[352][8] = l_cell_wire[193];							inform_L[97][8] = l_cell_wire[194];							inform_L[353][8] = l_cell_wire[195];							inform_L[98][8] = l_cell_wire[196];							inform_L[354][8] = l_cell_wire[197];							inform_L[99][8] = l_cell_wire[198];							inform_L[355][8] = l_cell_wire[199];							inform_L[100][8] = l_cell_wire[200];							inform_L[356][8] = l_cell_wire[201];							inform_L[101][8] = l_cell_wire[202];							inform_L[357][8] = l_cell_wire[203];							inform_L[102][8] = l_cell_wire[204];							inform_L[358][8] = l_cell_wire[205];							inform_L[103][8] = l_cell_wire[206];							inform_L[359][8] = l_cell_wire[207];							inform_L[104][8] = l_cell_wire[208];							inform_L[360][8] = l_cell_wire[209];							inform_L[105][8] = l_cell_wire[210];							inform_L[361][8] = l_cell_wire[211];							inform_L[106][8] = l_cell_wire[212];							inform_L[362][8] = l_cell_wire[213];							inform_L[107][8] = l_cell_wire[214];							inform_L[363][8] = l_cell_wire[215];							inform_L[108][8] = l_cell_wire[216];							inform_L[364][8] = l_cell_wire[217];							inform_L[109][8] = l_cell_wire[218];							inform_L[365][8] = l_cell_wire[219];							inform_L[110][8] = l_cell_wire[220];							inform_L[366][8] = l_cell_wire[221];							inform_L[111][8] = l_cell_wire[222];							inform_L[367][8] = l_cell_wire[223];							inform_L[112][8] = l_cell_wire[224];							inform_L[368][8] = l_cell_wire[225];							inform_L[113][8] = l_cell_wire[226];							inform_L[369][8] = l_cell_wire[227];							inform_L[114][8] = l_cell_wire[228];							inform_L[370][8] = l_cell_wire[229];							inform_L[115][8] = l_cell_wire[230];							inform_L[371][8] = l_cell_wire[231];							inform_L[116][8] = l_cell_wire[232];							inform_L[372][8] = l_cell_wire[233];							inform_L[117][8] = l_cell_wire[234];							inform_L[373][8] = l_cell_wire[235];							inform_L[118][8] = l_cell_wire[236];							inform_L[374][8] = l_cell_wire[237];							inform_L[119][8] = l_cell_wire[238];							inform_L[375][8] = l_cell_wire[239];							inform_L[120][8] = l_cell_wire[240];							inform_L[376][8] = l_cell_wire[241];							inform_L[121][8] = l_cell_wire[242];							inform_L[377][8] = l_cell_wire[243];							inform_L[122][8] = l_cell_wire[244];							inform_L[378][8] = l_cell_wire[245];							inform_L[123][8] = l_cell_wire[246];							inform_L[379][8] = l_cell_wire[247];							inform_L[124][8] = l_cell_wire[248];							inform_L[380][8] = l_cell_wire[249];							inform_L[125][8] = l_cell_wire[250];							inform_L[381][8] = l_cell_wire[251];							inform_L[126][8] = l_cell_wire[252];							inform_L[382][8] = l_cell_wire[253];							inform_L[127][8] = l_cell_wire[254];							inform_L[383][8] = l_cell_wire[255];							inform_L[128][8] = l_cell_wire[256];							inform_L[384][8] = l_cell_wire[257];							inform_L[129][8] = l_cell_wire[258];							inform_L[385][8] = l_cell_wire[259];							inform_L[130][8] = l_cell_wire[260];							inform_L[386][8] = l_cell_wire[261];							inform_L[131][8] = l_cell_wire[262];							inform_L[387][8] = l_cell_wire[263];							inform_L[132][8] = l_cell_wire[264];							inform_L[388][8] = l_cell_wire[265];							inform_L[133][8] = l_cell_wire[266];							inform_L[389][8] = l_cell_wire[267];							inform_L[134][8] = l_cell_wire[268];							inform_L[390][8] = l_cell_wire[269];							inform_L[135][8] = l_cell_wire[270];							inform_L[391][8] = l_cell_wire[271];							inform_L[136][8] = l_cell_wire[272];							inform_L[392][8] = l_cell_wire[273];							inform_L[137][8] = l_cell_wire[274];							inform_L[393][8] = l_cell_wire[275];							inform_L[138][8] = l_cell_wire[276];							inform_L[394][8] = l_cell_wire[277];							inform_L[139][8] = l_cell_wire[278];							inform_L[395][8] = l_cell_wire[279];							inform_L[140][8] = l_cell_wire[280];							inform_L[396][8] = l_cell_wire[281];							inform_L[141][8] = l_cell_wire[282];							inform_L[397][8] = l_cell_wire[283];							inform_L[142][8] = l_cell_wire[284];							inform_L[398][8] = l_cell_wire[285];							inform_L[143][8] = l_cell_wire[286];							inform_L[399][8] = l_cell_wire[287];							inform_L[144][8] = l_cell_wire[288];							inform_L[400][8] = l_cell_wire[289];							inform_L[145][8] = l_cell_wire[290];							inform_L[401][8] = l_cell_wire[291];							inform_L[146][8] = l_cell_wire[292];							inform_L[402][8] = l_cell_wire[293];							inform_L[147][8] = l_cell_wire[294];							inform_L[403][8] = l_cell_wire[295];							inform_L[148][8] = l_cell_wire[296];							inform_L[404][8] = l_cell_wire[297];							inform_L[149][8] = l_cell_wire[298];							inform_L[405][8] = l_cell_wire[299];							inform_L[150][8] = l_cell_wire[300];							inform_L[406][8] = l_cell_wire[301];							inform_L[151][8] = l_cell_wire[302];							inform_L[407][8] = l_cell_wire[303];							inform_L[152][8] = l_cell_wire[304];							inform_L[408][8] = l_cell_wire[305];							inform_L[153][8] = l_cell_wire[306];							inform_L[409][8] = l_cell_wire[307];							inform_L[154][8] = l_cell_wire[308];							inform_L[410][8] = l_cell_wire[309];							inform_L[155][8] = l_cell_wire[310];							inform_L[411][8] = l_cell_wire[311];							inform_L[156][8] = l_cell_wire[312];							inform_L[412][8] = l_cell_wire[313];							inform_L[157][8] = l_cell_wire[314];							inform_L[413][8] = l_cell_wire[315];							inform_L[158][8] = l_cell_wire[316];							inform_L[414][8] = l_cell_wire[317];							inform_L[159][8] = l_cell_wire[318];							inform_L[415][8] = l_cell_wire[319];							inform_L[160][8] = l_cell_wire[320];							inform_L[416][8] = l_cell_wire[321];							inform_L[161][8] = l_cell_wire[322];							inform_L[417][8] = l_cell_wire[323];							inform_L[162][8] = l_cell_wire[324];							inform_L[418][8] = l_cell_wire[325];							inform_L[163][8] = l_cell_wire[326];							inform_L[419][8] = l_cell_wire[327];							inform_L[164][8] = l_cell_wire[328];							inform_L[420][8] = l_cell_wire[329];							inform_L[165][8] = l_cell_wire[330];							inform_L[421][8] = l_cell_wire[331];							inform_L[166][8] = l_cell_wire[332];							inform_L[422][8] = l_cell_wire[333];							inform_L[167][8] = l_cell_wire[334];							inform_L[423][8] = l_cell_wire[335];							inform_L[168][8] = l_cell_wire[336];							inform_L[424][8] = l_cell_wire[337];							inform_L[169][8] = l_cell_wire[338];							inform_L[425][8] = l_cell_wire[339];							inform_L[170][8] = l_cell_wire[340];							inform_L[426][8] = l_cell_wire[341];							inform_L[171][8] = l_cell_wire[342];							inform_L[427][8] = l_cell_wire[343];							inform_L[172][8] = l_cell_wire[344];							inform_L[428][8] = l_cell_wire[345];							inform_L[173][8] = l_cell_wire[346];							inform_L[429][8] = l_cell_wire[347];							inform_L[174][8] = l_cell_wire[348];							inform_L[430][8] = l_cell_wire[349];							inform_L[175][8] = l_cell_wire[350];							inform_L[431][8] = l_cell_wire[351];							inform_L[176][8] = l_cell_wire[352];							inform_L[432][8] = l_cell_wire[353];							inform_L[177][8] = l_cell_wire[354];							inform_L[433][8] = l_cell_wire[355];							inform_L[178][8] = l_cell_wire[356];							inform_L[434][8] = l_cell_wire[357];							inform_L[179][8] = l_cell_wire[358];							inform_L[435][8] = l_cell_wire[359];							inform_L[180][8] = l_cell_wire[360];							inform_L[436][8] = l_cell_wire[361];							inform_L[181][8] = l_cell_wire[362];							inform_L[437][8] = l_cell_wire[363];							inform_L[182][8] = l_cell_wire[364];							inform_L[438][8] = l_cell_wire[365];							inform_L[183][8] = l_cell_wire[366];							inform_L[439][8] = l_cell_wire[367];							inform_L[184][8] = l_cell_wire[368];							inform_L[440][8] = l_cell_wire[369];							inform_L[185][8] = l_cell_wire[370];							inform_L[441][8] = l_cell_wire[371];							inform_L[186][8] = l_cell_wire[372];							inform_L[442][8] = l_cell_wire[373];							inform_L[187][8] = l_cell_wire[374];							inform_L[443][8] = l_cell_wire[375];							inform_L[188][8] = l_cell_wire[376];							inform_L[444][8] = l_cell_wire[377];							inform_L[189][8] = l_cell_wire[378];							inform_L[445][8] = l_cell_wire[379];							inform_L[190][8] = l_cell_wire[380];							inform_L[446][8] = l_cell_wire[381];							inform_L[191][8] = l_cell_wire[382];							inform_L[447][8] = l_cell_wire[383];							inform_L[192][8] = l_cell_wire[384];							inform_L[448][8] = l_cell_wire[385];							inform_L[193][8] = l_cell_wire[386];							inform_L[449][8] = l_cell_wire[387];							inform_L[194][8] = l_cell_wire[388];							inform_L[450][8] = l_cell_wire[389];							inform_L[195][8] = l_cell_wire[390];							inform_L[451][8] = l_cell_wire[391];							inform_L[196][8] = l_cell_wire[392];							inform_L[452][8] = l_cell_wire[393];							inform_L[197][8] = l_cell_wire[394];							inform_L[453][8] = l_cell_wire[395];							inform_L[198][8] = l_cell_wire[396];							inform_L[454][8] = l_cell_wire[397];							inform_L[199][8] = l_cell_wire[398];							inform_L[455][8] = l_cell_wire[399];							inform_L[200][8] = l_cell_wire[400];							inform_L[456][8] = l_cell_wire[401];							inform_L[201][8] = l_cell_wire[402];							inform_L[457][8] = l_cell_wire[403];							inform_L[202][8] = l_cell_wire[404];							inform_L[458][8] = l_cell_wire[405];							inform_L[203][8] = l_cell_wire[406];							inform_L[459][8] = l_cell_wire[407];							inform_L[204][8] = l_cell_wire[408];							inform_L[460][8] = l_cell_wire[409];							inform_L[205][8] = l_cell_wire[410];							inform_L[461][8] = l_cell_wire[411];							inform_L[206][8] = l_cell_wire[412];							inform_L[462][8] = l_cell_wire[413];							inform_L[207][8] = l_cell_wire[414];							inform_L[463][8] = l_cell_wire[415];							inform_L[208][8] = l_cell_wire[416];							inform_L[464][8] = l_cell_wire[417];							inform_L[209][8] = l_cell_wire[418];							inform_L[465][8] = l_cell_wire[419];							inform_L[210][8] = l_cell_wire[420];							inform_L[466][8] = l_cell_wire[421];							inform_L[211][8] = l_cell_wire[422];							inform_L[467][8] = l_cell_wire[423];							inform_L[212][8] = l_cell_wire[424];							inform_L[468][8] = l_cell_wire[425];							inform_L[213][8] = l_cell_wire[426];							inform_L[469][8] = l_cell_wire[427];							inform_L[214][8] = l_cell_wire[428];							inform_L[470][8] = l_cell_wire[429];							inform_L[215][8] = l_cell_wire[430];							inform_L[471][8] = l_cell_wire[431];							inform_L[216][8] = l_cell_wire[432];							inform_L[472][8] = l_cell_wire[433];							inform_L[217][8] = l_cell_wire[434];							inform_L[473][8] = l_cell_wire[435];							inform_L[218][8] = l_cell_wire[436];							inform_L[474][8] = l_cell_wire[437];							inform_L[219][8] = l_cell_wire[438];							inform_L[475][8] = l_cell_wire[439];							inform_L[220][8] = l_cell_wire[440];							inform_L[476][8] = l_cell_wire[441];							inform_L[221][8] = l_cell_wire[442];							inform_L[477][8] = l_cell_wire[443];							inform_L[222][8] = l_cell_wire[444];							inform_L[478][8] = l_cell_wire[445];							inform_L[223][8] = l_cell_wire[446];							inform_L[479][8] = l_cell_wire[447];							inform_L[224][8] = l_cell_wire[448];							inform_L[480][8] = l_cell_wire[449];							inform_L[225][8] = l_cell_wire[450];							inform_L[481][8] = l_cell_wire[451];							inform_L[226][8] = l_cell_wire[452];							inform_L[482][8] = l_cell_wire[453];							inform_L[227][8] = l_cell_wire[454];							inform_L[483][8] = l_cell_wire[455];							inform_L[228][8] = l_cell_wire[456];							inform_L[484][8] = l_cell_wire[457];							inform_L[229][8] = l_cell_wire[458];							inform_L[485][8] = l_cell_wire[459];							inform_L[230][8] = l_cell_wire[460];							inform_L[486][8] = l_cell_wire[461];							inform_L[231][8] = l_cell_wire[462];							inform_L[487][8] = l_cell_wire[463];							inform_L[232][8] = l_cell_wire[464];							inform_L[488][8] = l_cell_wire[465];							inform_L[233][8] = l_cell_wire[466];							inform_L[489][8] = l_cell_wire[467];							inform_L[234][8] = l_cell_wire[468];							inform_L[490][8] = l_cell_wire[469];							inform_L[235][8] = l_cell_wire[470];							inform_L[491][8] = l_cell_wire[471];							inform_L[236][8] = l_cell_wire[472];							inform_L[492][8] = l_cell_wire[473];							inform_L[237][8] = l_cell_wire[474];							inform_L[493][8] = l_cell_wire[475];							inform_L[238][8] = l_cell_wire[476];							inform_L[494][8] = l_cell_wire[477];							inform_L[239][8] = l_cell_wire[478];							inform_L[495][8] = l_cell_wire[479];							inform_L[240][8] = l_cell_wire[480];							inform_L[496][8] = l_cell_wire[481];							inform_L[241][8] = l_cell_wire[482];							inform_L[497][8] = l_cell_wire[483];							inform_L[242][8] = l_cell_wire[484];							inform_L[498][8] = l_cell_wire[485];							inform_L[243][8] = l_cell_wire[486];							inform_L[499][8] = l_cell_wire[487];							inform_L[244][8] = l_cell_wire[488];							inform_L[500][8] = l_cell_wire[489];							inform_L[245][8] = l_cell_wire[490];							inform_L[501][8] = l_cell_wire[491];							inform_L[246][8] = l_cell_wire[492];							inform_L[502][8] = l_cell_wire[493];							inform_L[247][8] = l_cell_wire[494];							inform_L[503][8] = l_cell_wire[495];							inform_L[248][8] = l_cell_wire[496];							inform_L[504][8] = l_cell_wire[497];							inform_L[249][8] = l_cell_wire[498];							inform_L[505][8] = l_cell_wire[499];							inform_L[250][8] = l_cell_wire[500];							inform_L[506][8] = l_cell_wire[501];							inform_L[251][8] = l_cell_wire[502];							inform_L[507][8] = l_cell_wire[503];							inform_L[252][8] = l_cell_wire[504];							inform_L[508][8] = l_cell_wire[505];							inform_L[253][8] = l_cell_wire[506];							inform_L[509][8] = l_cell_wire[507];							inform_L[254][8] = l_cell_wire[508];							inform_L[510][8] = l_cell_wire[509];							inform_L[255][8] = l_cell_wire[510];							inform_L[511][8] = l_cell_wire[511];							inform_L[512][8] = l_cell_wire[512];							inform_L[768][8] = l_cell_wire[513];							inform_L[513][8] = l_cell_wire[514];							inform_L[769][8] = l_cell_wire[515];							inform_L[514][8] = l_cell_wire[516];							inform_L[770][8] = l_cell_wire[517];							inform_L[515][8] = l_cell_wire[518];							inform_L[771][8] = l_cell_wire[519];							inform_L[516][8] = l_cell_wire[520];							inform_L[772][8] = l_cell_wire[521];							inform_L[517][8] = l_cell_wire[522];							inform_L[773][8] = l_cell_wire[523];							inform_L[518][8] = l_cell_wire[524];							inform_L[774][8] = l_cell_wire[525];							inform_L[519][8] = l_cell_wire[526];							inform_L[775][8] = l_cell_wire[527];							inform_L[520][8] = l_cell_wire[528];							inform_L[776][8] = l_cell_wire[529];							inform_L[521][8] = l_cell_wire[530];							inform_L[777][8] = l_cell_wire[531];							inform_L[522][8] = l_cell_wire[532];							inform_L[778][8] = l_cell_wire[533];							inform_L[523][8] = l_cell_wire[534];							inform_L[779][8] = l_cell_wire[535];							inform_L[524][8] = l_cell_wire[536];							inform_L[780][8] = l_cell_wire[537];							inform_L[525][8] = l_cell_wire[538];							inform_L[781][8] = l_cell_wire[539];							inform_L[526][8] = l_cell_wire[540];							inform_L[782][8] = l_cell_wire[541];							inform_L[527][8] = l_cell_wire[542];							inform_L[783][8] = l_cell_wire[543];							inform_L[528][8] = l_cell_wire[544];							inform_L[784][8] = l_cell_wire[545];							inform_L[529][8] = l_cell_wire[546];							inform_L[785][8] = l_cell_wire[547];							inform_L[530][8] = l_cell_wire[548];							inform_L[786][8] = l_cell_wire[549];							inform_L[531][8] = l_cell_wire[550];							inform_L[787][8] = l_cell_wire[551];							inform_L[532][8] = l_cell_wire[552];							inform_L[788][8] = l_cell_wire[553];							inform_L[533][8] = l_cell_wire[554];							inform_L[789][8] = l_cell_wire[555];							inform_L[534][8] = l_cell_wire[556];							inform_L[790][8] = l_cell_wire[557];							inform_L[535][8] = l_cell_wire[558];							inform_L[791][8] = l_cell_wire[559];							inform_L[536][8] = l_cell_wire[560];							inform_L[792][8] = l_cell_wire[561];							inform_L[537][8] = l_cell_wire[562];							inform_L[793][8] = l_cell_wire[563];							inform_L[538][8] = l_cell_wire[564];							inform_L[794][8] = l_cell_wire[565];							inform_L[539][8] = l_cell_wire[566];							inform_L[795][8] = l_cell_wire[567];							inform_L[540][8] = l_cell_wire[568];							inform_L[796][8] = l_cell_wire[569];							inform_L[541][8] = l_cell_wire[570];							inform_L[797][8] = l_cell_wire[571];							inform_L[542][8] = l_cell_wire[572];							inform_L[798][8] = l_cell_wire[573];							inform_L[543][8] = l_cell_wire[574];							inform_L[799][8] = l_cell_wire[575];							inform_L[544][8] = l_cell_wire[576];							inform_L[800][8] = l_cell_wire[577];							inform_L[545][8] = l_cell_wire[578];							inform_L[801][8] = l_cell_wire[579];							inform_L[546][8] = l_cell_wire[580];							inform_L[802][8] = l_cell_wire[581];							inform_L[547][8] = l_cell_wire[582];							inform_L[803][8] = l_cell_wire[583];							inform_L[548][8] = l_cell_wire[584];							inform_L[804][8] = l_cell_wire[585];							inform_L[549][8] = l_cell_wire[586];							inform_L[805][8] = l_cell_wire[587];							inform_L[550][8] = l_cell_wire[588];							inform_L[806][8] = l_cell_wire[589];							inform_L[551][8] = l_cell_wire[590];							inform_L[807][8] = l_cell_wire[591];							inform_L[552][8] = l_cell_wire[592];							inform_L[808][8] = l_cell_wire[593];							inform_L[553][8] = l_cell_wire[594];							inform_L[809][8] = l_cell_wire[595];							inform_L[554][8] = l_cell_wire[596];							inform_L[810][8] = l_cell_wire[597];							inform_L[555][8] = l_cell_wire[598];							inform_L[811][8] = l_cell_wire[599];							inform_L[556][8] = l_cell_wire[600];							inform_L[812][8] = l_cell_wire[601];							inform_L[557][8] = l_cell_wire[602];							inform_L[813][8] = l_cell_wire[603];							inform_L[558][8] = l_cell_wire[604];							inform_L[814][8] = l_cell_wire[605];							inform_L[559][8] = l_cell_wire[606];							inform_L[815][8] = l_cell_wire[607];							inform_L[560][8] = l_cell_wire[608];							inform_L[816][8] = l_cell_wire[609];							inform_L[561][8] = l_cell_wire[610];							inform_L[817][8] = l_cell_wire[611];							inform_L[562][8] = l_cell_wire[612];							inform_L[818][8] = l_cell_wire[613];							inform_L[563][8] = l_cell_wire[614];							inform_L[819][8] = l_cell_wire[615];							inform_L[564][8] = l_cell_wire[616];							inform_L[820][8] = l_cell_wire[617];							inform_L[565][8] = l_cell_wire[618];							inform_L[821][8] = l_cell_wire[619];							inform_L[566][8] = l_cell_wire[620];							inform_L[822][8] = l_cell_wire[621];							inform_L[567][8] = l_cell_wire[622];							inform_L[823][8] = l_cell_wire[623];							inform_L[568][8] = l_cell_wire[624];							inform_L[824][8] = l_cell_wire[625];							inform_L[569][8] = l_cell_wire[626];							inform_L[825][8] = l_cell_wire[627];							inform_L[570][8] = l_cell_wire[628];							inform_L[826][8] = l_cell_wire[629];							inform_L[571][8] = l_cell_wire[630];							inform_L[827][8] = l_cell_wire[631];							inform_L[572][8] = l_cell_wire[632];							inform_L[828][8] = l_cell_wire[633];							inform_L[573][8] = l_cell_wire[634];							inform_L[829][8] = l_cell_wire[635];							inform_L[574][8] = l_cell_wire[636];							inform_L[830][8] = l_cell_wire[637];							inform_L[575][8] = l_cell_wire[638];							inform_L[831][8] = l_cell_wire[639];							inform_L[576][8] = l_cell_wire[640];							inform_L[832][8] = l_cell_wire[641];							inform_L[577][8] = l_cell_wire[642];							inform_L[833][8] = l_cell_wire[643];							inform_L[578][8] = l_cell_wire[644];							inform_L[834][8] = l_cell_wire[645];							inform_L[579][8] = l_cell_wire[646];							inform_L[835][8] = l_cell_wire[647];							inform_L[580][8] = l_cell_wire[648];							inform_L[836][8] = l_cell_wire[649];							inform_L[581][8] = l_cell_wire[650];							inform_L[837][8] = l_cell_wire[651];							inform_L[582][8] = l_cell_wire[652];							inform_L[838][8] = l_cell_wire[653];							inform_L[583][8] = l_cell_wire[654];							inform_L[839][8] = l_cell_wire[655];							inform_L[584][8] = l_cell_wire[656];							inform_L[840][8] = l_cell_wire[657];							inform_L[585][8] = l_cell_wire[658];							inform_L[841][8] = l_cell_wire[659];							inform_L[586][8] = l_cell_wire[660];							inform_L[842][8] = l_cell_wire[661];							inform_L[587][8] = l_cell_wire[662];							inform_L[843][8] = l_cell_wire[663];							inform_L[588][8] = l_cell_wire[664];							inform_L[844][8] = l_cell_wire[665];							inform_L[589][8] = l_cell_wire[666];							inform_L[845][8] = l_cell_wire[667];							inform_L[590][8] = l_cell_wire[668];							inform_L[846][8] = l_cell_wire[669];							inform_L[591][8] = l_cell_wire[670];							inform_L[847][8] = l_cell_wire[671];							inform_L[592][8] = l_cell_wire[672];							inform_L[848][8] = l_cell_wire[673];							inform_L[593][8] = l_cell_wire[674];							inform_L[849][8] = l_cell_wire[675];							inform_L[594][8] = l_cell_wire[676];							inform_L[850][8] = l_cell_wire[677];							inform_L[595][8] = l_cell_wire[678];							inform_L[851][8] = l_cell_wire[679];							inform_L[596][8] = l_cell_wire[680];							inform_L[852][8] = l_cell_wire[681];							inform_L[597][8] = l_cell_wire[682];							inform_L[853][8] = l_cell_wire[683];							inform_L[598][8] = l_cell_wire[684];							inform_L[854][8] = l_cell_wire[685];							inform_L[599][8] = l_cell_wire[686];							inform_L[855][8] = l_cell_wire[687];							inform_L[600][8] = l_cell_wire[688];							inform_L[856][8] = l_cell_wire[689];							inform_L[601][8] = l_cell_wire[690];							inform_L[857][8] = l_cell_wire[691];							inform_L[602][8] = l_cell_wire[692];							inform_L[858][8] = l_cell_wire[693];							inform_L[603][8] = l_cell_wire[694];							inform_L[859][8] = l_cell_wire[695];							inform_L[604][8] = l_cell_wire[696];							inform_L[860][8] = l_cell_wire[697];							inform_L[605][8] = l_cell_wire[698];							inform_L[861][8] = l_cell_wire[699];							inform_L[606][8] = l_cell_wire[700];							inform_L[862][8] = l_cell_wire[701];							inform_L[607][8] = l_cell_wire[702];							inform_L[863][8] = l_cell_wire[703];							inform_L[608][8] = l_cell_wire[704];							inform_L[864][8] = l_cell_wire[705];							inform_L[609][8] = l_cell_wire[706];							inform_L[865][8] = l_cell_wire[707];							inform_L[610][8] = l_cell_wire[708];							inform_L[866][8] = l_cell_wire[709];							inform_L[611][8] = l_cell_wire[710];							inform_L[867][8] = l_cell_wire[711];							inform_L[612][8] = l_cell_wire[712];							inform_L[868][8] = l_cell_wire[713];							inform_L[613][8] = l_cell_wire[714];							inform_L[869][8] = l_cell_wire[715];							inform_L[614][8] = l_cell_wire[716];							inform_L[870][8] = l_cell_wire[717];							inform_L[615][8] = l_cell_wire[718];							inform_L[871][8] = l_cell_wire[719];							inform_L[616][8] = l_cell_wire[720];							inform_L[872][8] = l_cell_wire[721];							inform_L[617][8] = l_cell_wire[722];							inform_L[873][8] = l_cell_wire[723];							inform_L[618][8] = l_cell_wire[724];							inform_L[874][8] = l_cell_wire[725];							inform_L[619][8] = l_cell_wire[726];							inform_L[875][8] = l_cell_wire[727];							inform_L[620][8] = l_cell_wire[728];							inform_L[876][8] = l_cell_wire[729];							inform_L[621][8] = l_cell_wire[730];							inform_L[877][8] = l_cell_wire[731];							inform_L[622][8] = l_cell_wire[732];							inform_L[878][8] = l_cell_wire[733];							inform_L[623][8] = l_cell_wire[734];							inform_L[879][8] = l_cell_wire[735];							inform_L[624][8] = l_cell_wire[736];							inform_L[880][8] = l_cell_wire[737];							inform_L[625][8] = l_cell_wire[738];							inform_L[881][8] = l_cell_wire[739];							inform_L[626][8] = l_cell_wire[740];							inform_L[882][8] = l_cell_wire[741];							inform_L[627][8] = l_cell_wire[742];							inform_L[883][8] = l_cell_wire[743];							inform_L[628][8] = l_cell_wire[744];							inform_L[884][8] = l_cell_wire[745];							inform_L[629][8] = l_cell_wire[746];							inform_L[885][8] = l_cell_wire[747];							inform_L[630][8] = l_cell_wire[748];							inform_L[886][8] = l_cell_wire[749];							inform_L[631][8] = l_cell_wire[750];							inform_L[887][8] = l_cell_wire[751];							inform_L[632][8] = l_cell_wire[752];							inform_L[888][8] = l_cell_wire[753];							inform_L[633][8] = l_cell_wire[754];							inform_L[889][8] = l_cell_wire[755];							inform_L[634][8] = l_cell_wire[756];							inform_L[890][8] = l_cell_wire[757];							inform_L[635][8] = l_cell_wire[758];							inform_L[891][8] = l_cell_wire[759];							inform_L[636][8] = l_cell_wire[760];							inform_L[892][8] = l_cell_wire[761];							inform_L[637][8] = l_cell_wire[762];							inform_L[893][8] = l_cell_wire[763];							inform_L[638][8] = l_cell_wire[764];							inform_L[894][8] = l_cell_wire[765];							inform_L[639][8] = l_cell_wire[766];							inform_L[895][8] = l_cell_wire[767];							inform_L[640][8] = l_cell_wire[768];							inform_L[896][8] = l_cell_wire[769];							inform_L[641][8] = l_cell_wire[770];							inform_L[897][8] = l_cell_wire[771];							inform_L[642][8] = l_cell_wire[772];							inform_L[898][8] = l_cell_wire[773];							inform_L[643][8] = l_cell_wire[774];							inform_L[899][8] = l_cell_wire[775];							inform_L[644][8] = l_cell_wire[776];							inform_L[900][8] = l_cell_wire[777];							inform_L[645][8] = l_cell_wire[778];							inform_L[901][8] = l_cell_wire[779];							inform_L[646][8] = l_cell_wire[780];							inform_L[902][8] = l_cell_wire[781];							inform_L[647][8] = l_cell_wire[782];							inform_L[903][8] = l_cell_wire[783];							inform_L[648][8] = l_cell_wire[784];							inform_L[904][8] = l_cell_wire[785];							inform_L[649][8] = l_cell_wire[786];							inform_L[905][8] = l_cell_wire[787];							inform_L[650][8] = l_cell_wire[788];							inform_L[906][8] = l_cell_wire[789];							inform_L[651][8] = l_cell_wire[790];							inform_L[907][8] = l_cell_wire[791];							inform_L[652][8] = l_cell_wire[792];							inform_L[908][8] = l_cell_wire[793];							inform_L[653][8] = l_cell_wire[794];							inform_L[909][8] = l_cell_wire[795];							inform_L[654][8] = l_cell_wire[796];							inform_L[910][8] = l_cell_wire[797];							inform_L[655][8] = l_cell_wire[798];							inform_L[911][8] = l_cell_wire[799];							inform_L[656][8] = l_cell_wire[800];							inform_L[912][8] = l_cell_wire[801];							inform_L[657][8] = l_cell_wire[802];							inform_L[913][8] = l_cell_wire[803];							inform_L[658][8] = l_cell_wire[804];							inform_L[914][8] = l_cell_wire[805];							inform_L[659][8] = l_cell_wire[806];							inform_L[915][8] = l_cell_wire[807];							inform_L[660][8] = l_cell_wire[808];							inform_L[916][8] = l_cell_wire[809];							inform_L[661][8] = l_cell_wire[810];							inform_L[917][8] = l_cell_wire[811];							inform_L[662][8] = l_cell_wire[812];							inform_L[918][8] = l_cell_wire[813];							inform_L[663][8] = l_cell_wire[814];							inform_L[919][8] = l_cell_wire[815];							inform_L[664][8] = l_cell_wire[816];							inform_L[920][8] = l_cell_wire[817];							inform_L[665][8] = l_cell_wire[818];							inform_L[921][8] = l_cell_wire[819];							inform_L[666][8] = l_cell_wire[820];							inform_L[922][8] = l_cell_wire[821];							inform_L[667][8] = l_cell_wire[822];							inform_L[923][8] = l_cell_wire[823];							inform_L[668][8] = l_cell_wire[824];							inform_L[924][8] = l_cell_wire[825];							inform_L[669][8] = l_cell_wire[826];							inform_L[925][8] = l_cell_wire[827];							inform_L[670][8] = l_cell_wire[828];							inform_L[926][8] = l_cell_wire[829];							inform_L[671][8] = l_cell_wire[830];							inform_L[927][8] = l_cell_wire[831];							inform_L[672][8] = l_cell_wire[832];							inform_L[928][8] = l_cell_wire[833];							inform_L[673][8] = l_cell_wire[834];							inform_L[929][8] = l_cell_wire[835];							inform_L[674][8] = l_cell_wire[836];							inform_L[930][8] = l_cell_wire[837];							inform_L[675][8] = l_cell_wire[838];							inform_L[931][8] = l_cell_wire[839];							inform_L[676][8] = l_cell_wire[840];							inform_L[932][8] = l_cell_wire[841];							inform_L[677][8] = l_cell_wire[842];							inform_L[933][8] = l_cell_wire[843];							inform_L[678][8] = l_cell_wire[844];							inform_L[934][8] = l_cell_wire[845];							inform_L[679][8] = l_cell_wire[846];							inform_L[935][8] = l_cell_wire[847];							inform_L[680][8] = l_cell_wire[848];							inform_L[936][8] = l_cell_wire[849];							inform_L[681][8] = l_cell_wire[850];							inform_L[937][8] = l_cell_wire[851];							inform_L[682][8] = l_cell_wire[852];							inform_L[938][8] = l_cell_wire[853];							inform_L[683][8] = l_cell_wire[854];							inform_L[939][8] = l_cell_wire[855];							inform_L[684][8] = l_cell_wire[856];							inform_L[940][8] = l_cell_wire[857];							inform_L[685][8] = l_cell_wire[858];							inform_L[941][8] = l_cell_wire[859];							inform_L[686][8] = l_cell_wire[860];							inform_L[942][8] = l_cell_wire[861];							inform_L[687][8] = l_cell_wire[862];							inform_L[943][8] = l_cell_wire[863];							inform_L[688][8] = l_cell_wire[864];							inform_L[944][8] = l_cell_wire[865];							inform_L[689][8] = l_cell_wire[866];							inform_L[945][8] = l_cell_wire[867];							inform_L[690][8] = l_cell_wire[868];							inform_L[946][8] = l_cell_wire[869];							inform_L[691][8] = l_cell_wire[870];							inform_L[947][8] = l_cell_wire[871];							inform_L[692][8] = l_cell_wire[872];							inform_L[948][8] = l_cell_wire[873];							inform_L[693][8] = l_cell_wire[874];							inform_L[949][8] = l_cell_wire[875];							inform_L[694][8] = l_cell_wire[876];							inform_L[950][8] = l_cell_wire[877];							inform_L[695][8] = l_cell_wire[878];							inform_L[951][8] = l_cell_wire[879];							inform_L[696][8] = l_cell_wire[880];							inform_L[952][8] = l_cell_wire[881];							inform_L[697][8] = l_cell_wire[882];							inform_L[953][8] = l_cell_wire[883];							inform_L[698][8] = l_cell_wire[884];							inform_L[954][8] = l_cell_wire[885];							inform_L[699][8] = l_cell_wire[886];							inform_L[955][8] = l_cell_wire[887];							inform_L[700][8] = l_cell_wire[888];							inform_L[956][8] = l_cell_wire[889];							inform_L[701][8] = l_cell_wire[890];							inform_L[957][8] = l_cell_wire[891];							inform_L[702][8] = l_cell_wire[892];							inform_L[958][8] = l_cell_wire[893];							inform_L[703][8] = l_cell_wire[894];							inform_L[959][8] = l_cell_wire[895];							inform_L[704][8] = l_cell_wire[896];							inform_L[960][8] = l_cell_wire[897];							inform_L[705][8] = l_cell_wire[898];							inform_L[961][8] = l_cell_wire[899];							inform_L[706][8] = l_cell_wire[900];							inform_L[962][8] = l_cell_wire[901];							inform_L[707][8] = l_cell_wire[902];							inform_L[963][8] = l_cell_wire[903];							inform_L[708][8] = l_cell_wire[904];							inform_L[964][8] = l_cell_wire[905];							inform_L[709][8] = l_cell_wire[906];							inform_L[965][8] = l_cell_wire[907];							inform_L[710][8] = l_cell_wire[908];							inform_L[966][8] = l_cell_wire[909];							inform_L[711][8] = l_cell_wire[910];							inform_L[967][8] = l_cell_wire[911];							inform_L[712][8] = l_cell_wire[912];							inform_L[968][8] = l_cell_wire[913];							inform_L[713][8] = l_cell_wire[914];							inform_L[969][8] = l_cell_wire[915];							inform_L[714][8] = l_cell_wire[916];							inform_L[970][8] = l_cell_wire[917];							inform_L[715][8] = l_cell_wire[918];							inform_L[971][8] = l_cell_wire[919];							inform_L[716][8] = l_cell_wire[920];							inform_L[972][8] = l_cell_wire[921];							inform_L[717][8] = l_cell_wire[922];							inform_L[973][8] = l_cell_wire[923];							inform_L[718][8] = l_cell_wire[924];							inform_L[974][8] = l_cell_wire[925];							inform_L[719][8] = l_cell_wire[926];							inform_L[975][8] = l_cell_wire[927];							inform_L[720][8] = l_cell_wire[928];							inform_L[976][8] = l_cell_wire[929];							inform_L[721][8] = l_cell_wire[930];							inform_L[977][8] = l_cell_wire[931];							inform_L[722][8] = l_cell_wire[932];							inform_L[978][8] = l_cell_wire[933];							inform_L[723][8] = l_cell_wire[934];							inform_L[979][8] = l_cell_wire[935];							inform_L[724][8] = l_cell_wire[936];							inform_L[980][8] = l_cell_wire[937];							inform_L[725][8] = l_cell_wire[938];							inform_L[981][8] = l_cell_wire[939];							inform_L[726][8] = l_cell_wire[940];							inform_L[982][8] = l_cell_wire[941];							inform_L[727][8] = l_cell_wire[942];							inform_L[983][8] = l_cell_wire[943];							inform_L[728][8] = l_cell_wire[944];							inform_L[984][8] = l_cell_wire[945];							inform_L[729][8] = l_cell_wire[946];							inform_L[985][8] = l_cell_wire[947];							inform_L[730][8] = l_cell_wire[948];							inform_L[986][8] = l_cell_wire[949];							inform_L[731][8] = l_cell_wire[950];							inform_L[987][8] = l_cell_wire[951];							inform_L[732][8] = l_cell_wire[952];							inform_L[988][8] = l_cell_wire[953];							inform_L[733][8] = l_cell_wire[954];							inform_L[989][8] = l_cell_wire[955];							inform_L[734][8] = l_cell_wire[956];							inform_L[990][8] = l_cell_wire[957];							inform_L[735][8] = l_cell_wire[958];							inform_L[991][8] = l_cell_wire[959];							inform_L[736][8] = l_cell_wire[960];							inform_L[992][8] = l_cell_wire[961];							inform_L[737][8] = l_cell_wire[962];							inform_L[993][8] = l_cell_wire[963];							inform_L[738][8] = l_cell_wire[964];							inform_L[994][8] = l_cell_wire[965];							inform_L[739][8] = l_cell_wire[966];							inform_L[995][8] = l_cell_wire[967];							inform_L[740][8] = l_cell_wire[968];							inform_L[996][8] = l_cell_wire[969];							inform_L[741][8] = l_cell_wire[970];							inform_L[997][8] = l_cell_wire[971];							inform_L[742][8] = l_cell_wire[972];							inform_L[998][8] = l_cell_wire[973];							inform_L[743][8] = l_cell_wire[974];							inform_L[999][8] = l_cell_wire[975];							inform_L[744][8] = l_cell_wire[976];							inform_L[1000][8] = l_cell_wire[977];							inform_L[745][8] = l_cell_wire[978];							inform_L[1001][8] = l_cell_wire[979];							inform_L[746][8] = l_cell_wire[980];							inform_L[1002][8] = l_cell_wire[981];							inform_L[747][8] = l_cell_wire[982];							inform_L[1003][8] = l_cell_wire[983];							inform_L[748][8] = l_cell_wire[984];							inform_L[1004][8] = l_cell_wire[985];							inform_L[749][8] = l_cell_wire[986];							inform_L[1005][8] = l_cell_wire[987];							inform_L[750][8] = l_cell_wire[988];							inform_L[1006][8] = l_cell_wire[989];							inform_L[751][8] = l_cell_wire[990];							inform_L[1007][8] = l_cell_wire[991];							inform_L[752][8] = l_cell_wire[992];							inform_L[1008][8] = l_cell_wire[993];							inform_L[753][8] = l_cell_wire[994];							inform_L[1009][8] = l_cell_wire[995];							inform_L[754][8] = l_cell_wire[996];							inform_L[1010][8] = l_cell_wire[997];							inform_L[755][8] = l_cell_wire[998];							inform_L[1011][8] = l_cell_wire[999];							inform_L[756][8] = l_cell_wire[1000];							inform_L[1012][8] = l_cell_wire[1001];							inform_L[757][8] = l_cell_wire[1002];							inform_L[1013][8] = l_cell_wire[1003];							inform_L[758][8] = l_cell_wire[1004];							inform_L[1014][8] = l_cell_wire[1005];							inform_L[759][8] = l_cell_wire[1006];							inform_L[1015][8] = l_cell_wire[1007];							inform_L[760][8] = l_cell_wire[1008];							inform_L[1016][8] = l_cell_wire[1009];							inform_L[761][8] = l_cell_wire[1010];							inform_L[1017][8] = l_cell_wire[1011];							inform_L[762][8] = l_cell_wire[1012];							inform_L[1018][8] = l_cell_wire[1013];							inform_L[763][8] = l_cell_wire[1014];							inform_L[1019][8] = l_cell_wire[1015];							inform_L[764][8] = l_cell_wire[1016];							inform_L[1020][8] = l_cell_wire[1017];							inform_L[765][8] = l_cell_wire[1018];							inform_L[1021][8] = l_cell_wire[1019];							inform_L[766][8] = l_cell_wire[1020];							inform_L[1022][8] = l_cell_wire[1021];							inform_L[767][8] = l_cell_wire[1022];							inform_L[1023][8] = l_cell_wire[1023];						end
						10:						begin							inform_R[0][10] = r_cell_wire[0];							inform_R[512][10] = r_cell_wire[1];							inform_R[1][10] = r_cell_wire[2];							inform_R[513][10] = r_cell_wire[3];							inform_R[2][10] = r_cell_wire[4];							inform_R[514][10] = r_cell_wire[5];							inform_R[3][10] = r_cell_wire[6];							inform_R[515][10] = r_cell_wire[7];							inform_R[4][10] = r_cell_wire[8];							inform_R[516][10] = r_cell_wire[9];							inform_R[5][10] = r_cell_wire[10];							inform_R[517][10] = r_cell_wire[11];							inform_R[6][10] = r_cell_wire[12];							inform_R[518][10] = r_cell_wire[13];							inform_R[7][10] = r_cell_wire[14];							inform_R[519][10] = r_cell_wire[15];							inform_R[8][10] = r_cell_wire[16];							inform_R[520][10] = r_cell_wire[17];							inform_R[9][10] = r_cell_wire[18];							inform_R[521][10] = r_cell_wire[19];							inform_R[10][10] = r_cell_wire[20];							inform_R[522][10] = r_cell_wire[21];							inform_R[11][10] = r_cell_wire[22];							inform_R[523][10] = r_cell_wire[23];							inform_R[12][10] = r_cell_wire[24];							inform_R[524][10] = r_cell_wire[25];							inform_R[13][10] = r_cell_wire[26];							inform_R[525][10] = r_cell_wire[27];							inform_R[14][10] = r_cell_wire[28];							inform_R[526][10] = r_cell_wire[29];							inform_R[15][10] = r_cell_wire[30];							inform_R[527][10] = r_cell_wire[31];							inform_R[16][10] = r_cell_wire[32];							inform_R[528][10] = r_cell_wire[33];							inform_R[17][10] = r_cell_wire[34];							inform_R[529][10] = r_cell_wire[35];							inform_R[18][10] = r_cell_wire[36];							inform_R[530][10] = r_cell_wire[37];							inform_R[19][10] = r_cell_wire[38];							inform_R[531][10] = r_cell_wire[39];							inform_R[20][10] = r_cell_wire[40];							inform_R[532][10] = r_cell_wire[41];							inform_R[21][10] = r_cell_wire[42];							inform_R[533][10] = r_cell_wire[43];							inform_R[22][10] = r_cell_wire[44];							inform_R[534][10] = r_cell_wire[45];							inform_R[23][10] = r_cell_wire[46];							inform_R[535][10] = r_cell_wire[47];							inform_R[24][10] = r_cell_wire[48];							inform_R[536][10] = r_cell_wire[49];							inform_R[25][10] = r_cell_wire[50];							inform_R[537][10] = r_cell_wire[51];							inform_R[26][10] = r_cell_wire[52];							inform_R[538][10] = r_cell_wire[53];							inform_R[27][10] = r_cell_wire[54];							inform_R[539][10] = r_cell_wire[55];							inform_R[28][10] = r_cell_wire[56];							inform_R[540][10] = r_cell_wire[57];							inform_R[29][10] = r_cell_wire[58];							inform_R[541][10] = r_cell_wire[59];							inform_R[30][10] = r_cell_wire[60];							inform_R[542][10] = r_cell_wire[61];							inform_R[31][10] = r_cell_wire[62];							inform_R[543][10] = r_cell_wire[63];							inform_R[32][10] = r_cell_wire[64];							inform_R[544][10] = r_cell_wire[65];							inform_R[33][10] = r_cell_wire[66];							inform_R[545][10] = r_cell_wire[67];							inform_R[34][10] = r_cell_wire[68];							inform_R[546][10] = r_cell_wire[69];							inform_R[35][10] = r_cell_wire[70];							inform_R[547][10] = r_cell_wire[71];							inform_R[36][10] = r_cell_wire[72];							inform_R[548][10] = r_cell_wire[73];							inform_R[37][10] = r_cell_wire[74];							inform_R[549][10] = r_cell_wire[75];							inform_R[38][10] = r_cell_wire[76];							inform_R[550][10] = r_cell_wire[77];							inform_R[39][10] = r_cell_wire[78];							inform_R[551][10] = r_cell_wire[79];							inform_R[40][10] = r_cell_wire[80];							inform_R[552][10] = r_cell_wire[81];							inform_R[41][10] = r_cell_wire[82];							inform_R[553][10] = r_cell_wire[83];							inform_R[42][10] = r_cell_wire[84];							inform_R[554][10] = r_cell_wire[85];							inform_R[43][10] = r_cell_wire[86];							inform_R[555][10] = r_cell_wire[87];							inform_R[44][10] = r_cell_wire[88];							inform_R[556][10] = r_cell_wire[89];							inform_R[45][10] = r_cell_wire[90];							inform_R[557][10] = r_cell_wire[91];							inform_R[46][10] = r_cell_wire[92];							inform_R[558][10] = r_cell_wire[93];							inform_R[47][10] = r_cell_wire[94];							inform_R[559][10] = r_cell_wire[95];							inform_R[48][10] = r_cell_wire[96];							inform_R[560][10] = r_cell_wire[97];							inform_R[49][10] = r_cell_wire[98];							inform_R[561][10] = r_cell_wire[99];							inform_R[50][10] = r_cell_wire[100];							inform_R[562][10] = r_cell_wire[101];							inform_R[51][10] = r_cell_wire[102];							inform_R[563][10] = r_cell_wire[103];							inform_R[52][10] = r_cell_wire[104];							inform_R[564][10] = r_cell_wire[105];							inform_R[53][10] = r_cell_wire[106];							inform_R[565][10] = r_cell_wire[107];							inform_R[54][10] = r_cell_wire[108];							inform_R[566][10] = r_cell_wire[109];							inform_R[55][10] = r_cell_wire[110];							inform_R[567][10] = r_cell_wire[111];							inform_R[56][10] = r_cell_wire[112];							inform_R[568][10] = r_cell_wire[113];							inform_R[57][10] = r_cell_wire[114];							inform_R[569][10] = r_cell_wire[115];							inform_R[58][10] = r_cell_wire[116];							inform_R[570][10] = r_cell_wire[117];							inform_R[59][10] = r_cell_wire[118];							inform_R[571][10] = r_cell_wire[119];							inform_R[60][10] = r_cell_wire[120];							inform_R[572][10] = r_cell_wire[121];							inform_R[61][10] = r_cell_wire[122];							inform_R[573][10] = r_cell_wire[123];							inform_R[62][10] = r_cell_wire[124];							inform_R[574][10] = r_cell_wire[125];							inform_R[63][10] = r_cell_wire[126];							inform_R[575][10] = r_cell_wire[127];							inform_R[64][10] = r_cell_wire[128];							inform_R[576][10] = r_cell_wire[129];							inform_R[65][10] = r_cell_wire[130];							inform_R[577][10] = r_cell_wire[131];							inform_R[66][10] = r_cell_wire[132];							inform_R[578][10] = r_cell_wire[133];							inform_R[67][10] = r_cell_wire[134];							inform_R[579][10] = r_cell_wire[135];							inform_R[68][10] = r_cell_wire[136];							inform_R[580][10] = r_cell_wire[137];							inform_R[69][10] = r_cell_wire[138];							inform_R[581][10] = r_cell_wire[139];							inform_R[70][10] = r_cell_wire[140];							inform_R[582][10] = r_cell_wire[141];							inform_R[71][10] = r_cell_wire[142];							inform_R[583][10] = r_cell_wire[143];							inform_R[72][10] = r_cell_wire[144];							inform_R[584][10] = r_cell_wire[145];							inform_R[73][10] = r_cell_wire[146];							inform_R[585][10] = r_cell_wire[147];							inform_R[74][10] = r_cell_wire[148];							inform_R[586][10] = r_cell_wire[149];							inform_R[75][10] = r_cell_wire[150];							inform_R[587][10] = r_cell_wire[151];							inform_R[76][10] = r_cell_wire[152];							inform_R[588][10] = r_cell_wire[153];							inform_R[77][10] = r_cell_wire[154];							inform_R[589][10] = r_cell_wire[155];							inform_R[78][10] = r_cell_wire[156];							inform_R[590][10] = r_cell_wire[157];							inform_R[79][10] = r_cell_wire[158];							inform_R[591][10] = r_cell_wire[159];							inform_R[80][10] = r_cell_wire[160];							inform_R[592][10] = r_cell_wire[161];							inform_R[81][10] = r_cell_wire[162];							inform_R[593][10] = r_cell_wire[163];							inform_R[82][10] = r_cell_wire[164];							inform_R[594][10] = r_cell_wire[165];							inform_R[83][10] = r_cell_wire[166];							inform_R[595][10] = r_cell_wire[167];							inform_R[84][10] = r_cell_wire[168];							inform_R[596][10] = r_cell_wire[169];							inform_R[85][10] = r_cell_wire[170];							inform_R[597][10] = r_cell_wire[171];							inform_R[86][10] = r_cell_wire[172];							inform_R[598][10] = r_cell_wire[173];							inform_R[87][10] = r_cell_wire[174];							inform_R[599][10] = r_cell_wire[175];							inform_R[88][10] = r_cell_wire[176];							inform_R[600][10] = r_cell_wire[177];							inform_R[89][10] = r_cell_wire[178];							inform_R[601][10] = r_cell_wire[179];							inform_R[90][10] = r_cell_wire[180];							inform_R[602][10] = r_cell_wire[181];							inform_R[91][10] = r_cell_wire[182];							inform_R[603][10] = r_cell_wire[183];							inform_R[92][10] = r_cell_wire[184];							inform_R[604][10] = r_cell_wire[185];							inform_R[93][10] = r_cell_wire[186];							inform_R[605][10] = r_cell_wire[187];							inform_R[94][10] = r_cell_wire[188];							inform_R[606][10] = r_cell_wire[189];							inform_R[95][10] = r_cell_wire[190];							inform_R[607][10] = r_cell_wire[191];							inform_R[96][10] = r_cell_wire[192];							inform_R[608][10] = r_cell_wire[193];							inform_R[97][10] = r_cell_wire[194];							inform_R[609][10] = r_cell_wire[195];							inform_R[98][10] = r_cell_wire[196];							inform_R[610][10] = r_cell_wire[197];							inform_R[99][10] = r_cell_wire[198];							inform_R[611][10] = r_cell_wire[199];							inform_R[100][10] = r_cell_wire[200];							inform_R[612][10] = r_cell_wire[201];							inform_R[101][10] = r_cell_wire[202];							inform_R[613][10] = r_cell_wire[203];							inform_R[102][10] = r_cell_wire[204];							inform_R[614][10] = r_cell_wire[205];							inform_R[103][10] = r_cell_wire[206];							inform_R[615][10] = r_cell_wire[207];							inform_R[104][10] = r_cell_wire[208];							inform_R[616][10] = r_cell_wire[209];							inform_R[105][10] = r_cell_wire[210];							inform_R[617][10] = r_cell_wire[211];							inform_R[106][10] = r_cell_wire[212];							inform_R[618][10] = r_cell_wire[213];							inform_R[107][10] = r_cell_wire[214];							inform_R[619][10] = r_cell_wire[215];							inform_R[108][10] = r_cell_wire[216];							inform_R[620][10] = r_cell_wire[217];							inform_R[109][10] = r_cell_wire[218];							inform_R[621][10] = r_cell_wire[219];							inform_R[110][10] = r_cell_wire[220];							inform_R[622][10] = r_cell_wire[221];							inform_R[111][10] = r_cell_wire[222];							inform_R[623][10] = r_cell_wire[223];							inform_R[112][10] = r_cell_wire[224];							inform_R[624][10] = r_cell_wire[225];							inform_R[113][10] = r_cell_wire[226];							inform_R[625][10] = r_cell_wire[227];							inform_R[114][10] = r_cell_wire[228];							inform_R[626][10] = r_cell_wire[229];							inform_R[115][10] = r_cell_wire[230];							inform_R[627][10] = r_cell_wire[231];							inform_R[116][10] = r_cell_wire[232];							inform_R[628][10] = r_cell_wire[233];							inform_R[117][10] = r_cell_wire[234];							inform_R[629][10] = r_cell_wire[235];							inform_R[118][10] = r_cell_wire[236];							inform_R[630][10] = r_cell_wire[237];							inform_R[119][10] = r_cell_wire[238];							inform_R[631][10] = r_cell_wire[239];							inform_R[120][10] = r_cell_wire[240];							inform_R[632][10] = r_cell_wire[241];							inform_R[121][10] = r_cell_wire[242];							inform_R[633][10] = r_cell_wire[243];							inform_R[122][10] = r_cell_wire[244];							inform_R[634][10] = r_cell_wire[245];							inform_R[123][10] = r_cell_wire[246];							inform_R[635][10] = r_cell_wire[247];							inform_R[124][10] = r_cell_wire[248];							inform_R[636][10] = r_cell_wire[249];							inform_R[125][10] = r_cell_wire[250];							inform_R[637][10] = r_cell_wire[251];							inform_R[126][10] = r_cell_wire[252];							inform_R[638][10] = r_cell_wire[253];							inform_R[127][10] = r_cell_wire[254];							inform_R[639][10] = r_cell_wire[255];							inform_R[128][10] = r_cell_wire[256];							inform_R[640][10] = r_cell_wire[257];							inform_R[129][10] = r_cell_wire[258];							inform_R[641][10] = r_cell_wire[259];							inform_R[130][10] = r_cell_wire[260];							inform_R[642][10] = r_cell_wire[261];							inform_R[131][10] = r_cell_wire[262];							inform_R[643][10] = r_cell_wire[263];							inform_R[132][10] = r_cell_wire[264];							inform_R[644][10] = r_cell_wire[265];							inform_R[133][10] = r_cell_wire[266];							inform_R[645][10] = r_cell_wire[267];							inform_R[134][10] = r_cell_wire[268];							inform_R[646][10] = r_cell_wire[269];							inform_R[135][10] = r_cell_wire[270];							inform_R[647][10] = r_cell_wire[271];							inform_R[136][10] = r_cell_wire[272];							inform_R[648][10] = r_cell_wire[273];							inform_R[137][10] = r_cell_wire[274];							inform_R[649][10] = r_cell_wire[275];							inform_R[138][10] = r_cell_wire[276];							inform_R[650][10] = r_cell_wire[277];							inform_R[139][10] = r_cell_wire[278];							inform_R[651][10] = r_cell_wire[279];							inform_R[140][10] = r_cell_wire[280];							inform_R[652][10] = r_cell_wire[281];							inform_R[141][10] = r_cell_wire[282];							inform_R[653][10] = r_cell_wire[283];							inform_R[142][10] = r_cell_wire[284];							inform_R[654][10] = r_cell_wire[285];							inform_R[143][10] = r_cell_wire[286];							inform_R[655][10] = r_cell_wire[287];							inform_R[144][10] = r_cell_wire[288];							inform_R[656][10] = r_cell_wire[289];							inform_R[145][10] = r_cell_wire[290];							inform_R[657][10] = r_cell_wire[291];							inform_R[146][10] = r_cell_wire[292];							inform_R[658][10] = r_cell_wire[293];							inform_R[147][10] = r_cell_wire[294];							inform_R[659][10] = r_cell_wire[295];							inform_R[148][10] = r_cell_wire[296];							inform_R[660][10] = r_cell_wire[297];							inform_R[149][10] = r_cell_wire[298];							inform_R[661][10] = r_cell_wire[299];							inform_R[150][10] = r_cell_wire[300];							inform_R[662][10] = r_cell_wire[301];							inform_R[151][10] = r_cell_wire[302];							inform_R[663][10] = r_cell_wire[303];							inform_R[152][10] = r_cell_wire[304];							inform_R[664][10] = r_cell_wire[305];							inform_R[153][10] = r_cell_wire[306];							inform_R[665][10] = r_cell_wire[307];							inform_R[154][10] = r_cell_wire[308];							inform_R[666][10] = r_cell_wire[309];							inform_R[155][10] = r_cell_wire[310];							inform_R[667][10] = r_cell_wire[311];							inform_R[156][10] = r_cell_wire[312];							inform_R[668][10] = r_cell_wire[313];							inform_R[157][10] = r_cell_wire[314];							inform_R[669][10] = r_cell_wire[315];							inform_R[158][10] = r_cell_wire[316];							inform_R[670][10] = r_cell_wire[317];							inform_R[159][10] = r_cell_wire[318];							inform_R[671][10] = r_cell_wire[319];							inform_R[160][10] = r_cell_wire[320];							inform_R[672][10] = r_cell_wire[321];							inform_R[161][10] = r_cell_wire[322];							inform_R[673][10] = r_cell_wire[323];							inform_R[162][10] = r_cell_wire[324];							inform_R[674][10] = r_cell_wire[325];							inform_R[163][10] = r_cell_wire[326];							inform_R[675][10] = r_cell_wire[327];							inform_R[164][10] = r_cell_wire[328];							inform_R[676][10] = r_cell_wire[329];							inform_R[165][10] = r_cell_wire[330];							inform_R[677][10] = r_cell_wire[331];							inform_R[166][10] = r_cell_wire[332];							inform_R[678][10] = r_cell_wire[333];							inform_R[167][10] = r_cell_wire[334];							inform_R[679][10] = r_cell_wire[335];							inform_R[168][10] = r_cell_wire[336];							inform_R[680][10] = r_cell_wire[337];							inform_R[169][10] = r_cell_wire[338];							inform_R[681][10] = r_cell_wire[339];							inform_R[170][10] = r_cell_wire[340];							inform_R[682][10] = r_cell_wire[341];							inform_R[171][10] = r_cell_wire[342];							inform_R[683][10] = r_cell_wire[343];							inform_R[172][10] = r_cell_wire[344];							inform_R[684][10] = r_cell_wire[345];							inform_R[173][10] = r_cell_wire[346];							inform_R[685][10] = r_cell_wire[347];							inform_R[174][10] = r_cell_wire[348];							inform_R[686][10] = r_cell_wire[349];							inform_R[175][10] = r_cell_wire[350];							inform_R[687][10] = r_cell_wire[351];							inform_R[176][10] = r_cell_wire[352];							inform_R[688][10] = r_cell_wire[353];							inform_R[177][10] = r_cell_wire[354];							inform_R[689][10] = r_cell_wire[355];							inform_R[178][10] = r_cell_wire[356];							inform_R[690][10] = r_cell_wire[357];							inform_R[179][10] = r_cell_wire[358];							inform_R[691][10] = r_cell_wire[359];							inform_R[180][10] = r_cell_wire[360];							inform_R[692][10] = r_cell_wire[361];							inform_R[181][10] = r_cell_wire[362];							inform_R[693][10] = r_cell_wire[363];							inform_R[182][10] = r_cell_wire[364];							inform_R[694][10] = r_cell_wire[365];							inform_R[183][10] = r_cell_wire[366];							inform_R[695][10] = r_cell_wire[367];							inform_R[184][10] = r_cell_wire[368];							inform_R[696][10] = r_cell_wire[369];							inform_R[185][10] = r_cell_wire[370];							inform_R[697][10] = r_cell_wire[371];							inform_R[186][10] = r_cell_wire[372];							inform_R[698][10] = r_cell_wire[373];							inform_R[187][10] = r_cell_wire[374];							inform_R[699][10] = r_cell_wire[375];							inform_R[188][10] = r_cell_wire[376];							inform_R[700][10] = r_cell_wire[377];							inform_R[189][10] = r_cell_wire[378];							inform_R[701][10] = r_cell_wire[379];							inform_R[190][10] = r_cell_wire[380];							inform_R[702][10] = r_cell_wire[381];							inform_R[191][10] = r_cell_wire[382];							inform_R[703][10] = r_cell_wire[383];							inform_R[192][10] = r_cell_wire[384];							inform_R[704][10] = r_cell_wire[385];							inform_R[193][10] = r_cell_wire[386];							inform_R[705][10] = r_cell_wire[387];							inform_R[194][10] = r_cell_wire[388];							inform_R[706][10] = r_cell_wire[389];							inform_R[195][10] = r_cell_wire[390];							inform_R[707][10] = r_cell_wire[391];							inform_R[196][10] = r_cell_wire[392];							inform_R[708][10] = r_cell_wire[393];							inform_R[197][10] = r_cell_wire[394];							inform_R[709][10] = r_cell_wire[395];							inform_R[198][10] = r_cell_wire[396];							inform_R[710][10] = r_cell_wire[397];							inform_R[199][10] = r_cell_wire[398];							inform_R[711][10] = r_cell_wire[399];							inform_R[200][10] = r_cell_wire[400];							inform_R[712][10] = r_cell_wire[401];							inform_R[201][10] = r_cell_wire[402];							inform_R[713][10] = r_cell_wire[403];							inform_R[202][10] = r_cell_wire[404];							inform_R[714][10] = r_cell_wire[405];							inform_R[203][10] = r_cell_wire[406];							inform_R[715][10] = r_cell_wire[407];							inform_R[204][10] = r_cell_wire[408];							inform_R[716][10] = r_cell_wire[409];							inform_R[205][10] = r_cell_wire[410];							inform_R[717][10] = r_cell_wire[411];							inform_R[206][10] = r_cell_wire[412];							inform_R[718][10] = r_cell_wire[413];							inform_R[207][10] = r_cell_wire[414];							inform_R[719][10] = r_cell_wire[415];							inform_R[208][10] = r_cell_wire[416];							inform_R[720][10] = r_cell_wire[417];							inform_R[209][10] = r_cell_wire[418];							inform_R[721][10] = r_cell_wire[419];							inform_R[210][10] = r_cell_wire[420];							inform_R[722][10] = r_cell_wire[421];							inform_R[211][10] = r_cell_wire[422];							inform_R[723][10] = r_cell_wire[423];							inform_R[212][10] = r_cell_wire[424];							inform_R[724][10] = r_cell_wire[425];							inform_R[213][10] = r_cell_wire[426];							inform_R[725][10] = r_cell_wire[427];							inform_R[214][10] = r_cell_wire[428];							inform_R[726][10] = r_cell_wire[429];							inform_R[215][10] = r_cell_wire[430];							inform_R[727][10] = r_cell_wire[431];							inform_R[216][10] = r_cell_wire[432];							inform_R[728][10] = r_cell_wire[433];							inform_R[217][10] = r_cell_wire[434];							inform_R[729][10] = r_cell_wire[435];							inform_R[218][10] = r_cell_wire[436];							inform_R[730][10] = r_cell_wire[437];							inform_R[219][10] = r_cell_wire[438];							inform_R[731][10] = r_cell_wire[439];							inform_R[220][10] = r_cell_wire[440];							inform_R[732][10] = r_cell_wire[441];							inform_R[221][10] = r_cell_wire[442];							inform_R[733][10] = r_cell_wire[443];							inform_R[222][10] = r_cell_wire[444];							inform_R[734][10] = r_cell_wire[445];							inform_R[223][10] = r_cell_wire[446];							inform_R[735][10] = r_cell_wire[447];							inform_R[224][10] = r_cell_wire[448];							inform_R[736][10] = r_cell_wire[449];							inform_R[225][10] = r_cell_wire[450];							inform_R[737][10] = r_cell_wire[451];							inform_R[226][10] = r_cell_wire[452];							inform_R[738][10] = r_cell_wire[453];							inform_R[227][10] = r_cell_wire[454];							inform_R[739][10] = r_cell_wire[455];							inform_R[228][10] = r_cell_wire[456];							inform_R[740][10] = r_cell_wire[457];							inform_R[229][10] = r_cell_wire[458];							inform_R[741][10] = r_cell_wire[459];							inform_R[230][10] = r_cell_wire[460];							inform_R[742][10] = r_cell_wire[461];							inform_R[231][10] = r_cell_wire[462];							inform_R[743][10] = r_cell_wire[463];							inform_R[232][10] = r_cell_wire[464];							inform_R[744][10] = r_cell_wire[465];							inform_R[233][10] = r_cell_wire[466];							inform_R[745][10] = r_cell_wire[467];							inform_R[234][10] = r_cell_wire[468];							inform_R[746][10] = r_cell_wire[469];							inform_R[235][10] = r_cell_wire[470];							inform_R[747][10] = r_cell_wire[471];							inform_R[236][10] = r_cell_wire[472];							inform_R[748][10] = r_cell_wire[473];							inform_R[237][10] = r_cell_wire[474];							inform_R[749][10] = r_cell_wire[475];							inform_R[238][10] = r_cell_wire[476];							inform_R[750][10] = r_cell_wire[477];							inform_R[239][10] = r_cell_wire[478];							inform_R[751][10] = r_cell_wire[479];							inform_R[240][10] = r_cell_wire[480];							inform_R[752][10] = r_cell_wire[481];							inform_R[241][10] = r_cell_wire[482];							inform_R[753][10] = r_cell_wire[483];							inform_R[242][10] = r_cell_wire[484];							inform_R[754][10] = r_cell_wire[485];							inform_R[243][10] = r_cell_wire[486];							inform_R[755][10] = r_cell_wire[487];							inform_R[244][10] = r_cell_wire[488];							inform_R[756][10] = r_cell_wire[489];							inform_R[245][10] = r_cell_wire[490];							inform_R[757][10] = r_cell_wire[491];							inform_R[246][10] = r_cell_wire[492];							inform_R[758][10] = r_cell_wire[493];							inform_R[247][10] = r_cell_wire[494];							inform_R[759][10] = r_cell_wire[495];							inform_R[248][10] = r_cell_wire[496];							inform_R[760][10] = r_cell_wire[497];							inform_R[249][10] = r_cell_wire[498];							inform_R[761][10] = r_cell_wire[499];							inform_R[250][10] = r_cell_wire[500];							inform_R[762][10] = r_cell_wire[501];							inform_R[251][10] = r_cell_wire[502];							inform_R[763][10] = r_cell_wire[503];							inform_R[252][10] = r_cell_wire[504];							inform_R[764][10] = r_cell_wire[505];							inform_R[253][10] = r_cell_wire[506];							inform_R[765][10] = r_cell_wire[507];							inform_R[254][10] = r_cell_wire[508];							inform_R[766][10] = r_cell_wire[509];							inform_R[255][10] = r_cell_wire[510];							inform_R[767][10] = r_cell_wire[511];							inform_R[256][10] = r_cell_wire[512];							inform_R[768][10] = r_cell_wire[513];							inform_R[257][10] = r_cell_wire[514];							inform_R[769][10] = r_cell_wire[515];							inform_R[258][10] = r_cell_wire[516];							inform_R[770][10] = r_cell_wire[517];							inform_R[259][10] = r_cell_wire[518];							inform_R[771][10] = r_cell_wire[519];							inform_R[260][10] = r_cell_wire[520];							inform_R[772][10] = r_cell_wire[521];							inform_R[261][10] = r_cell_wire[522];							inform_R[773][10] = r_cell_wire[523];							inform_R[262][10] = r_cell_wire[524];							inform_R[774][10] = r_cell_wire[525];							inform_R[263][10] = r_cell_wire[526];							inform_R[775][10] = r_cell_wire[527];							inform_R[264][10] = r_cell_wire[528];							inform_R[776][10] = r_cell_wire[529];							inform_R[265][10] = r_cell_wire[530];							inform_R[777][10] = r_cell_wire[531];							inform_R[266][10] = r_cell_wire[532];							inform_R[778][10] = r_cell_wire[533];							inform_R[267][10] = r_cell_wire[534];							inform_R[779][10] = r_cell_wire[535];							inform_R[268][10] = r_cell_wire[536];							inform_R[780][10] = r_cell_wire[537];							inform_R[269][10] = r_cell_wire[538];							inform_R[781][10] = r_cell_wire[539];							inform_R[270][10] = r_cell_wire[540];							inform_R[782][10] = r_cell_wire[541];							inform_R[271][10] = r_cell_wire[542];							inform_R[783][10] = r_cell_wire[543];							inform_R[272][10] = r_cell_wire[544];							inform_R[784][10] = r_cell_wire[545];							inform_R[273][10] = r_cell_wire[546];							inform_R[785][10] = r_cell_wire[547];							inform_R[274][10] = r_cell_wire[548];							inform_R[786][10] = r_cell_wire[549];							inform_R[275][10] = r_cell_wire[550];							inform_R[787][10] = r_cell_wire[551];							inform_R[276][10] = r_cell_wire[552];							inform_R[788][10] = r_cell_wire[553];							inform_R[277][10] = r_cell_wire[554];							inform_R[789][10] = r_cell_wire[555];							inform_R[278][10] = r_cell_wire[556];							inform_R[790][10] = r_cell_wire[557];							inform_R[279][10] = r_cell_wire[558];							inform_R[791][10] = r_cell_wire[559];							inform_R[280][10] = r_cell_wire[560];							inform_R[792][10] = r_cell_wire[561];							inform_R[281][10] = r_cell_wire[562];							inform_R[793][10] = r_cell_wire[563];							inform_R[282][10] = r_cell_wire[564];							inform_R[794][10] = r_cell_wire[565];							inform_R[283][10] = r_cell_wire[566];							inform_R[795][10] = r_cell_wire[567];							inform_R[284][10] = r_cell_wire[568];							inform_R[796][10] = r_cell_wire[569];							inform_R[285][10] = r_cell_wire[570];							inform_R[797][10] = r_cell_wire[571];							inform_R[286][10] = r_cell_wire[572];							inform_R[798][10] = r_cell_wire[573];							inform_R[287][10] = r_cell_wire[574];							inform_R[799][10] = r_cell_wire[575];							inform_R[288][10] = r_cell_wire[576];							inform_R[800][10] = r_cell_wire[577];							inform_R[289][10] = r_cell_wire[578];							inform_R[801][10] = r_cell_wire[579];							inform_R[290][10] = r_cell_wire[580];							inform_R[802][10] = r_cell_wire[581];							inform_R[291][10] = r_cell_wire[582];							inform_R[803][10] = r_cell_wire[583];							inform_R[292][10] = r_cell_wire[584];							inform_R[804][10] = r_cell_wire[585];							inform_R[293][10] = r_cell_wire[586];							inform_R[805][10] = r_cell_wire[587];							inform_R[294][10] = r_cell_wire[588];							inform_R[806][10] = r_cell_wire[589];							inform_R[295][10] = r_cell_wire[590];							inform_R[807][10] = r_cell_wire[591];							inform_R[296][10] = r_cell_wire[592];							inform_R[808][10] = r_cell_wire[593];							inform_R[297][10] = r_cell_wire[594];							inform_R[809][10] = r_cell_wire[595];							inform_R[298][10] = r_cell_wire[596];							inform_R[810][10] = r_cell_wire[597];							inform_R[299][10] = r_cell_wire[598];							inform_R[811][10] = r_cell_wire[599];							inform_R[300][10] = r_cell_wire[600];							inform_R[812][10] = r_cell_wire[601];							inform_R[301][10] = r_cell_wire[602];							inform_R[813][10] = r_cell_wire[603];							inform_R[302][10] = r_cell_wire[604];							inform_R[814][10] = r_cell_wire[605];							inform_R[303][10] = r_cell_wire[606];							inform_R[815][10] = r_cell_wire[607];							inform_R[304][10] = r_cell_wire[608];							inform_R[816][10] = r_cell_wire[609];							inform_R[305][10] = r_cell_wire[610];							inform_R[817][10] = r_cell_wire[611];							inform_R[306][10] = r_cell_wire[612];							inform_R[818][10] = r_cell_wire[613];							inform_R[307][10] = r_cell_wire[614];							inform_R[819][10] = r_cell_wire[615];							inform_R[308][10] = r_cell_wire[616];							inform_R[820][10] = r_cell_wire[617];							inform_R[309][10] = r_cell_wire[618];							inform_R[821][10] = r_cell_wire[619];							inform_R[310][10] = r_cell_wire[620];							inform_R[822][10] = r_cell_wire[621];							inform_R[311][10] = r_cell_wire[622];							inform_R[823][10] = r_cell_wire[623];							inform_R[312][10] = r_cell_wire[624];							inform_R[824][10] = r_cell_wire[625];							inform_R[313][10] = r_cell_wire[626];							inform_R[825][10] = r_cell_wire[627];							inform_R[314][10] = r_cell_wire[628];							inform_R[826][10] = r_cell_wire[629];							inform_R[315][10] = r_cell_wire[630];							inform_R[827][10] = r_cell_wire[631];							inform_R[316][10] = r_cell_wire[632];							inform_R[828][10] = r_cell_wire[633];							inform_R[317][10] = r_cell_wire[634];							inform_R[829][10] = r_cell_wire[635];							inform_R[318][10] = r_cell_wire[636];							inform_R[830][10] = r_cell_wire[637];							inform_R[319][10] = r_cell_wire[638];							inform_R[831][10] = r_cell_wire[639];							inform_R[320][10] = r_cell_wire[640];							inform_R[832][10] = r_cell_wire[641];							inform_R[321][10] = r_cell_wire[642];							inform_R[833][10] = r_cell_wire[643];							inform_R[322][10] = r_cell_wire[644];							inform_R[834][10] = r_cell_wire[645];							inform_R[323][10] = r_cell_wire[646];							inform_R[835][10] = r_cell_wire[647];							inform_R[324][10] = r_cell_wire[648];							inform_R[836][10] = r_cell_wire[649];							inform_R[325][10] = r_cell_wire[650];							inform_R[837][10] = r_cell_wire[651];							inform_R[326][10] = r_cell_wire[652];							inform_R[838][10] = r_cell_wire[653];							inform_R[327][10] = r_cell_wire[654];							inform_R[839][10] = r_cell_wire[655];							inform_R[328][10] = r_cell_wire[656];							inform_R[840][10] = r_cell_wire[657];							inform_R[329][10] = r_cell_wire[658];							inform_R[841][10] = r_cell_wire[659];							inform_R[330][10] = r_cell_wire[660];							inform_R[842][10] = r_cell_wire[661];							inform_R[331][10] = r_cell_wire[662];							inform_R[843][10] = r_cell_wire[663];							inform_R[332][10] = r_cell_wire[664];							inform_R[844][10] = r_cell_wire[665];							inform_R[333][10] = r_cell_wire[666];							inform_R[845][10] = r_cell_wire[667];							inform_R[334][10] = r_cell_wire[668];							inform_R[846][10] = r_cell_wire[669];							inform_R[335][10] = r_cell_wire[670];							inform_R[847][10] = r_cell_wire[671];							inform_R[336][10] = r_cell_wire[672];							inform_R[848][10] = r_cell_wire[673];							inform_R[337][10] = r_cell_wire[674];							inform_R[849][10] = r_cell_wire[675];							inform_R[338][10] = r_cell_wire[676];							inform_R[850][10] = r_cell_wire[677];							inform_R[339][10] = r_cell_wire[678];							inform_R[851][10] = r_cell_wire[679];							inform_R[340][10] = r_cell_wire[680];							inform_R[852][10] = r_cell_wire[681];							inform_R[341][10] = r_cell_wire[682];							inform_R[853][10] = r_cell_wire[683];							inform_R[342][10] = r_cell_wire[684];							inform_R[854][10] = r_cell_wire[685];							inform_R[343][10] = r_cell_wire[686];							inform_R[855][10] = r_cell_wire[687];							inform_R[344][10] = r_cell_wire[688];							inform_R[856][10] = r_cell_wire[689];							inform_R[345][10] = r_cell_wire[690];							inform_R[857][10] = r_cell_wire[691];							inform_R[346][10] = r_cell_wire[692];							inform_R[858][10] = r_cell_wire[693];							inform_R[347][10] = r_cell_wire[694];							inform_R[859][10] = r_cell_wire[695];							inform_R[348][10] = r_cell_wire[696];							inform_R[860][10] = r_cell_wire[697];							inform_R[349][10] = r_cell_wire[698];							inform_R[861][10] = r_cell_wire[699];							inform_R[350][10] = r_cell_wire[700];							inform_R[862][10] = r_cell_wire[701];							inform_R[351][10] = r_cell_wire[702];							inform_R[863][10] = r_cell_wire[703];							inform_R[352][10] = r_cell_wire[704];							inform_R[864][10] = r_cell_wire[705];							inform_R[353][10] = r_cell_wire[706];							inform_R[865][10] = r_cell_wire[707];							inform_R[354][10] = r_cell_wire[708];							inform_R[866][10] = r_cell_wire[709];							inform_R[355][10] = r_cell_wire[710];							inform_R[867][10] = r_cell_wire[711];							inform_R[356][10] = r_cell_wire[712];							inform_R[868][10] = r_cell_wire[713];							inform_R[357][10] = r_cell_wire[714];							inform_R[869][10] = r_cell_wire[715];							inform_R[358][10] = r_cell_wire[716];							inform_R[870][10] = r_cell_wire[717];							inform_R[359][10] = r_cell_wire[718];							inform_R[871][10] = r_cell_wire[719];							inform_R[360][10] = r_cell_wire[720];							inform_R[872][10] = r_cell_wire[721];							inform_R[361][10] = r_cell_wire[722];							inform_R[873][10] = r_cell_wire[723];							inform_R[362][10] = r_cell_wire[724];							inform_R[874][10] = r_cell_wire[725];							inform_R[363][10] = r_cell_wire[726];							inform_R[875][10] = r_cell_wire[727];							inform_R[364][10] = r_cell_wire[728];							inform_R[876][10] = r_cell_wire[729];							inform_R[365][10] = r_cell_wire[730];							inform_R[877][10] = r_cell_wire[731];							inform_R[366][10] = r_cell_wire[732];							inform_R[878][10] = r_cell_wire[733];							inform_R[367][10] = r_cell_wire[734];							inform_R[879][10] = r_cell_wire[735];							inform_R[368][10] = r_cell_wire[736];							inform_R[880][10] = r_cell_wire[737];							inform_R[369][10] = r_cell_wire[738];							inform_R[881][10] = r_cell_wire[739];							inform_R[370][10] = r_cell_wire[740];							inform_R[882][10] = r_cell_wire[741];							inform_R[371][10] = r_cell_wire[742];							inform_R[883][10] = r_cell_wire[743];							inform_R[372][10] = r_cell_wire[744];							inform_R[884][10] = r_cell_wire[745];							inform_R[373][10] = r_cell_wire[746];							inform_R[885][10] = r_cell_wire[747];							inform_R[374][10] = r_cell_wire[748];							inform_R[886][10] = r_cell_wire[749];							inform_R[375][10] = r_cell_wire[750];							inform_R[887][10] = r_cell_wire[751];							inform_R[376][10] = r_cell_wire[752];							inform_R[888][10] = r_cell_wire[753];							inform_R[377][10] = r_cell_wire[754];							inform_R[889][10] = r_cell_wire[755];							inform_R[378][10] = r_cell_wire[756];							inform_R[890][10] = r_cell_wire[757];							inform_R[379][10] = r_cell_wire[758];							inform_R[891][10] = r_cell_wire[759];							inform_R[380][10] = r_cell_wire[760];							inform_R[892][10] = r_cell_wire[761];							inform_R[381][10] = r_cell_wire[762];							inform_R[893][10] = r_cell_wire[763];							inform_R[382][10] = r_cell_wire[764];							inform_R[894][10] = r_cell_wire[765];							inform_R[383][10] = r_cell_wire[766];							inform_R[895][10] = r_cell_wire[767];							inform_R[384][10] = r_cell_wire[768];							inform_R[896][10] = r_cell_wire[769];							inform_R[385][10] = r_cell_wire[770];							inform_R[897][10] = r_cell_wire[771];							inform_R[386][10] = r_cell_wire[772];							inform_R[898][10] = r_cell_wire[773];							inform_R[387][10] = r_cell_wire[774];							inform_R[899][10] = r_cell_wire[775];							inform_R[388][10] = r_cell_wire[776];							inform_R[900][10] = r_cell_wire[777];							inform_R[389][10] = r_cell_wire[778];							inform_R[901][10] = r_cell_wire[779];							inform_R[390][10] = r_cell_wire[780];							inform_R[902][10] = r_cell_wire[781];							inform_R[391][10] = r_cell_wire[782];							inform_R[903][10] = r_cell_wire[783];							inform_R[392][10] = r_cell_wire[784];							inform_R[904][10] = r_cell_wire[785];							inform_R[393][10] = r_cell_wire[786];							inform_R[905][10] = r_cell_wire[787];							inform_R[394][10] = r_cell_wire[788];							inform_R[906][10] = r_cell_wire[789];							inform_R[395][10] = r_cell_wire[790];							inform_R[907][10] = r_cell_wire[791];							inform_R[396][10] = r_cell_wire[792];							inform_R[908][10] = r_cell_wire[793];							inform_R[397][10] = r_cell_wire[794];							inform_R[909][10] = r_cell_wire[795];							inform_R[398][10] = r_cell_wire[796];							inform_R[910][10] = r_cell_wire[797];							inform_R[399][10] = r_cell_wire[798];							inform_R[911][10] = r_cell_wire[799];							inform_R[400][10] = r_cell_wire[800];							inform_R[912][10] = r_cell_wire[801];							inform_R[401][10] = r_cell_wire[802];							inform_R[913][10] = r_cell_wire[803];							inform_R[402][10] = r_cell_wire[804];							inform_R[914][10] = r_cell_wire[805];							inform_R[403][10] = r_cell_wire[806];							inform_R[915][10] = r_cell_wire[807];							inform_R[404][10] = r_cell_wire[808];							inform_R[916][10] = r_cell_wire[809];							inform_R[405][10] = r_cell_wire[810];							inform_R[917][10] = r_cell_wire[811];							inform_R[406][10] = r_cell_wire[812];							inform_R[918][10] = r_cell_wire[813];							inform_R[407][10] = r_cell_wire[814];							inform_R[919][10] = r_cell_wire[815];							inform_R[408][10] = r_cell_wire[816];							inform_R[920][10] = r_cell_wire[817];							inform_R[409][10] = r_cell_wire[818];							inform_R[921][10] = r_cell_wire[819];							inform_R[410][10] = r_cell_wire[820];							inform_R[922][10] = r_cell_wire[821];							inform_R[411][10] = r_cell_wire[822];							inform_R[923][10] = r_cell_wire[823];							inform_R[412][10] = r_cell_wire[824];							inform_R[924][10] = r_cell_wire[825];							inform_R[413][10] = r_cell_wire[826];							inform_R[925][10] = r_cell_wire[827];							inform_R[414][10] = r_cell_wire[828];							inform_R[926][10] = r_cell_wire[829];							inform_R[415][10] = r_cell_wire[830];							inform_R[927][10] = r_cell_wire[831];							inform_R[416][10] = r_cell_wire[832];							inform_R[928][10] = r_cell_wire[833];							inform_R[417][10] = r_cell_wire[834];							inform_R[929][10] = r_cell_wire[835];							inform_R[418][10] = r_cell_wire[836];							inform_R[930][10] = r_cell_wire[837];							inform_R[419][10] = r_cell_wire[838];							inform_R[931][10] = r_cell_wire[839];							inform_R[420][10] = r_cell_wire[840];							inform_R[932][10] = r_cell_wire[841];							inform_R[421][10] = r_cell_wire[842];							inform_R[933][10] = r_cell_wire[843];							inform_R[422][10] = r_cell_wire[844];							inform_R[934][10] = r_cell_wire[845];							inform_R[423][10] = r_cell_wire[846];							inform_R[935][10] = r_cell_wire[847];							inform_R[424][10] = r_cell_wire[848];							inform_R[936][10] = r_cell_wire[849];							inform_R[425][10] = r_cell_wire[850];							inform_R[937][10] = r_cell_wire[851];							inform_R[426][10] = r_cell_wire[852];							inform_R[938][10] = r_cell_wire[853];							inform_R[427][10] = r_cell_wire[854];							inform_R[939][10] = r_cell_wire[855];							inform_R[428][10] = r_cell_wire[856];							inform_R[940][10] = r_cell_wire[857];							inform_R[429][10] = r_cell_wire[858];							inform_R[941][10] = r_cell_wire[859];							inform_R[430][10] = r_cell_wire[860];							inform_R[942][10] = r_cell_wire[861];							inform_R[431][10] = r_cell_wire[862];							inform_R[943][10] = r_cell_wire[863];							inform_R[432][10] = r_cell_wire[864];							inform_R[944][10] = r_cell_wire[865];							inform_R[433][10] = r_cell_wire[866];							inform_R[945][10] = r_cell_wire[867];							inform_R[434][10] = r_cell_wire[868];							inform_R[946][10] = r_cell_wire[869];							inform_R[435][10] = r_cell_wire[870];							inform_R[947][10] = r_cell_wire[871];							inform_R[436][10] = r_cell_wire[872];							inform_R[948][10] = r_cell_wire[873];							inform_R[437][10] = r_cell_wire[874];							inform_R[949][10] = r_cell_wire[875];							inform_R[438][10] = r_cell_wire[876];							inform_R[950][10] = r_cell_wire[877];							inform_R[439][10] = r_cell_wire[878];							inform_R[951][10] = r_cell_wire[879];							inform_R[440][10] = r_cell_wire[880];							inform_R[952][10] = r_cell_wire[881];							inform_R[441][10] = r_cell_wire[882];							inform_R[953][10] = r_cell_wire[883];							inform_R[442][10] = r_cell_wire[884];							inform_R[954][10] = r_cell_wire[885];							inform_R[443][10] = r_cell_wire[886];							inform_R[955][10] = r_cell_wire[887];							inform_R[444][10] = r_cell_wire[888];							inform_R[956][10] = r_cell_wire[889];							inform_R[445][10] = r_cell_wire[890];							inform_R[957][10] = r_cell_wire[891];							inform_R[446][10] = r_cell_wire[892];							inform_R[958][10] = r_cell_wire[893];							inform_R[447][10] = r_cell_wire[894];							inform_R[959][10] = r_cell_wire[895];							inform_R[448][10] = r_cell_wire[896];							inform_R[960][10] = r_cell_wire[897];							inform_R[449][10] = r_cell_wire[898];							inform_R[961][10] = r_cell_wire[899];							inform_R[450][10] = r_cell_wire[900];							inform_R[962][10] = r_cell_wire[901];							inform_R[451][10] = r_cell_wire[902];							inform_R[963][10] = r_cell_wire[903];							inform_R[452][10] = r_cell_wire[904];							inform_R[964][10] = r_cell_wire[905];							inform_R[453][10] = r_cell_wire[906];							inform_R[965][10] = r_cell_wire[907];							inform_R[454][10] = r_cell_wire[908];							inform_R[966][10] = r_cell_wire[909];							inform_R[455][10] = r_cell_wire[910];							inform_R[967][10] = r_cell_wire[911];							inform_R[456][10] = r_cell_wire[912];							inform_R[968][10] = r_cell_wire[913];							inform_R[457][10] = r_cell_wire[914];							inform_R[969][10] = r_cell_wire[915];							inform_R[458][10] = r_cell_wire[916];							inform_R[970][10] = r_cell_wire[917];							inform_R[459][10] = r_cell_wire[918];							inform_R[971][10] = r_cell_wire[919];							inform_R[460][10] = r_cell_wire[920];							inform_R[972][10] = r_cell_wire[921];							inform_R[461][10] = r_cell_wire[922];							inform_R[973][10] = r_cell_wire[923];							inform_R[462][10] = r_cell_wire[924];							inform_R[974][10] = r_cell_wire[925];							inform_R[463][10] = r_cell_wire[926];							inform_R[975][10] = r_cell_wire[927];							inform_R[464][10] = r_cell_wire[928];							inform_R[976][10] = r_cell_wire[929];							inform_R[465][10] = r_cell_wire[930];							inform_R[977][10] = r_cell_wire[931];							inform_R[466][10] = r_cell_wire[932];							inform_R[978][10] = r_cell_wire[933];							inform_R[467][10] = r_cell_wire[934];							inform_R[979][10] = r_cell_wire[935];							inform_R[468][10] = r_cell_wire[936];							inform_R[980][10] = r_cell_wire[937];							inform_R[469][10] = r_cell_wire[938];							inform_R[981][10] = r_cell_wire[939];							inform_R[470][10] = r_cell_wire[940];							inform_R[982][10] = r_cell_wire[941];							inform_R[471][10] = r_cell_wire[942];							inform_R[983][10] = r_cell_wire[943];							inform_R[472][10] = r_cell_wire[944];							inform_R[984][10] = r_cell_wire[945];							inform_R[473][10] = r_cell_wire[946];							inform_R[985][10] = r_cell_wire[947];							inform_R[474][10] = r_cell_wire[948];							inform_R[986][10] = r_cell_wire[949];							inform_R[475][10] = r_cell_wire[950];							inform_R[987][10] = r_cell_wire[951];							inform_R[476][10] = r_cell_wire[952];							inform_R[988][10] = r_cell_wire[953];							inform_R[477][10] = r_cell_wire[954];							inform_R[989][10] = r_cell_wire[955];							inform_R[478][10] = r_cell_wire[956];							inform_R[990][10] = r_cell_wire[957];							inform_R[479][10] = r_cell_wire[958];							inform_R[991][10] = r_cell_wire[959];							inform_R[480][10] = r_cell_wire[960];							inform_R[992][10] = r_cell_wire[961];							inform_R[481][10] = r_cell_wire[962];							inform_R[993][10] = r_cell_wire[963];							inform_R[482][10] = r_cell_wire[964];							inform_R[994][10] = r_cell_wire[965];							inform_R[483][10] = r_cell_wire[966];							inform_R[995][10] = r_cell_wire[967];							inform_R[484][10] = r_cell_wire[968];							inform_R[996][10] = r_cell_wire[969];							inform_R[485][10] = r_cell_wire[970];							inform_R[997][10] = r_cell_wire[971];							inform_R[486][10] = r_cell_wire[972];							inform_R[998][10] = r_cell_wire[973];							inform_R[487][10] = r_cell_wire[974];							inform_R[999][10] = r_cell_wire[975];							inform_R[488][10] = r_cell_wire[976];							inform_R[1000][10] = r_cell_wire[977];							inform_R[489][10] = r_cell_wire[978];							inform_R[1001][10] = r_cell_wire[979];							inform_R[490][10] = r_cell_wire[980];							inform_R[1002][10] = r_cell_wire[981];							inform_R[491][10] = r_cell_wire[982];							inform_R[1003][10] = r_cell_wire[983];							inform_R[492][10] = r_cell_wire[984];							inform_R[1004][10] = r_cell_wire[985];							inform_R[493][10] = r_cell_wire[986];							inform_R[1005][10] = r_cell_wire[987];							inform_R[494][10] = r_cell_wire[988];							inform_R[1006][10] = r_cell_wire[989];							inform_R[495][10] = r_cell_wire[990];							inform_R[1007][10] = r_cell_wire[991];							inform_R[496][10] = r_cell_wire[992];							inform_R[1008][10] = r_cell_wire[993];							inform_R[497][10] = r_cell_wire[994];							inform_R[1009][10] = r_cell_wire[995];							inform_R[498][10] = r_cell_wire[996];							inform_R[1010][10] = r_cell_wire[997];							inform_R[499][10] = r_cell_wire[998];							inform_R[1011][10] = r_cell_wire[999];							inform_R[500][10] = r_cell_wire[1000];							inform_R[1012][10] = r_cell_wire[1001];							inform_R[501][10] = r_cell_wire[1002];							inform_R[1013][10] = r_cell_wire[1003];							inform_R[502][10] = r_cell_wire[1004];							inform_R[1014][10] = r_cell_wire[1005];							inform_R[503][10] = r_cell_wire[1006];							inform_R[1015][10] = r_cell_wire[1007];							inform_R[504][10] = r_cell_wire[1008];							inform_R[1016][10] = r_cell_wire[1009];							inform_R[505][10] = r_cell_wire[1010];							inform_R[1017][10] = r_cell_wire[1011];							inform_R[506][10] = r_cell_wire[1012];							inform_R[1018][10] = r_cell_wire[1013];							inform_R[507][10] = r_cell_wire[1014];							inform_R[1019][10] = r_cell_wire[1015];							inform_R[508][10] = r_cell_wire[1016];							inform_R[1020][10] = r_cell_wire[1017];							inform_R[509][10] = r_cell_wire[1018];							inform_R[1021][10] = r_cell_wire[1019];							inform_R[510][10] = r_cell_wire[1020];							inform_R[1022][10] = r_cell_wire[1021];							inform_R[511][10] = r_cell_wire[1022];							inform_R[1023][10] = r_cell_wire[1023];							inform_L[0][9] = l_cell_wire[0];							inform_L[512][9] = l_cell_wire[1];							inform_L[1][9] = l_cell_wire[2];							inform_L[513][9] = l_cell_wire[3];							inform_L[2][9] = l_cell_wire[4];							inform_L[514][9] = l_cell_wire[5];							inform_L[3][9] = l_cell_wire[6];							inform_L[515][9] = l_cell_wire[7];							inform_L[4][9] = l_cell_wire[8];							inform_L[516][9] = l_cell_wire[9];							inform_L[5][9] = l_cell_wire[10];							inform_L[517][9] = l_cell_wire[11];							inform_L[6][9] = l_cell_wire[12];							inform_L[518][9] = l_cell_wire[13];							inform_L[7][9] = l_cell_wire[14];							inform_L[519][9] = l_cell_wire[15];							inform_L[8][9] = l_cell_wire[16];							inform_L[520][9] = l_cell_wire[17];							inform_L[9][9] = l_cell_wire[18];							inform_L[521][9] = l_cell_wire[19];							inform_L[10][9] = l_cell_wire[20];							inform_L[522][9] = l_cell_wire[21];							inform_L[11][9] = l_cell_wire[22];							inform_L[523][9] = l_cell_wire[23];							inform_L[12][9] = l_cell_wire[24];							inform_L[524][9] = l_cell_wire[25];							inform_L[13][9] = l_cell_wire[26];							inform_L[525][9] = l_cell_wire[27];							inform_L[14][9] = l_cell_wire[28];							inform_L[526][9] = l_cell_wire[29];							inform_L[15][9] = l_cell_wire[30];							inform_L[527][9] = l_cell_wire[31];							inform_L[16][9] = l_cell_wire[32];							inform_L[528][9] = l_cell_wire[33];							inform_L[17][9] = l_cell_wire[34];							inform_L[529][9] = l_cell_wire[35];							inform_L[18][9] = l_cell_wire[36];							inform_L[530][9] = l_cell_wire[37];							inform_L[19][9] = l_cell_wire[38];							inform_L[531][9] = l_cell_wire[39];							inform_L[20][9] = l_cell_wire[40];							inform_L[532][9] = l_cell_wire[41];							inform_L[21][9] = l_cell_wire[42];							inform_L[533][9] = l_cell_wire[43];							inform_L[22][9] = l_cell_wire[44];							inform_L[534][9] = l_cell_wire[45];							inform_L[23][9] = l_cell_wire[46];							inform_L[535][9] = l_cell_wire[47];							inform_L[24][9] = l_cell_wire[48];							inform_L[536][9] = l_cell_wire[49];							inform_L[25][9] = l_cell_wire[50];							inform_L[537][9] = l_cell_wire[51];							inform_L[26][9] = l_cell_wire[52];							inform_L[538][9] = l_cell_wire[53];							inform_L[27][9] = l_cell_wire[54];							inform_L[539][9] = l_cell_wire[55];							inform_L[28][9] = l_cell_wire[56];							inform_L[540][9] = l_cell_wire[57];							inform_L[29][9] = l_cell_wire[58];							inform_L[541][9] = l_cell_wire[59];							inform_L[30][9] = l_cell_wire[60];							inform_L[542][9] = l_cell_wire[61];							inform_L[31][9] = l_cell_wire[62];							inform_L[543][9] = l_cell_wire[63];							inform_L[32][9] = l_cell_wire[64];							inform_L[544][9] = l_cell_wire[65];							inform_L[33][9] = l_cell_wire[66];							inform_L[545][9] = l_cell_wire[67];							inform_L[34][9] = l_cell_wire[68];							inform_L[546][9] = l_cell_wire[69];							inform_L[35][9] = l_cell_wire[70];							inform_L[547][9] = l_cell_wire[71];							inform_L[36][9] = l_cell_wire[72];							inform_L[548][9] = l_cell_wire[73];							inform_L[37][9] = l_cell_wire[74];							inform_L[549][9] = l_cell_wire[75];							inform_L[38][9] = l_cell_wire[76];							inform_L[550][9] = l_cell_wire[77];							inform_L[39][9] = l_cell_wire[78];							inform_L[551][9] = l_cell_wire[79];							inform_L[40][9] = l_cell_wire[80];							inform_L[552][9] = l_cell_wire[81];							inform_L[41][9] = l_cell_wire[82];							inform_L[553][9] = l_cell_wire[83];							inform_L[42][9] = l_cell_wire[84];							inform_L[554][9] = l_cell_wire[85];							inform_L[43][9] = l_cell_wire[86];							inform_L[555][9] = l_cell_wire[87];							inform_L[44][9] = l_cell_wire[88];							inform_L[556][9] = l_cell_wire[89];							inform_L[45][9] = l_cell_wire[90];							inform_L[557][9] = l_cell_wire[91];							inform_L[46][9] = l_cell_wire[92];							inform_L[558][9] = l_cell_wire[93];							inform_L[47][9] = l_cell_wire[94];							inform_L[559][9] = l_cell_wire[95];							inform_L[48][9] = l_cell_wire[96];							inform_L[560][9] = l_cell_wire[97];							inform_L[49][9] = l_cell_wire[98];							inform_L[561][9] = l_cell_wire[99];							inform_L[50][9] = l_cell_wire[100];							inform_L[562][9] = l_cell_wire[101];							inform_L[51][9] = l_cell_wire[102];							inform_L[563][9] = l_cell_wire[103];							inform_L[52][9] = l_cell_wire[104];							inform_L[564][9] = l_cell_wire[105];							inform_L[53][9] = l_cell_wire[106];							inform_L[565][9] = l_cell_wire[107];							inform_L[54][9] = l_cell_wire[108];							inform_L[566][9] = l_cell_wire[109];							inform_L[55][9] = l_cell_wire[110];							inform_L[567][9] = l_cell_wire[111];							inform_L[56][9] = l_cell_wire[112];							inform_L[568][9] = l_cell_wire[113];							inform_L[57][9] = l_cell_wire[114];							inform_L[569][9] = l_cell_wire[115];							inform_L[58][9] = l_cell_wire[116];							inform_L[570][9] = l_cell_wire[117];							inform_L[59][9] = l_cell_wire[118];							inform_L[571][9] = l_cell_wire[119];							inform_L[60][9] = l_cell_wire[120];							inform_L[572][9] = l_cell_wire[121];							inform_L[61][9] = l_cell_wire[122];							inform_L[573][9] = l_cell_wire[123];							inform_L[62][9] = l_cell_wire[124];							inform_L[574][9] = l_cell_wire[125];							inform_L[63][9] = l_cell_wire[126];							inform_L[575][9] = l_cell_wire[127];							inform_L[64][9] = l_cell_wire[128];							inform_L[576][9] = l_cell_wire[129];							inform_L[65][9] = l_cell_wire[130];							inform_L[577][9] = l_cell_wire[131];							inform_L[66][9] = l_cell_wire[132];							inform_L[578][9] = l_cell_wire[133];							inform_L[67][9] = l_cell_wire[134];							inform_L[579][9] = l_cell_wire[135];							inform_L[68][9] = l_cell_wire[136];							inform_L[580][9] = l_cell_wire[137];							inform_L[69][9] = l_cell_wire[138];							inform_L[581][9] = l_cell_wire[139];							inform_L[70][9] = l_cell_wire[140];							inform_L[582][9] = l_cell_wire[141];							inform_L[71][9] = l_cell_wire[142];							inform_L[583][9] = l_cell_wire[143];							inform_L[72][9] = l_cell_wire[144];							inform_L[584][9] = l_cell_wire[145];							inform_L[73][9] = l_cell_wire[146];							inform_L[585][9] = l_cell_wire[147];							inform_L[74][9] = l_cell_wire[148];							inform_L[586][9] = l_cell_wire[149];							inform_L[75][9] = l_cell_wire[150];							inform_L[587][9] = l_cell_wire[151];							inform_L[76][9] = l_cell_wire[152];							inform_L[588][9] = l_cell_wire[153];							inform_L[77][9] = l_cell_wire[154];							inform_L[589][9] = l_cell_wire[155];							inform_L[78][9] = l_cell_wire[156];							inform_L[590][9] = l_cell_wire[157];							inform_L[79][9] = l_cell_wire[158];							inform_L[591][9] = l_cell_wire[159];							inform_L[80][9] = l_cell_wire[160];							inform_L[592][9] = l_cell_wire[161];							inform_L[81][9] = l_cell_wire[162];							inform_L[593][9] = l_cell_wire[163];							inform_L[82][9] = l_cell_wire[164];							inform_L[594][9] = l_cell_wire[165];							inform_L[83][9] = l_cell_wire[166];							inform_L[595][9] = l_cell_wire[167];							inform_L[84][9] = l_cell_wire[168];							inform_L[596][9] = l_cell_wire[169];							inform_L[85][9] = l_cell_wire[170];							inform_L[597][9] = l_cell_wire[171];							inform_L[86][9] = l_cell_wire[172];							inform_L[598][9] = l_cell_wire[173];							inform_L[87][9] = l_cell_wire[174];							inform_L[599][9] = l_cell_wire[175];							inform_L[88][9] = l_cell_wire[176];							inform_L[600][9] = l_cell_wire[177];							inform_L[89][9] = l_cell_wire[178];							inform_L[601][9] = l_cell_wire[179];							inform_L[90][9] = l_cell_wire[180];							inform_L[602][9] = l_cell_wire[181];							inform_L[91][9] = l_cell_wire[182];							inform_L[603][9] = l_cell_wire[183];							inform_L[92][9] = l_cell_wire[184];							inform_L[604][9] = l_cell_wire[185];							inform_L[93][9] = l_cell_wire[186];							inform_L[605][9] = l_cell_wire[187];							inform_L[94][9] = l_cell_wire[188];							inform_L[606][9] = l_cell_wire[189];							inform_L[95][9] = l_cell_wire[190];							inform_L[607][9] = l_cell_wire[191];							inform_L[96][9] = l_cell_wire[192];							inform_L[608][9] = l_cell_wire[193];							inform_L[97][9] = l_cell_wire[194];							inform_L[609][9] = l_cell_wire[195];							inform_L[98][9] = l_cell_wire[196];							inform_L[610][9] = l_cell_wire[197];							inform_L[99][9] = l_cell_wire[198];							inform_L[611][9] = l_cell_wire[199];							inform_L[100][9] = l_cell_wire[200];							inform_L[612][9] = l_cell_wire[201];							inform_L[101][9] = l_cell_wire[202];							inform_L[613][9] = l_cell_wire[203];							inform_L[102][9] = l_cell_wire[204];							inform_L[614][9] = l_cell_wire[205];							inform_L[103][9] = l_cell_wire[206];							inform_L[615][9] = l_cell_wire[207];							inform_L[104][9] = l_cell_wire[208];							inform_L[616][9] = l_cell_wire[209];							inform_L[105][9] = l_cell_wire[210];							inform_L[617][9] = l_cell_wire[211];							inform_L[106][9] = l_cell_wire[212];							inform_L[618][9] = l_cell_wire[213];							inform_L[107][9] = l_cell_wire[214];							inform_L[619][9] = l_cell_wire[215];							inform_L[108][9] = l_cell_wire[216];							inform_L[620][9] = l_cell_wire[217];							inform_L[109][9] = l_cell_wire[218];							inform_L[621][9] = l_cell_wire[219];							inform_L[110][9] = l_cell_wire[220];							inform_L[622][9] = l_cell_wire[221];							inform_L[111][9] = l_cell_wire[222];							inform_L[623][9] = l_cell_wire[223];							inform_L[112][9] = l_cell_wire[224];							inform_L[624][9] = l_cell_wire[225];							inform_L[113][9] = l_cell_wire[226];							inform_L[625][9] = l_cell_wire[227];							inform_L[114][9] = l_cell_wire[228];							inform_L[626][9] = l_cell_wire[229];							inform_L[115][9] = l_cell_wire[230];							inform_L[627][9] = l_cell_wire[231];							inform_L[116][9] = l_cell_wire[232];							inform_L[628][9] = l_cell_wire[233];							inform_L[117][9] = l_cell_wire[234];							inform_L[629][9] = l_cell_wire[235];							inform_L[118][9] = l_cell_wire[236];							inform_L[630][9] = l_cell_wire[237];							inform_L[119][9] = l_cell_wire[238];							inform_L[631][9] = l_cell_wire[239];							inform_L[120][9] = l_cell_wire[240];							inform_L[632][9] = l_cell_wire[241];							inform_L[121][9] = l_cell_wire[242];							inform_L[633][9] = l_cell_wire[243];							inform_L[122][9] = l_cell_wire[244];							inform_L[634][9] = l_cell_wire[245];							inform_L[123][9] = l_cell_wire[246];							inform_L[635][9] = l_cell_wire[247];							inform_L[124][9] = l_cell_wire[248];							inform_L[636][9] = l_cell_wire[249];							inform_L[125][9] = l_cell_wire[250];							inform_L[637][9] = l_cell_wire[251];							inform_L[126][9] = l_cell_wire[252];							inform_L[638][9] = l_cell_wire[253];							inform_L[127][9] = l_cell_wire[254];							inform_L[639][9] = l_cell_wire[255];							inform_L[128][9] = l_cell_wire[256];							inform_L[640][9] = l_cell_wire[257];							inform_L[129][9] = l_cell_wire[258];							inform_L[641][9] = l_cell_wire[259];							inform_L[130][9] = l_cell_wire[260];							inform_L[642][9] = l_cell_wire[261];							inform_L[131][9] = l_cell_wire[262];							inform_L[643][9] = l_cell_wire[263];							inform_L[132][9] = l_cell_wire[264];							inform_L[644][9] = l_cell_wire[265];							inform_L[133][9] = l_cell_wire[266];							inform_L[645][9] = l_cell_wire[267];							inform_L[134][9] = l_cell_wire[268];							inform_L[646][9] = l_cell_wire[269];							inform_L[135][9] = l_cell_wire[270];							inform_L[647][9] = l_cell_wire[271];							inform_L[136][9] = l_cell_wire[272];							inform_L[648][9] = l_cell_wire[273];							inform_L[137][9] = l_cell_wire[274];							inform_L[649][9] = l_cell_wire[275];							inform_L[138][9] = l_cell_wire[276];							inform_L[650][9] = l_cell_wire[277];							inform_L[139][9] = l_cell_wire[278];							inform_L[651][9] = l_cell_wire[279];							inform_L[140][9] = l_cell_wire[280];							inform_L[652][9] = l_cell_wire[281];							inform_L[141][9] = l_cell_wire[282];							inform_L[653][9] = l_cell_wire[283];							inform_L[142][9] = l_cell_wire[284];							inform_L[654][9] = l_cell_wire[285];							inform_L[143][9] = l_cell_wire[286];							inform_L[655][9] = l_cell_wire[287];							inform_L[144][9] = l_cell_wire[288];							inform_L[656][9] = l_cell_wire[289];							inform_L[145][9] = l_cell_wire[290];							inform_L[657][9] = l_cell_wire[291];							inform_L[146][9] = l_cell_wire[292];							inform_L[658][9] = l_cell_wire[293];							inform_L[147][9] = l_cell_wire[294];							inform_L[659][9] = l_cell_wire[295];							inform_L[148][9] = l_cell_wire[296];							inform_L[660][9] = l_cell_wire[297];							inform_L[149][9] = l_cell_wire[298];							inform_L[661][9] = l_cell_wire[299];							inform_L[150][9] = l_cell_wire[300];							inform_L[662][9] = l_cell_wire[301];							inform_L[151][9] = l_cell_wire[302];							inform_L[663][9] = l_cell_wire[303];							inform_L[152][9] = l_cell_wire[304];							inform_L[664][9] = l_cell_wire[305];							inform_L[153][9] = l_cell_wire[306];							inform_L[665][9] = l_cell_wire[307];							inform_L[154][9] = l_cell_wire[308];							inform_L[666][9] = l_cell_wire[309];							inform_L[155][9] = l_cell_wire[310];							inform_L[667][9] = l_cell_wire[311];							inform_L[156][9] = l_cell_wire[312];							inform_L[668][9] = l_cell_wire[313];							inform_L[157][9] = l_cell_wire[314];							inform_L[669][9] = l_cell_wire[315];							inform_L[158][9] = l_cell_wire[316];							inform_L[670][9] = l_cell_wire[317];							inform_L[159][9] = l_cell_wire[318];							inform_L[671][9] = l_cell_wire[319];							inform_L[160][9] = l_cell_wire[320];							inform_L[672][9] = l_cell_wire[321];							inform_L[161][9] = l_cell_wire[322];							inform_L[673][9] = l_cell_wire[323];							inform_L[162][9] = l_cell_wire[324];							inform_L[674][9] = l_cell_wire[325];							inform_L[163][9] = l_cell_wire[326];							inform_L[675][9] = l_cell_wire[327];							inform_L[164][9] = l_cell_wire[328];							inform_L[676][9] = l_cell_wire[329];							inform_L[165][9] = l_cell_wire[330];							inform_L[677][9] = l_cell_wire[331];							inform_L[166][9] = l_cell_wire[332];							inform_L[678][9] = l_cell_wire[333];							inform_L[167][9] = l_cell_wire[334];							inform_L[679][9] = l_cell_wire[335];							inform_L[168][9] = l_cell_wire[336];							inform_L[680][9] = l_cell_wire[337];							inform_L[169][9] = l_cell_wire[338];							inform_L[681][9] = l_cell_wire[339];							inform_L[170][9] = l_cell_wire[340];							inform_L[682][9] = l_cell_wire[341];							inform_L[171][9] = l_cell_wire[342];							inform_L[683][9] = l_cell_wire[343];							inform_L[172][9] = l_cell_wire[344];							inform_L[684][9] = l_cell_wire[345];							inform_L[173][9] = l_cell_wire[346];							inform_L[685][9] = l_cell_wire[347];							inform_L[174][9] = l_cell_wire[348];							inform_L[686][9] = l_cell_wire[349];							inform_L[175][9] = l_cell_wire[350];							inform_L[687][9] = l_cell_wire[351];							inform_L[176][9] = l_cell_wire[352];							inform_L[688][9] = l_cell_wire[353];							inform_L[177][9] = l_cell_wire[354];							inform_L[689][9] = l_cell_wire[355];							inform_L[178][9] = l_cell_wire[356];							inform_L[690][9] = l_cell_wire[357];							inform_L[179][9] = l_cell_wire[358];							inform_L[691][9] = l_cell_wire[359];							inform_L[180][9] = l_cell_wire[360];							inform_L[692][9] = l_cell_wire[361];							inform_L[181][9] = l_cell_wire[362];							inform_L[693][9] = l_cell_wire[363];							inform_L[182][9] = l_cell_wire[364];							inform_L[694][9] = l_cell_wire[365];							inform_L[183][9] = l_cell_wire[366];							inform_L[695][9] = l_cell_wire[367];							inform_L[184][9] = l_cell_wire[368];							inform_L[696][9] = l_cell_wire[369];							inform_L[185][9] = l_cell_wire[370];							inform_L[697][9] = l_cell_wire[371];							inform_L[186][9] = l_cell_wire[372];							inform_L[698][9] = l_cell_wire[373];							inform_L[187][9] = l_cell_wire[374];							inform_L[699][9] = l_cell_wire[375];							inform_L[188][9] = l_cell_wire[376];							inform_L[700][9] = l_cell_wire[377];							inform_L[189][9] = l_cell_wire[378];							inform_L[701][9] = l_cell_wire[379];							inform_L[190][9] = l_cell_wire[380];							inform_L[702][9] = l_cell_wire[381];							inform_L[191][9] = l_cell_wire[382];							inform_L[703][9] = l_cell_wire[383];							inform_L[192][9] = l_cell_wire[384];							inform_L[704][9] = l_cell_wire[385];							inform_L[193][9] = l_cell_wire[386];							inform_L[705][9] = l_cell_wire[387];							inform_L[194][9] = l_cell_wire[388];							inform_L[706][9] = l_cell_wire[389];							inform_L[195][9] = l_cell_wire[390];							inform_L[707][9] = l_cell_wire[391];							inform_L[196][9] = l_cell_wire[392];							inform_L[708][9] = l_cell_wire[393];							inform_L[197][9] = l_cell_wire[394];							inform_L[709][9] = l_cell_wire[395];							inform_L[198][9] = l_cell_wire[396];							inform_L[710][9] = l_cell_wire[397];							inform_L[199][9] = l_cell_wire[398];							inform_L[711][9] = l_cell_wire[399];							inform_L[200][9] = l_cell_wire[400];							inform_L[712][9] = l_cell_wire[401];							inform_L[201][9] = l_cell_wire[402];							inform_L[713][9] = l_cell_wire[403];							inform_L[202][9] = l_cell_wire[404];							inform_L[714][9] = l_cell_wire[405];							inform_L[203][9] = l_cell_wire[406];							inform_L[715][9] = l_cell_wire[407];							inform_L[204][9] = l_cell_wire[408];							inform_L[716][9] = l_cell_wire[409];							inform_L[205][9] = l_cell_wire[410];							inform_L[717][9] = l_cell_wire[411];							inform_L[206][9] = l_cell_wire[412];							inform_L[718][9] = l_cell_wire[413];							inform_L[207][9] = l_cell_wire[414];							inform_L[719][9] = l_cell_wire[415];							inform_L[208][9] = l_cell_wire[416];							inform_L[720][9] = l_cell_wire[417];							inform_L[209][9] = l_cell_wire[418];							inform_L[721][9] = l_cell_wire[419];							inform_L[210][9] = l_cell_wire[420];							inform_L[722][9] = l_cell_wire[421];							inform_L[211][9] = l_cell_wire[422];							inform_L[723][9] = l_cell_wire[423];							inform_L[212][9] = l_cell_wire[424];							inform_L[724][9] = l_cell_wire[425];							inform_L[213][9] = l_cell_wire[426];							inform_L[725][9] = l_cell_wire[427];							inform_L[214][9] = l_cell_wire[428];							inform_L[726][9] = l_cell_wire[429];							inform_L[215][9] = l_cell_wire[430];							inform_L[727][9] = l_cell_wire[431];							inform_L[216][9] = l_cell_wire[432];							inform_L[728][9] = l_cell_wire[433];							inform_L[217][9] = l_cell_wire[434];							inform_L[729][9] = l_cell_wire[435];							inform_L[218][9] = l_cell_wire[436];							inform_L[730][9] = l_cell_wire[437];							inform_L[219][9] = l_cell_wire[438];							inform_L[731][9] = l_cell_wire[439];							inform_L[220][9] = l_cell_wire[440];							inform_L[732][9] = l_cell_wire[441];							inform_L[221][9] = l_cell_wire[442];							inform_L[733][9] = l_cell_wire[443];							inform_L[222][9] = l_cell_wire[444];							inform_L[734][9] = l_cell_wire[445];							inform_L[223][9] = l_cell_wire[446];							inform_L[735][9] = l_cell_wire[447];							inform_L[224][9] = l_cell_wire[448];							inform_L[736][9] = l_cell_wire[449];							inform_L[225][9] = l_cell_wire[450];							inform_L[737][9] = l_cell_wire[451];							inform_L[226][9] = l_cell_wire[452];							inform_L[738][9] = l_cell_wire[453];							inform_L[227][9] = l_cell_wire[454];							inform_L[739][9] = l_cell_wire[455];							inform_L[228][9] = l_cell_wire[456];							inform_L[740][9] = l_cell_wire[457];							inform_L[229][9] = l_cell_wire[458];							inform_L[741][9] = l_cell_wire[459];							inform_L[230][9] = l_cell_wire[460];							inform_L[742][9] = l_cell_wire[461];							inform_L[231][9] = l_cell_wire[462];							inform_L[743][9] = l_cell_wire[463];							inform_L[232][9] = l_cell_wire[464];							inform_L[744][9] = l_cell_wire[465];							inform_L[233][9] = l_cell_wire[466];							inform_L[745][9] = l_cell_wire[467];							inform_L[234][9] = l_cell_wire[468];							inform_L[746][9] = l_cell_wire[469];							inform_L[235][9] = l_cell_wire[470];							inform_L[747][9] = l_cell_wire[471];							inform_L[236][9] = l_cell_wire[472];							inform_L[748][9] = l_cell_wire[473];							inform_L[237][9] = l_cell_wire[474];							inform_L[749][9] = l_cell_wire[475];							inform_L[238][9] = l_cell_wire[476];							inform_L[750][9] = l_cell_wire[477];							inform_L[239][9] = l_cell_wire[478];							inform_L[751][9] = l_cell_wire[479];							inform_L[240][9] = l_cell_wire[480];							inform_L[752][9] = l_cell_wire[481];							inform_L[241][9] = l_cell_wire[482];							inform_L[753][9] = l_cell_wire[483];							inform_L[242][9] = l_cell_wire[484];							inform_L[754][9] = l_cell_wire[485];							inform_L[243][9] = l_cell_wire[486];							inform_L[755][9] = l_cell_wire[487];							inform_L[244][9] = l_cell_wire[488];							inform_L[756][9] = l_cell_wire[489];							inform_L[245][9] = l_cell_wire[490];							inform_L[757][9] = l_cell_wire[491];							inform_L[246][9] = l_cell_wire[492];							inform_L[758][9] = l_cell_wire[493];							inform_L[247][9] = l_cell_wire[494];							inform_L[759][9] = l_cell_wire[495];							inform_L[248][9] = l_cell_wire[496];							inform_L[760][9] = l_cell_wire[497];							inform_L[249][9] = l_cell_wire[498];							inform_L[761][9] = l_cell_wire[499];							inform_L[250][9] = l_cell_wire[500];							inform_L[762][9] = l_cell_wire[501];							inform_L[251][9] = l_cell_wire[502];							inform_L[763][9] = l_cell_wire[503];							inform_L[252][9] = l_cell_wire[504];							inform_L[764][9] = l_cell_wire[505];							inform_L[253][9] = l_cell_wire[506];							inform_L[765][9] = l_cell_wire[507];							inform_L[254][9] = l_cell_wire[508];							inform_L[766][9] = l_cell_wire[509];							inform_L[255][9] = l_cell_wire[510];							inform_L[767][9] = l_cell_wire[511];							inform_L[256][9] = l_cell_wire[512];							inform_L[768][9] = l_cell_wire[513];							inform_L[257][9] = l_cell_wire[514];							inform_L[769][9] = l_cell_wire[515];							inform_L[258][9] = l_cell_wire[516];							inform_L[770][9] = l_cell_wire[517];							inform_L[259][9] = l_cell_wire[518];							inform_L[771][9] = l_cell_wire[519];							inform_L[260][9] = l_cell_wire[520];							inform_L[772][9] = l_cell_wire[521];							inform_L[261][9] = l_cell_wire[522];							inform_L[773][9] = l_cell_wire[523];							inform_L[262][9] = l_cell_wire[524];							inform_L[774][9] = l_cell_wire[525];							inform_L[263][9] = l_cell_wire[526];							inform_L[775][9] = l_cell_wire[527];							inform_L[264][9] = l_cell_wire[528];							inform_L[776][9] = l_cell_wire[529];							inform_L[265][9] = l_cell_wire[530];							inform_L[777][9] = l_cell_wire[531];							inform_L[266][9] = l_cell_wire[532];							inform_L[778][9] = l_cell_wire[533];							inform_L[267][9] = l_cell_wire[534];							inform_L[779][9] = l_cell_wire[535];							inform_L[268][9] = l_cell_wire[536];							inform_L[780][9] = l_cell_wire[537];							inform_L[269][9] = l_cell_wire[538];							inform_L[781][9] = l_cell_wire[539];							inform_L[270][9] = l_cell_wire[540];							inform_L[782][9] = l_cell_wire[541];							inform_L[271][9] = l_cell_wire[542];							inform_L[783][9] = l_cell_wire[543];							inform_L[272][9] = l_cell_wire[544];							inform_L[784][9] = l_cell_wire[545];							inform_L[273][9] = l_cell_wire[546];							inform_L[785][9] = l_cell_wire[547];							inform_L[274][9] = l_cell_wire[548];							inform_L[786][9] = l_cell_wire[549];							inform_L[275][9] = l_cell_wire[550];							inform_L[787][9] = l_cell_wire[551];							inform_L[276][9] = l_cell_wire[552];							inform_L[788][9] = l_cell_wire[553];							inform_L[277][9] = l_cell_wire[554];							inform_L[789][9] = l_cell_wire[555];							inform_L[278][9] = l_cell_wire[556];							inform_L[790][9] = l_cell_wire[557];							inform_L[279][9] = l_cell_wire[558];							inform_L[791][9] = l_cell_wire[559];							inform_L[280][9] = l_cell_wire[560];							inform_L[792][9] = l_cell_wire[561];							inform_L[281][9] = l_cell_wire[562];							inform_L[793][9] = l_cell_wire[563];							inform_L[282][9] = l_cell_wire[564];							inform_L[794][9] = l_cell_wire[565];							inform_L[283][9] = l_cell_wire[566];							inform_L[795][9] = l_cell_wire[567];							inform_L[284][9] = l_cell_wire[568];							inform_L[796][9] = l_cell_wire[569];							inform_L[285][9] = l_cell_wire[570];							inform_L[797][9] = l_cell_wire[571];							inform_L[286][9] = l_cell_wire[572];							inform_L[798][9] = l_cell_wire[573];							inform_L[287][9] = l_cell_wire[574];							inform_L[799][9] = l_cell_wire[575];							inform_L[288][9] = l_cell_wire[576];							inform_L[800][9] = l_cell_wire[577];							inform_L[289][9] = l_cell_wire[578];							inform_L[801][9] = l_cell_wire[579];							inform_L[290][9] = l_cell_wire[580];							inform_L[802][9] = l_cell_wire[581];							inform_L[291][9] = l_cell_wire[582];							inform_L[803][9] = l_cell_wire[583];							inform_L[292][9] = l_cell_wire[584];							inform_L[804][9] = l_cell_wire[585];							inform_L[293][9] = l_cell_wire[586];							inform_L[805][9] = l_cell_wire[587];							inform_L[294][9] = l_cell_wire[588];							inform_L[806][9] = l_cell_wire[589];							inform_L[295][9] = l_cell_wire[590];							inform_L[807][9] = l_cell_wire[591];							inform_L[296][9] = l_cell_wire[592];							inform_L[808][9] = l_cell_wire[593];							inform_L[297][9] = l_cell_wire[594];							inform_L[809][9] = l_cell_wire[595];							inform_L[298][9] = l_cell_wire[596];							inform_L[810][9] = l_cell_wire[597];							inform_L[299][9] = l_cell_wire[598];							inform_L[811][9] = l_cell_wire[599];							inform_L[300][9] = l_cell_wire[600];							inform_L[812][9] = l_cell_wire[601];							inform_L[301][9] = l_cell_wire[602];							inform_L[813][9] = l_cell_wire[603];							inform_L[302][9] = l_cell_wire[604];							inform_L[814][9] = l_cell_wire[605];							inform_L[303][9] = l_cell_wire[606];							inform_L[815][9] = l_cell_wire[607];							inform_L[304][9] = l_cell_wire[608];							inform_L[816][9] = l_cell_wire[609];							inform_L[305][9] = l_cell_wire[610];							inform_L[817][9] = l_cell_wire[611];							inform_L[306][9] = l_cell_wire[612];							inform_L[818][9] = l_cell_wire[613];							inform_L[307][9] = l_cell_wire[614];							inform_L[819][9] = l_cell_wire[615];							inform_L[308][9] = l_cell_wire[616];							inform_L[820][9] = l_cell_wire[617];							inform_L[309][9] = l_cell_wire[618];							inform_L[821][9] = l_cell_wire[619];							inform_L[310][9] = l_cell_wire[620];							inform_L[822][9] = l_cell_wire[621];							inform_L[311][9] = l_cell_wire[622];							inform_L[823][9] = l_cell_wire[623];							inform_L[312][9] = l_cell_wire[624];							inform_L[824][9] = l_cell_wire[625];							inform_L[313][9] = l_cell_wire[626];							inform_L[825][9] = l_cell_wire[627];							inform_L[314][9] = l_cell_wire[628];							inform_L[826][9] = l_cell_wire[629];							inform_L[315][9] = l_cell_wire[630];							inform_L[827][9] = l_cell_wire[631];							inform_L[316][9] = l_cell_wire[632];							inform_L[828][9] = l_cell_wire[633];							inform_L[317][9] = l_cell_wire[634];							inform_L[829][9] = l_cell_wire[635];							inform_L[318][9] = l_cell_wire[636];							inform_L[830][9] = l_cell_wire[637];							inform_L[319][9] = l_cell_wire[638];							inform_L[831][9] = l_cell_wire[639];							inform_L[320][9] = l_cell_wire[640];							inform_L[832][9] = l_cell_wire[641];							inform_L[321][9] = l_cell_wire[642];							inform_L[833][9] = l_cell_wire[643];							inform_L[322][9] = l_cell_wire[644];							inform_L[834][9] = l_cell_wire[645];							inform_L[323][9] = l_cell_wire[646];							inform_L[835][9] = l_cell_wire[647];							inform_L[324][9] = l_cell_wire[648];							inform_L[836][9] = l_cell_wire[649];							inform_L[325][9] = l_cell_wire[650];							inform_L[837][9] = l_cell_wire[651];							inform_L[326][9] = l_cell_wire[652];							inform_L[838][9] = l_cell_wire[653];							inform_L[327][9] = l_cell_wire[654];							inform_L[839][9] = l_cell_wire[655];							inform_L[328][9] = l_cell_wire[656];							inform_L[840][9] = l_cell_wire[657];							inform_L[329][9] = l_cell_wire[658];							inform_L[841][9] = l_cell_wire[659];							inform_L[330][9] = l_cell_wire[660];							inform_L[842][9] = l_cell_wire[661];							inform_L[331][9] = l_cell_wire[662];							inform_L[843][9] = l_cell_wire[663];							inform_L[332][9] = l_cell_wire[664];							inform_L[844][9] = l_cell_wire[665];							inform_L[333][9] = l_cell_wire[666];							inform_L[845][9] = l_cell_wire[667];							inform_L[334][9] = l_cell_wire[668];							inform_L[846][9] = l_cell_wire[669];							inform_L[335][9] = l_cell_wire[670];							inform_L[847][9] = l_cell_wire[671];							inform_L[336][9] = l_cell_wire[672];							inform_L[848][9] = l_cell_wire[673];							inform_L[337][9] = l_cell_wire[674];							inform_L[849][9] = l_cell_wire[675];							inform_L[338][9] = l_cell_wire[676];							inform_L[850][9] = l_cell_wire[677];							inform_L[339][9] = l_cell_wire[678];							inform_L[851][9] = l_cell_wire[679];							inform_L[340][9] = l_cell_wire[680];							inform_L[852][9] = l_cell_wire[681];							inform_L[341][9] = l_cell_wire[682];							inform_L[853][9] = l_cell_wire[683];							inform_L[342][9] = l_cell_wire[684];							inform_L[854][9] = l_cell_wire[685];							inform_L[343][9] = l_cell_wire[686];							inform_L[855][9] = l_cell_wire[687];							inform_L[344][9] = l_cell_wire[688];							inform_L[856][9] = l_cell_wire[689];							inform_L[345][9] = l_cell_wire[690];							inform_L[857][9] = l_cell_wire[691];							inform_L[346][9] = l_cell_wire[692];							inform_L[858][9] = l_cell_wire[693];							inform_L[347][9] = l_cell_wire[694];							inform_L[859][9] = l_cell_wire[695];							inform_L[348][9] = l_cell_wire[696];							inform_L[860][9] = l_cell_wire[697];							inform_L[349][9] = l_cell_wire[698];							inform_L[861][9] = l_cell_wire[699];							inform_L[350][9] = l_cell_wire[700];							inform_L[862][9] = l_cell_wire[701];							inform_L[351][9] = l_cell_wire[702];							inform_L[863][9] = l_cell_wire[703];							inform_L[352][9] = l_cell_wire[704];							inform_L[864][9] = l_cell_wire[705];							inform_L[353][9] = l_cell_wire[706];							inform_L[865][9] = l_cell_wire[707];							inform_L[354][9] = l_cell_wire[708];							inform_L[866][9] = l_cell_wire[709];							inform_L[355][9] = l_cell_wire[710];							inform_L[867][9] = l_cell_wire[711];							inform_L[356][9] = l_cell_wire[712];							inform_L[868][9] = l_cell_wire[713];							inform_L[357][9] = l_cell_wire[714];							inform_L[869][9] = l_cell_wire[715];							inform_L[358][9] = l_cell_wire[716];							inform_L[870][9] = l_cell_wire[717];							inform_L[359][9] = l_cell_wire[718];							inform_L[871][9] = l_cell_wire[719];							inform_L[360][9] = l_cell_wire[720];							inform_L[872][9] = l_cell_wire[721];							inform_L[361][9] = l_cell_wire[722];							inform_L[873][9] = l_cell_wire[723];							inform_L[362][9] = l_cell_wire[724];							inform_L[874][9] = l_cell_wire[725];							inform_L[363][9] = l_cell_wire[726];							inform_L[875][9] = l_cell_wire[727];							inform_L[364][9] = l_cell_wire[728];							inform_L[876][9] = l_cell_wire[729];							inform_L[365][9] = l_cell_wire[730];							inform_L[877][9] = l_cell_wire[731];							inform_L[366][9] = l_cell_wire[732];							inform_L[878][9] = l_cell_wire[733];							inform_L[367][9] = l_cell_wire[734];							inform_L[879][9] = l_cell_wire[735];							inform_L[368][9] = l_cell_wire[736];							inform_L[880][9] = l_cell_wire[737];							inform_L[369][9] = l_cell_wire[738];							inform_L[881][9] = l_cell_wire[739];							inform_L[370][9] = l_cell_wire[740];							inform_L[882][9] = l_cell_wire[741];							inform_L[371][9] = l_cell_wire[742];							inform_L[883][9] = l_cell_wire[743];							inform_L[372][9] = l_cell_wire[744];							inform_L[884][9] = l_cell_wire[745];							inform_L[373][9] = l_cell_wire[746];							inform_L[885][9] = l_cell_wire[747];							inform_L[374][9] = l_cell_wire[748];							inform_L[886][9] = l_cell_wire[749];							inform_L[375][9] = l_cell_wire[750];							inform_L[887][9] = l_cell_wire[751];							inform_L[376][9] = l_cell_wire[752];							inform_L[888][9] = l_cell_wire[753];							inform_L[377][9] = l_cell_wire[754];							inform_L[889][9] = l_cell_wire[755];							inform_L[378][9] = l_cell_wire[756];							inform_L[890][9] = l_cell_wire[757];							inform_L[379][9] = l_cell_wire[758];							inform_L[891][9] = l_cell_wire[759];							inform_L[380][9] = l_cell_wire[760];							inform_L[892][9] = l_cell_wire[761];							inform_L[381][9] = l_cell_wire[762];							inform_L[893][9] = l_cell_wire[763];							inform_L[382][9] = l_cell_wire[764];							inform_L[894][9] = l_cell_wire[765];							inform_L[383][9] = l_cell_wire[766];							inform_L[895][9] = l_cell_wire[767];							inform_L[384][9] = l_cell_wire[768];							inform_L[896][9] = l_cell_wire[769];							inform_L[385][9] = l_cell_wire[770];							inform_L[897][9] = l_cell_wire[771];							inform_L[386][9] = l_cell_wire[772];							inform_L[898][9] = l_cell_wire[773];							inform_L[387][9] = l_cell_wire[774];							inform_L[899][9] = l_cell_wire[775];							inform_L[388][9] = l_cell_wire[776];							inform_L[900][9] = l_cell_wire[777];							inform_L[389][9] = l_cell_wire[778];							inform_L[901][9] = l_cell_wire[779];							inform_L[390][9] = l_cell_wire[780];							inform_L[902][9] = l_cell_wire[781];							inform_L[391][9] = l_cell_wire[782];							inform_L[903][9] = l_cell_wire[783];							inform_L[392][9] = l_cell_wire[784];							inform_L[904][9] = l_cell_wire[785];							inform_L[393][9] = l_cell_wire[786];							inform_L[905][9] = l_cell_wire[787];							inform_L[394][9] = l_cell_wire[788];							inform_L[906][9] = l_cell_wire[789];							inform_L[395][9] = l_cell_wire[790];							inform_L[907][9] = l_cell_wire[791];							inform_L[396][9] = l_cell_wire[792];							inform_L[908][9] = l_cell_wire[793];							inform_L[397][9] = l_cell_wire[794];							inform_L[909][9] = l_cell_wire[795];							inform_L[398][9] = l_cell_wire[796];							inform_L[910][9] = l_cell_wire[797];							inform_L[399][9] = l_cell_wire[798];							inform_L[911][9] = l_cell_wire[799];							inform_L[400][9] = l_cell_wire[800];							inform_L[912][9] = l_cell_wire[801];							inform_L[401][9] = l_cell_wire[802];							inform_L[913][9] = l_cell_wire[803];							inform_L[402][9] = l_cell_wire[804];							inform_L[914][9] = l_cell_wire[805];							inform_L[403][9] = l_cell_wire[806];							inform_L[915][9] = l_cell_wire[807];							inform_L[404][9] = l_cell_wire[808];							inform_L[916][9] = l_cell_wire[809];							inform_L[405][9] = l_cell_wire[810];							inform_L[917][9] = l_cell_wire[811];							inform_L[406][9] = l_cell_wire[812];							inform_L[918][9] = l_cell_wire[813];							inform_L[407][9] = l_cell_wire[814];							inform_L[919][9] = l_cell_wire[815];							inform_L[408][9] = l_cell_wire[816];							inform_L[920][9] = l_cell_wire[817];							inform_L[409][9] = l_cell_wire[818];							inform_L[921][9] = l_cell_wire[819];							inform_L[410][9] = l_cell_wire[820];							inform_L[922][9] = l_cell_wire[821];							inform_L[411][9] = l_cell_wire[822];							inform_L[923][9] = l_cell_wire[823];							inform_L[412][9] = l_cell_wire[824];							inform_L[924][9] = l_cell_wire[825];							inform_L[413][9] = l_cell_wire[826];							inform_L[925][9] = l_cell_wire[827];							inform_L[414][9] = l_cell_wire[828];							inform_L[926][9] = l_cell_wire[829];							inform_L[415][9] = l_cell_wire[830];							inform_L[927][9] = l_cell_wire[831];							inform_L[416][9] = l_cell_wire[832];							inform_L[928][9] = l_cell_wire[833];							inform_L[417][9] = l_cell_wire[834];							inform_L[929][9] = l_cell_wire[835];							inform_L[418][9] = l_cell_wire[836];							inform_L[930][9] = l_cell_wire[837];							inform_L[419][9] = l_cell_wire[838];							inform_L[931][9] = l_cell_wire[839];							inform_L[420][9] = l_cell_wire[840];							inform_L[932][9] = l_cell_wire[841];							inform_L[421][9] = l_cell_wire[842];							inform_L[933][9] = l_cell_wire[843];							inform_L[422][9] = l_cell_wire[844];							inform_L[934][9] = l_cell_wire[845];							inform_L[423][9] = l_cell_wire[846];							inform_L[935][9] = l_cell_wire[847];							inform_L[424][9] = l_cell_wire[848];							inform_L[936][9] = l_cell_wire[849];							inform_L[425][9] = l_cell_wire[850];							inform_L[937][9] = l_cell_wire[851];							inform_L[426][9] = l_cell_wire[852];							inform_L[938][9] = l_cell_wire[853];							inform_L[427][9] = l_cell_wire[854];							inform_L[939][9] = l_cell_wire[855];							inform_L[428][9] = l_cell_wire[856];							inform_L[940][9] = l_cell_wire[857];							inform_L[429][9] = l_cell_wire[858];							inform_L[941][9] = l_cell_wire[859];							inform_L[430][9] = l_cell_wire[860];							inform_L[942][9] = l_cell_wire[861];							inform_L[431][9] = l_cell_wire[862];							inform_L[943][9] = l_cell_wire[863];							inform_L[432][9] = l_cell_wire[864];							inform_L[944][9] = l_cell_wire[865];							inform_L[433][9] = l_cell_wire[866];							inform_L[945][9] = l_cell_wire[867];							inform_L[434][9] = l_cell_wire[868];							inform_L[946][9] = l_cell_wire[869];							inform_L[435][9] = l_cell_wire[870];							inform_L[947][9] = l_cell_wire[871];							inform_L[436][9] = l_cell_wire[872];							inform_L[948][9] = l_cell_wire[873];							inform_L[437][9] = l_cell_wire[874];							inform_L[949][9] = l_cell_wire[875];							inform_L[438][9] = l_cell_wire[876];							inform_L[950][9] = l_cell_wire[877];							inform_L[439][9] = l_cell_wire[878];							inform_L[951][9] = l_cell_wire[879];							inform_L[440][9] = l_cell_wire[880];							inform_L[952][9] = l_cell_wire[881];							inform_L[441][9] = l_cell_wire[882];							inform_L[953][9] = l_cell_wire[883];							inform_L[442][9] = l_cell_wire[884];							inform_L[954][9] = l_cell_wire[885];							inform_L[443][9] = l_cell_wire[886];							inform_L[955][9] = l_cell_wire[887];							inform_L[444][9] = l_cell_wire[888];							inform_L[956][9] = l_cell_wire[889];							inform_L[445][9] = l_cell_wire[890];							inform_L[957][9] = l_cell_wire[891];							inform_L[446][9] = l_cell_wire[892];							inform_L[958][9] = l_cell_wire[893];							inform_L[447][9] = l_cell_wire[894];							inform_L[959][9] = l_cell_wire[895];							inform_L[448][9] = l_cell_wire[896];							inform_L[960][9] = l_cell_wire[897];							inform_L[449][9] = l_cell_wire[898];							inform_L[961][9] = l_cell_wire[899];							inform_L[450][9] = l_cell_wire[900];							inform_L[962][9] = l_cell_wire[901];							inform_L[451][9] = l_cell_wire[902];							inform_L[963][9] = l_cell_wire[903];							inform_L[452][9] = l_cell_wire[904];							inform_L[964][9] = l_cell_wire[905];							inform_L[453][9] = l_cell_wire[906];							inform_L[965][9] = l_cell_wire[907];							inform_L[454][9] = l_cell_wire[908];							inform_L[966][9] = l_cell_wire[909];							inform_L[455][9] = l_cell_wire[910];							inform_L[967][9] = l_cell_wire[911];							inform_L[456][9] = l_cell_wire[912];							inform_L[968][9] = l_cell_wire[913];							inform_L[457][9] = l_cell_wire[914];							inform_L[969][9] = l_cell_wire[915];							inform_L[458][9] = l_cell_wire[916];							inform_L[970][9] = l_cell_wire[917];							inform_L[459][9] = l_cell_wire[918];							inform_L[971][9] = l_cell_wire[919];							inform_L[460][9] = l_cell_wire[920];							inform_L[972][9] = l_cell_wire[921];							inform_L[461][9] = l_cell_wire[922];							inform_L[973][9] = l_cell_wire[923];							inform_L[462][9] = l_cell_wire[924];							inform_L[974][9] = l_cell_wire[925];							inform_L[463][9] = l_cell_wire[926];							inform_L[975][9] = l_cell_wire[927];							inform_L[464][9] = l_cell_wire[928];							inform_L[976][9] = l_cell_wire[929];							inform_L[465][9] = l_cell_wire[930];							inform_L[977][9] = l_cell_wire[931];							inform_L[466][9] = l_cell_wire[932];							inform_L[978][9] = l_cell_wire[933];							inform_L[467][9] = l_cell_wire[934];							inform_L[979][9] = l_cell_wire[935];							inform_L[468][9] = l_cell_wire[936];							inform_L[980][9] = l_cell_wire[937];							inform_L[469][9] = l_cell_wire[938];							inform_L[981][9] = l_cell_wire[939];							inform_L[470][9] = l_cell_wire[940];							inform_L[982][9] = l_cell_wire[941];							inform_L[471][9] = l_cell_wire[942];							inform_L[983][9] = l_cell_wire[943];							inform_L[472][9] = l_cell_wire[944];							inform_L[984][9] = l_cell_wire[945];							inform_L[473][9] = l_cell_wire[946];							inform_L[985][9] = l_cell_wire[947];							inform_L[474][9] = l_cell_wire[948];							inform_L[986][9] = l_cell_wire[949];							inform_L[475][9] = l_cell_wire[950];							inform_L[987][9] = l_cell_wire[951];							inform_L[476][9] = l_cell_wire[952];							inform_L[988][9] = l_cell_wire[953];							inform_L[477][9] = l_cell_wire[954];							inform_L[989][9] = l_cell_wire[955];							inform_L[478][9] = l_cell_wire[956];							inform_L[990][9] = l_cell_wire[957];							inform_L[479][9] = l_cell_wire[958];							inform_L[991][9] = l_cell_wire[959];							inform_L[480][9] = l_cell_wire[960];							inform_L[992][9] = l_cell_wire[961];							inform_L[481][9] = l_cell_wire[962];							inform_L[993][9] = l_cell_wire[963];							inform_L[482][9] = l_cell_wire[964];							inform_L[994][9] = l_cell_wire[965];							inform_L[483][9] = l_cell_wire[966];							inform_L[995][9] = l_cell_wire[967];							inform_L[484][9] = l_cell_wire[968];							inform_L[996][9] = l_cell_wire[969];							inform_L[485][9] = l_cell_wire[970];							inform_L[997][9] = l_cell_wire[971];							inform_L[486][9] = l_cell_wire[972];							inform_L[998][9] = l_cell_wire[973];							inform_L[487][9] = l_cell_wire[974];							inform_L[999][9] = l_cell_wire[975];							inform_L[488][9] = l_cell_wire[976];							inform_L[1000][9] = l_cell_wire[977];							inform_L[489][9] = l_cell_wire[978];							inform_L[1001][9] = l_cell_wire[979];							inform_L[490][9] = l_cell_wire[980];							inform_L[1002][9] = l_cell_wire[981];							inform_L[491][9] = l_cell_wire[982];							inform_L[1003][9] = l_cell_wire[983];							inform_L[492][9] = l_cell_wire[984];							inform_L[1004][9] = l_cell_wire[985];							inform_L[493][9] = l_cell_wire[986];							inform_L[1005][9] = l_cell_wire[987];							inform_L[494][9] = l_cell_wire[988];							inform_L[1006][9] = l_cell_wire[989];							inform_L[495][9] = l_cell_wire[990];							inform_L[1007][9] = l_cell_wire[991];							inform_L[496][9] = l_cell_wire[992];							inform_L[1008][9] = l_cell_wire[993];							inform_L[497][9] = l_cell_wire[994];							inform_L[1009][9] = l_cell_wire[995];							inform_L[498][9] = l_cell_wire[996];							inform_L[1010][9] = l_cell_wire[997];							inform_L[499][9] = l_cell_wire[998];							inform_L[1011][9] = l_cell_wire[999];							inform_L[500][9] = l_cell_wire[1000];							inform_L[1012][9] = l_cell_wire[1001];							inform_L[501][9] = l_cell_wire[1002];							inform_L[1013][9] = l_cell_wire[1003];							inform_L[502][9] = l_cell_wire[1004];							inform_L[1014][9] = l_cell_wire[1005];							inform_L[503][9] = l_cell_wire[1006];							inform_L[1015][9] = l_cell_wire[1007];							inform_L[504][9] = l_cell_wire[1008];							inform_L[1016][9] = l_cell_wire[1009];							inform_L[505][9] = l_cell_wire[1010];							inform_L[1017][9] = l_cell_wire[1011];							inform_L[506][9] = l_cell_wire[1012];							inform_L[1018][9] = l_cell_wire[1013];							inform_L[507][9] = l_cell_wire[1014];							inform_L[1019][9] = l_cell_wire[1015];							inform_L[508][9] = l_cell_wire[1016];							inform_L[1020][9] = l_cell_wire[1017];							inform_L[509][9] = l_cell_wire[1018];							inform_L[1021][9] = l_cell_wire[1019];							inform_L[510][9] = l_cell_wire[1020];							inform_L[1022][9] = l_cell_wire[1021];							inform_L[511][9] = l_cell_wire[1022];							inform_L[1023][9] = l_cell_wire[1023];						end
						default:							for (x = 0; x < 1024; x = x + 1)								for (y = 0; y < 10; y = y + 1)								begin									inform_R[x][y+1] <= 8'd0;									inform_L[x][y] <= 8'd0;								end					endcase				end			end
				default:				begin				if (start) begin					inform_R [0][0] <= 8'b0111_1111;					inform_R [1][0] <= 8'b0111_1111;					inform_R [2][0] <= 8'b0111_1111;					inform_R [3][0] <= 8'b0111_1111;					inform_R [4][0] <= 8'b0111_1111;					inform_R [5][0] <= 8'b0111_1111;					inform_R [6][0] <= 8'b0111_1111;					inform_R [7][0] <= 8'b0111_1111;					inform_R [8][0] <= 8'b0111_1111;					inform_R [9][0] <= 8'b0111_1111;					inform_R [10][0] <= 8'b0111_1111;					inform_R [11][0] <= 8'b0111_1111;					inform_R [12][0] <= 8'b0111_1111;					inform_R [13][0] <= 8'b0111_1111;					inform_R [14][0] <= 8'b0111_1111;					inform_R [15][0] <= 8'b0111_1111;					inform_R [16][0] <= 8'b0111_1111;					inform_R [17][0] <= 8'b0111_1111;					inform_R [18][0] <= 8'b0111_1111;					inform_R [19][0] <= 8'b0111_1111;					inform_R [20][0] <= 8'b0111_1111;					inform_R [21][0] <= 8'b0111_1111;					inform_R [22][0] <= 8'b0111_1111;					inform_R [23][0] <= 8'b0111_1111;					inform_R [24][0] <= 8'b0111_1111;					inform_R [25][0] <= 8'b0111_1111;					inform_R [26][0] <= 8'b0111_1111;					inform_R [27][0] <= 8'b0111_1111;					inform_R [28][0] <= 8'b0111_1111;					inform_R [29][0] <= 8'b0111_1111;					inform_R [30][0] <= 8'b0111_1111;					inform_R [31][0] <= 8'b0111_1111;					inform_R [32][0] <= 8'b0111_1111;					inform_R [33][0] <= 8'b0111_1111;					inform_R [34][0] <= 8'b0111_1111;					inform_R [35][0] <= 8'b0111_1111;					inform_R [36][0] <= 8'b0111_1111;					inform_R [37][0] <= 8'b0111_1111;					inform_R [38][0] <= 8'b0111_1111;					inform_R [39][0] <= 8'b0111_1111;					inform_R [40][0] <= 8'b0111_1111;					inform_R [41][0] <= 8'b0111_1111;					inform_R [42][0] <= 8'b0111_1111;					inform_R [43][0] <= 8'b0111_1111;					inform_R [44][0] <= 8'b0111_1111;					inform_R [45][0] <= 8'b0111_1111;					inform_R [46][0] <= 8'b0111_1111;					inform_R [47][0] <= 8'b0111_1111;					inform_R [48][0] <= 8'b0111_1111;					inform_R [49][0] <= 8'b0111_1111;					inform_R [50][0] <= 8'b0111_1111;					inform_R [51][0] <= 8'b0111_1111;					inform_R [52][0] <= 8'b0111_1111;					inform_R [53][0] <= 8'b0111_1111;					inform_R [54][0] <= 8'b0111_1111;					inform_R [55][0] <= 8'b0111_1111;					inform_R [56][0] <= 8'b0111_1111;					inform_R [57][0] <= 8'b0111_1111;					inform_R [58][0] <= 8'b0111_1111;					inform_R [59][0] <= 8'b0111_1111;					inform_R [60][0] <= 8'b0111_1111;					inform_R [61][0] <= 8'b0111_1111;					inform_R [62][0] <= 8'b0111_1111;					inform_R [63][0] <= 8'b0000_0000;					inform_R [64][0] <= 8'b0111_1111;					inform_R [65][0] <= 8'b0111_1111;					inform_R [66][0] <= 8'b0111_1111;					inform_R [67][0] <= 8'b0111_1111;					inform_R [68][0] <= 8'b0111_1111;					inform_R [69][0] <= 8'b0111_1111;					inform_R [70][0] <= 8'b0111_1111;					inform_R [71][0] <= 8'b0111_1111;					inform_R [72][0] <= 8'b0111_1111;					inform_R [73][0] <= 8'b0111_1111;					inform_R [74][0] <= 8'b0111_1111;					inform_R [75][0] <= 8'b0111_1111;					inform_R [76][0] <= 8'b0111_1111;					inform_R [77][0] <= 8'b0111_1111;					inform_R [78][0] <= 8'b0111_1111;					inform_R [79][0] <= 8'b0111_1111;					inform_R [80][0] <= 8'b0111_1111;					inform_R [81][0] <= 8'b0111_1111;					inform_R [82][0] <= 8'b0111_1111;					inform_R [83][0] <= 8'b0111_1111;					inform_R [84][0] <= 8'b0111_1111;					inform_R [85][0] <= 8'b0111_1111;					inform_R [86][0] <= 8'b0111_1111;					inform_R [87][0] <= 8'b0111_1111;					inform_R [88][0] <= 8'b0111_1111;					inform_R [89][0] <= 8'b0111_1111;					inform_R [90][0] <= 8'b0111_1111;					inform_R [91][0] <= 8'b0111_1111;					inform_R [92][0] <= 8'b0111_1111;					inform_R [93][0] <= 8'b0111_1111;					inform_R [94][0] <= 8'b0111_1111;					inform_R [95][0] <= 8'b0000_0000;					inform_R [96][0] <= 8'b0111_1111;					inform_R [97][0] <= 8'b0111_1111;					inform_R [98][0] <= 8'b0111_1111;					inform_R [99][0] <= 8'b0111_1111;					inform_R [100][0] <= 8'b0111_1111;					inform_R [101][0] <= 8'b0111_1111;					inform_R [102][0] <= 8'b0111_1111;					inform_R [103][0] <= 8'b0111_1111;					inform_R [104][0] <= 8'b0111_1111;					inform_R [105][0] <= 8'b0111_1111;					inform_R [106][0] <= 8'b0111_1111;					inform_R [107][0] <= 8'b0111_1111;					inform_R [108][0] <= 8'b0111_1111;					inform_R [109][0] <= 8'b0111_1111;					inform_R [110][0] <= 8'b0111_1111;					inform_R [111][0] <= 8'b0000_0000;					inform_R [112][0] <= 8'b0111_1111;					inform_R [113][0] <= 8'b0111_1111;					inform_R [114][0] <= 8'b0111_1111;					inform_R [115][0] <= 8'b0111_1111;					inform_R [116][0] <= 8'b0111_1111;					inform_R [117][0] <= 8'b0111_1111;					inform_R [118][0] <= 8'b0111_1111;					inform_R [119][0] <= 8'b0000_0000;					inform_R [120][0] <= 8'b0111_1111;					inform_R [121][0] <= 8'b0111_1111;					inform_R [122][0] <= 8'b0000_0000;					inform_R [123][0] <= 8'b0000_0000;					inform_R [124][0] <= 8'b0000_0000;					inform_R [125][0] <= 8'b0000_0000;					inform_R [126][0] <= 8'b0000_0000;					inform_R [127][0] <= 8'b0000_0000;					inform_R [128][0] <= 8'b0111_1111;					inform_R [129][0] <= 8'b0111_1111;					inform_R [130][0] <= 8'b0111_1111;					inform_R [131][0] <= 8'b0111_1111;					inform_R [132][0] <= 8'b0111_1111;					inform_R [133][0] <= 8'b0111_1111;					inform_R [134][0] <= 8'b0111_1111;					inform_R [135][0] <= 8'b0111_1111;					inform_R [136][0] <= 8'b0111_1111;					inform_R [137][0] <= 8'b0111_1111;					inform_R [138][0] <= 8'b0111_1111;					inform_R [139][0] <= 8'b0111_1111;					inform_R [140][0] <= 8'b0111_1111;					inform_R [141][0] <= 8'b0111_1111;					inform_R [142][0] <= 8'b0111_1111;					inform_R [143][0] <= 8'b0111_1111;					inform_R [144][0] <= 8'b0111_1111;					inform_R [145][0] <= 8'b0111_1111;					inform_R [146][0] <= 8'b0111_1111;					inform_R [147][0] <= 8'b0111_1111;					inform_R [148][0] <= 8'b0111_1111;					inform_R [149][0] <= 8'b0111_1111;					inform_R [150][0] <= 8'b0111_1111;					inform_R [151][0] <= 8'b0111_1111;					inform_R [152][0] <= 8'b0111_1111;					inform_R [153][0] <= 8'b0111_1111;					inform_R [154][0] <= 8'b0111_1111;					inform_R [155][0] <= 8'b0111_1111;					inform_R [156][0] <= 8'b0111_1111;					inform_R [157][0] <= 8'b0111_1111;					inform_R [158][0] <= 8'b0111_1111;					inform_R [159][0] <= 8'b0000_0000;					inform_R [160][0] <= 8'b0111_1111;					inform_R [161][0] <= 8'b0111_1111;					inform_R [162][0] <= 8'b0111_1111;					inform_R [163][0] <= 8'b0111_1111;					inform_R [164][0] <= 8'b0111_1111;					inform_R [165][0] <= 8'b0111_1111;					inform_R [166][0] <= 8'b0111_1111;					inform_R [167][0] <= 8'b0111_1111;					inform_R [168][0] <= 8'b0111_1111;					inform_R [169][0] <= 8'b0111_1111;					inform_R [170][0] <= 8'b0111_1111;					inform_R [171][0] <= 8'b0111_1111;					inform_R [172][0] <= 8'b0111_1111;					inform_R [173][0] <= 8'b0111_1111;					inform_R [174][0] <= 8'b0111_1111;					inform_R [175][0] <= 8'b0000_0000;					inform_R [176][0] <= 8'b0111_1111;					inform_R [177][0] <= 8'b0111_1111;					inform_R [178][0] <= 8'b0111_1111;					inform_R [179][0] <= 8'b0111_1111;					inform_R [180][0] <= 8'b0111_1111;					inform_R [181][0] <= 8'b0000_0000;					inform_R [182][0] <= 8'b0000_0000;					inform_R [183][0] <= 8'b0000_0000;					inform_R [184][0] <= 8'b0111_1111;					inform_R [185][0] <= 8'b0000_0000;					inform_R [186][0] <= 8'b0000_0000;					inform_R [187][0] <= 8'b0000_0000;					inform_R [188][0] <= 8'b0000_0000;					inform_R [189][0] <= 8'b0000_0000;					inform_R [190][0] <= 8'b0000_0000;					inform_R [191][0] <= 8'b0000_0000;					inform_R [192][0] <= 8'b0111_1111;					inform_R [193][0] <= 8'b0111_1111;					inform_R [194][0] <= 8'b0111_1111;					inform_R [195][0] <= 8'b0111_1111;					inform_R [196][0] <= 8'b0111_1111;					inform_R [197][0] <= 8'b0111_1111;					inform_R [198][0] <= 8'b0111_1111;					inform_R [199][0] <= 8'b0000_0000;					inform_R [200][0] <= 8'b0111_1111;					inform_R [201][0] <= 8'b0111_1111;					inform_R [202][0] <= 8'b0111_1111;					inform_R [203][0] <= 8'b0000_0000;					inform_R [204][0] <= 8'b0111_1111;					inform_R [205][0] <= 8'b0000_0000;					inform_R [206][0] <= 8'b0000_0000;					inform_R [207][0] <= 8'b0000_0000;					inform_R [208][0] <= 8'b0111_1111;					inform_R [209][0] <= 8'b0111_1111;					inform_R [210][0] <= 8'b0111_1111;					inform_R [211][0] <= 8'b0000_0000;					inform_R [212][0] <= 8'b0111_1111;					inform_R [213][0] <= 8'b0000_0000;					inform_R [214][0] <= 8'b0000_0000;					inform_R [215][0] <= 8'b0000_0000;					inform_R [216][0] <= 8'b0111_1111;					inform_R [217][0] <= 8'b0000_0000;					inform_R [218][0] <= 8'b0000_0000;					inform_R [219][0] <= 8'b0000_0000;					inform_R [220][0] <= 8'b0000_0000;					inform_R [221][0] <= 8'b0000_0000;					inform_R [222][0] <= 8'b0000_0000;					inform_R [223][0] <= 8'b0000_0000;					inform_R [224][0] <= 8'b0111_1111;					inform_R [225][0] <= 8'b0111_1111;					inform_R [226][0] <= 8'b0111_1111;					inform_R [227][0] <= 8'b0000_0000;					inform_R [228][0] <= 8'b0111_1111;					inform_R [229][0] <= 8'b0000_0000;					inform_R [230][0] <= 8'b0000_0000;					inform_R [231][0] <= 8'b0000_0000;					inform_R [232][0] <= 8'b0000_0000;					inform_R [233][0] <= 8'b0000_0000;					inform_R [234][0] <= 8'b0000_0000;					inform_R [235][0] <= 8'b0000_0000;					inform_R [236][0] <= 8'b0000_0000;					inform_R [237][0] <= 8'b0000_0000;					inform_R [238][0] <= 8'b0000_0000;					inform_R [239][0] <= 8'b0000_0000;					inform_R [240][0] <= 8'b0000_0000;					inform_R [241][0] <= 8'b0000_0000;					inform_R [242][0] <= 8'b0000_0000;					inform_R [243][0] <= 8'b0000_0000;					inform_R [244][0] <= 8'b0000_0000;					inform_R [245][0] <= 8'b0000_0000;					inform_R [246][0] <= 8'b0000_0000;					inform_R [247][0] <= 8'b0000_0000;					inform_R [248][0] <= 8'b0000_0000;					inform_R [249][0] <= 8'b0000_0000;					inform_R [250][0] <= 8'b0000_0000;					inform_R [251][0] <= 8'b0000_0000;					inform_R [252][0] <= 8'b0000_0000;					inform_R [253][0] <= 8'b0000_0000;					inform_R [254][0] <= 8'b0000_0000;					inform_R [255][0] <= 8'b0000_0000;					inform_R [256][0] <= 8'b0111_1111;					inform_R [257][0] <= 8'b0111_1111;					inform_R [258][0] <= 8'b0111_1111;					inform_R [259][0] <= 8'b0111_1111;					inform_R [260][0] <= 8'b0111_1111;					inform_R [261][0] <= 8'b0111_1111;					inform_R [262][0] <= 8'b0111_1111;					inform_R [263][0] <= 8'b0111_1111;					inform_R [264][0] <= 8'b0111_1111;					inform_R [265][0] <= 8'b0111_1111;					inform_R [266][0] <= 8'b0111_1111;					inform_R [267][0] <= 8'b0111_1111;					inform_R [268][0] <= 8'b0111_1111;					inform_R [269][0] <= 8'b0111_1111;					inform_R [270][0] <= 8'b0111_1111;					inform_R [271][0] <= 8'b0111_1111;					inform_R [272][0] <= 8'b0111_1111;					inform_R [273][0] <= 8'b0111_1111;					inform_R [274][0] <= 8'b0111_1111;					inform_R [275][0] <= 8'b0111_1111;					inform_R [276][0] <= 8'b0111_1111;					inform_R [277][0] <= 8'b0111_1111;					inform_R [278][0] <= 8'b0111_1111;					inform_R [279][0] <= 8'b0000_0000;					inform_R [280][0] <= 8'b0111_1111;					inform_R [281][0] <= 8'b0111_1111;					inform_R [282][0] <= 8'b0111_1111;					inform_R [283][0] <= 8'b0000_0000;					inform_R [284][0] <= 8'b0111_1111;					inform_R [285][0] <= 8'b0000_0000;					inform_R [286][0] <= 8'b0000_0000;					inform_R [287][0] <= 8'b0000_0000;					inform_R [288][0] <= 8'b0111_1111;					inform_R [289][0] <= 8'b0111_1111;					inform_R [290][0] <= 8'b0111_1111;					inform_R [291][0] <= 8'b0111_1111;					inform_R [292][0] <= 8'b0111_1111;					inform_R [293][0] <= 8'b0111_1111;					inform_R [294][0] <= 8'b0111_1111;					inform_R [295][0] <= 8'b0000_0000;					inform_R [296][0] <= 8'b0111_1111;					inform_R [297][0] <= 8'b0111_1111;					inform_R [298][0] <= 8'b0111_1111;					inform_R [299][0] <= 8'b0000_0000;					inform_R [300][0] <= 8'b0111_1111;					inform_R [301][0] <= 8'b0000_0000;					inform_R [302][0] <= 8'b0000_0000;					inform_R [303][0] <= 8'b0000_0000;					inform_R [304][0] <= 8'b0111_1111;					inform_R [305][0] <= 8'b0111_1111;					inform_R [306][0] <= 8'b0111_1111;					inform_R [307][0] <= 8'b0000_0000;					inform_R [308][0] <= 8'b0111_1111;					inform_R [309][0] <= 8'b0000_0000;					inform_R [310][0] <= 8'b0000_0000;					inform_R [311][0] <= 8'b0000_0000;					inform_R [312][0] <= 8'b0111_1111;					inform_R [313][0] <= 8'b0000_0000;					inform_R [314][0] <= 8'b0000_0000;					inform_R [315][0] <= 8'b0000_0000;					inform_R [316][0] <= 8'b0000_0000;					inform_R [317][0] <= 8'b0000_0000;					inform_R [318][0] <= 8'b0000_0000;					inform_R [319][0] <= 8'b0000_0000;					inform_R [320][0] <= 8'b0111_1111;					inform_R [321][0] <= 8'b0111_1111;					inform_R [322][0] <= 8'b0111_1111;					inform_R [323][0] <= 8'b0111_1111;					inform_R [324][0] <= 8'b0111_1111;					inform_R [325][0] <= 8'b0111_1111;					inform_R [326][0] <= 8'b0111_1111;					inform_R [327][0] <= 8'b0000_0000;					inform_R [328][0] <= 8'b0111_1111;					inform_R [329][0] <= 8'b0111_1111;					inform_R [330][0] <= 8'b0111_1111;					inform_R [331][0] <= 8'b0000_0000;					inform_R [332][0] <= 8'b0111_1111;					inform_R [333][0] <= 8'b0000_0000;					inform_R [334][0] <= 8'b0000_0000;					inform_R [335][0] <= 8'b0000_0000;					inform_R [336][0] <= 8'b0111_1111;					inform_R [337][0] <= 8'b0111_1111;					inform_R [338][0] <= 8'b0111_1111;					inform_R [339][0] <= 8'b0000_0000;					inform_R [340][0] <= 8'b0000_0000;					inform_R [341][0] <= 8'b0000_0000;					inform_R [342][0] <= 8'b0000_0000;					inform_R [343][0] <= 8'b0000_0000;					inform_R [344][0] <= 8'b0000_0000;					inform_R [345][0] <= 8'b0000_0000;					inform_R [346][0] <= 8'b0000_0000;					inform_R [347][0] <= 8'b0000_0000;					inform_R [348][0] <= 8'b0000_0000;					inform_R [349][0] <= 8'b0000_0000;					inform_R [350][0] <= 8'b0000_0000;					inform_R [351][0] <= 8'b0000_0000;					inform_R [352][0] <= 8'b0111_1111;					inform_R [353][0] <= 8'b0000_0000;					inform_R [354][0] <= 8'b0000_0000;					inform_R [355][0] <= 8'b0000_0000;					inform_R [356][0] <= 8'b0000_0000;					inform_R [357][0] <= 8'b0000_0000;					inform_R [358][0] <= 8'b0000_0000;					inform_R [359][0] <= 8'b0000_0000;					inform_R [360][0] <= 8'b0000_0000;					inform_R [361][0] <= 8'b0000_0000;					inform_R [362][0] <= 8'b0000_0000;					inform_R [363][0] <= 8'b0000_0000;					inform_R [364][0] <= 8'b0000_0000;					inform_R [365][0] <= 8'b0000_0000;					inform_R [366][0] <= 8'b0000_0000;					inform_R [367][0] <= 8'b0000_0000;					inform_R [368][0] <= 8'b0000_0000;					inform_R [369][0] <= 8'b0000_0000;					inform_R [370][0] <= 8'b0000_0000;					inform_R [371][0] <= 8'b0000_0000;					inform_R [372][0] <= 8'b0000_0000;					inform_R [373][0] <= 8'b0000_0000;					inform_R [374][0] <= 8'b0000_0000;					inform_R [375][0] <= 8'b0000_0000;					inform_R [376][0] <= 8'b0000_0000;					inform_R [377][0] <= 8'b0000_0000;					inform_R [378][0] <= 8'b0000_0000;					inform_R [379][0] <= 8'b0000_0000;					inform_R [380][0] <= 8'b0000_0000;					inform_R [381][0] <= 8'b0000_0000;					inform_R [382][0] <= 8'b0000_0000;					inform_R [383][0] <= 8'b0000_0000;					inform_R [384][0] <= 8'b0111_1111;					inform_R [385][0] <= 8'b0111_1111;					inform_R [386][0] <= 8'b0111_1111;					inform_R [387][0] <= 8'b0111_1111;					inform_R [388][0] <= 8'b0111_1111;					inform_R [389][0] <= 8'b0111_1111;					inform_R [390][0] <= 8'b0000_0000;					inform_R [391][0] <= 8'b0000_0000;					inform_R [392][0] <= 8'b0111_1111;					inform_R [393][0] <= 8'b0000_0000;					inform_R [394][0] <= 8'b0000_0000;					inform_R [395][0] <= 8'b0000_0000;					inform_R [396][0] <= 8'b0000_0000;					inform_R [397][0] <= 8'b0000_0000;					inform_R [398][0] <= 8'b0000_0000;					inform_R [399][0] <= 8'b0000_0000;					inform_R [400][0] <= 8'b0111_1111;					inform_R [401][0] <= 8'b0000_0000;					inform_R [402][0] <= 8'b0000_0000;					inform_R [403][0] <= 8'b0000_0000;					inform_R [404][0] <= 8'b0000_0000;					inform_R [405][0] <= 8'b0000_0000;					inform_R [406][0] <= 8'b0000_0000;					inform_R [407][0] <= 8'b0000_0000;					inform_R [408][0] <= 8'b0000_0000;					inform_R [409][0] <= 8'b0000_0000;					inform_R [410][0] <= 8'b0000_0000;					inform_R [411][0] <= 8'b0000_0000;					inform_R [412][0] <= 8'b0000_0000;					inform_R [413][0] <= 8'b0000_0000;					inform_R [414][0] <= 8'b0000_0000;					inform_R [415][0] <= 8'b0000_0000;					inform_R [416][0] <= 8'b0111_1111;					inform_R [417][0] <= 8'b0000_0000;					inform_R [418][0] <= 8'b0000_0000;					inform_R [419][0] <= 8'b0000_0000;					inform_R [420][0] <= 8'b0000_0000;					inform_R [421][0] <= 8'b0000_0000;					inform_R [422][0] <= 8'b0000_0000;					inform_R [423][0] <= 8'b0000_0000;					inform_R [424][0] <= 8'b0000_0000;					inform_R [425][0] <= 8'b0000_0000;					inform_R [426][0] <= 8'b0000_0000;					inform_R [427][0] <= 8'b0000_0000;					inform_R [428][0] <= 8'b0000_0000;					inform_R [429][0] <= 8'b0000_0000;					inform_R [430][0] <= 8'b0000_0000;					inform_R [431][0] <= 8'b0000_0000;					inform_R [432][0] <= 8'b0000_0000;					inform_R [433][0] <= 8'b0000_0000;					inform_R [434][0] <= 8'b0000_0000;					inform_R [435][0] <= 8'b0000_0000;					inform_R [436][0] <= 8'b0000_0000;					inform_R [437][0] <= 8'b0000_0000;					inform_R [438][0] <= 8'b0000_0000;					inform_R [439][0] <= 8'b0000_0000;					inform_R [440][0] <= 8'b0000_0000;					inform_R [441][0] <= 8'b0000_0000;					inform_R [442][0] <= 8'b0000_0000;					inform_R [443][0] <= 8'b0000_0000;					inform_R [444][0] <= 8'b0000_0000;					inform_R [445][0] <= 8'b0000_0000;					inform_R [446][0] <= 8'b0000_0000;					inform_R [447][0] <= 8'b0000_0000;					inform_R [448][0] <= 8'b0000_0000;					inform_R [449][0] <= 8'b0000_0000;					inform_R [450][0] <= 8'b0000_0000;					inform_R [451][0] <= 8'b0000_0000;					inform_R [452][0] <= 8'b0000_0000;					inform_R [453][0] <= 8'b0000_0000;					inform_R [454][0] <= 8'b0000_0000;					inform_R [455][0] <= 8'b0000_0000;					inform_R [456][0] <= 8'b0000_0000;					inform_R [457][0] <= 8'b0000_0000;					inform_R [458][0] <= 8'b0000_0000;					inform_R [459][0] <= 8'b0000_0000;					inform_R [460][0] <= 8'b0000_0000;					inform_R [461][0] <= 8'b0000_0000;					inform_R [462][0] <= 8'b0000_0000;					inform_R [463][0] <= 8'b0000_0000;					inform_R [464][0] <= 8'b0000_0000;					inform_R [465][0] <= 8'b0000_0000;					inform_R [466][0] <= 8'b0000_0000;					inform_R [467][0] <= 8'b0000_0000;					inform_R [468][0] <= 8'b0000_0000;					inform_R [469][0] <= 8'b0000_0000;					inform_R [470][0] <= 8'b0000_0000;					inform_R [471][0] <= 8'b0000_0000;					inform_R [472][0] <= 8'b0000_0000;					inform_R [473][0] <= 8'b0000_0000;					inform_R [474][0] <= 8'b0000_0000;					inform_R [475][0] <= 8'b0000_0000;					inform_R [476][0] <= 8'b0000_0000;					inform_R [477][0] <= 8'b0000_0000;					inform_R [478][0] <= 8'b0000_0000;					inform_R [479][0] <= 8'b0000_0000;					inform_R [480][0] <= 8'b0000_0000;					inform_R [481][0] <= 8'b0000_0000;					inform_R [482][0] <= 8'b0000_0000;					inform_R [483][0] <= 8'b0000_0000;					inform_R [484][0] <= 8'b0000_0000;					inform_R [485][0] <= 8'b0000_0000;					inform_R [486][0] <= 8'b0000_0000;					inform_R [487][0] <= 8'b0000_0000;					inform_R [488][0] <= 8'b0000_0000;					inform_R [489][0] <= 8'b0000_0000;					inform_R [490][0] <= 8'b0000_0000;					inform_R [491][0] <= 8'b0000_0000;					inform_R [492][0] <= 8'b0000_0000;					inform_R [493][0] <= 8'b0000_0000;					inform_R [494][0] <= 8'b0000_0000;					inform_R [495][0] <= 8'b0000_0000;					inform_R [496][0] <= 8'b0000_0000;					inform_R [497][0] <= 8'b0000_0000;					inform_R [498][0] <= 8'b0000_0000;					inform_R [499][0] <= 8'b0000_0000;					inform_R [500][0] <= 8'b0000_0000;					inform_R [501][0] <= 8'b0000_0000;					inform_R [502][0] <= 8'b0000_0000;					inform_R [503][0] <= 8'b0000_0000;					inform_R [504][0] <= 8'b0000_0000;					inform_R [505][0] <= 8'b0000_0000;					inform_R [506][0] <= 8'b0000_0000;					inform_R [507][0] <= 8'b0000_0000;					inform_R [508][0] <= 8'b0000_0000;					inform_R [509][0] <= 8'b0000_0000;					inform_R [510][0] <= 8'b0000_0000;					inform_R [511][0] <= 8'b0000_0000;					inform_R [512][0] <= 8'b0111_1111;					inform_R [513][0] <= 8'b0111_1111;					inform_R [514][0] <= 8'b0111_1111;					inform_R [515][0] <= 8'b0111_1111;					inform_R [516][0] <= 8'b0111_1111;					inform_R [517][0] <= 8'b0111_1111;					inform_R [518][0] <= 8'b0111_1111;					inform_R [519][0] <= 8'b0111_1111;					inform_R [520][0] <= 8'b0111_1111;					inform_R [521][0] <= 8'b0111_1111;					inform_R [522][0] <= 8'b0111_1111;					inform_R [523][0] <= 8'b0111_1111;					inform_R [524][0] <= 8'b0111_1111;					inform_R [525][0] <= 8'b0111_1111;					inform_R [526][0] <= 8'b0111_1111;					inform_R [527][0] <= 8'b0000_0000;					inform_R [528][0] <= 8'b0111_1111;					inform_R [529][0] <= 8'b0111_1111;					inform_R [530][0] <= 8'b0111_1111;					inform_R [531][0] <= 8'b0111_1111;					inform_R [532][0] <= 8'b0111_1111;					inform_R [533][0] <= 8'b0111_1111;					inform_R [534][0] <= 8'b0111_1111;					inform_R [535][0] <= 8'b0000_0000;					inform_R [536][0] <= 8'b0111_1111;					inform_R [537][0] <= 8'b0111_1111;					inform_R [538][0] <= 8'b0111_1111;					inform_R [539][0] <= 8'b0000_0000;					inform_R [540][0] <= 8'b0111_1111;					inform_R [541][0] <= 8'b0000_0000;					inform_R [542][0] <= 8'b0000_0000;					inform_R [543][0] <= 8'b0000_0000;					inform_R [544][0] <= 8'b0111_1111;					inform_R [545][0] <= 8'b0111_1111;					inform_R [546][0] <= 8'b0111_1111;					inform_R [547][0] <= 8'b0111_1111;					inform_R [548][0] <= 8'b0111_1111;					inform_R [549][0] <= 8'b0111_1111;					inform_R [550][0] <= 8'b0111_1111;					inform_R [551][0] <= 8'b0000_0000;					inform_R [552][0] <= 8'b0111_1111;					inform_R [553][0] <= 8'b0111_1111;					inform_R [554][0] <= 8'b0000_0000;					inform_R [555][0] <= 8'b0000_0000;					inform_R [556][0] <= 8'b0000_0000;					inform_R [557][0] <= 8'b0000_0000;					inform_R [558][0] <= 8'b0000_0000;					inform_R [559][0] <= 8'b0000_0000;					inform_R [560][0] <= 8'b0111_1111;					inform_R [561][0] <= 8'b0000_0000;					inform_R [562][0] <= 8'b0000_0000;					inform_R [563][0] <= 8'b0000_0000;					inform_R [564][0] <= 8'b0000_0000;					inform_R [565][0] <= 8'b0000_0000;					inform_R [566][0] <= 8'b0000_0000;					inform_R [567][0] <= 8'b0000_0000;					inform_R [568][0] <= 8'b0000_0000;					inform_R [569][0] <= 8'b0000_0000;					inform_R [570][0] <= 8'b0000_0000;					inform_R [571][0] <= 8'b0000_0000;					inform_R [572][0] <= 8'b0000_0000;					inform_R [573][0] <= 8'b0000_0000;					inform_R [574][0] <= 8'b0000_0000;					inform_R [575][0] <= 8'b0000_0000;					inform_R [576][0] <= 8'b0111_1111;					inform_R [577][0] <= 8'b0111_1111;					inform_R [578][0] <= 8'b0111_1111;					inform_R [579][0] <= 8'b0000_0000;					inform_R [580][0] <= 8'b0111_1111;					inform_R [581][0] <= 8'b0000_0000;					inform_R [582][0] <= 8'b0000_0000;					inform_R [583][0] <= 8'b0000_0000;					inform_R [584][0] <= 8'b0111_1111;					inform_R [585][0] <= 8'b0000_0000;					inform_R [586][0] <= 8'b0000_0000;					inform_R [587][0] <= 8'b0000_0000;					inform_R [588][0] <= 8'b0000_0000;					inform_R [589][0] <= 8'b0000_0000;					inform_R [590][0] <= 8'b0000_0000;					inform_R [591][0] <= 8'b0000_0000;					inform_R [592][0] <= 8'b0111_1111;					inform_R [593][0] <= 8'b0000_0000;					inform_R [594][0] <= 8'b0000_0000;					inform_R [595][0] <= 8'b0000_0000;					inform_R [596][0] <= 8'b0000_0000;					inform_R [597][0] <= 8'b0000_0000;					inform_R [598][0] <= 8'b0000_0000;					inform_R [599][0] <= 8'b0000_0000;					inform_R [600][0] <= 8'b0000_0000;					inform_R [601][0] <= 8'b0000_0000;					inform_R [602][0] <= 8'b0000_0000;					inform_R [603][0] <= 8'b0000_0000;					inform_R [604][0] <= 8'b0000_0000;					inform_R [605][0] <= 8'b0000_0000;					inform_R [606][0] <= 8'b0000_0000;					inform_R [607][0] <= 8'b0000_0000;					inform_R [608][0] <= 8'b0000_0000;					inform_R [609][0] <= 8'b0000_0000;					inform_R [610][0] <= 8'b0000_0000;					inform_R [611][0] <= 8'b0000_0000;					inform_R [612][0] <= 8'b0000_0000;					inform_R [613][0] <= 8'b0000_0000;					inform_R [614][0] <= 8'b0000_0000;					inform_R [615][0] <= 8'b0000_0000;					inform_R [616][0] <= 8'b0000_0000;					inform_R [617][0] <= 8'b0000_0000;					inform_R [618][0] <= 8'b0000_0000;					inform_R [619][0] <= 8'b0000_0000;					inform_R [620][0] <= 8'b0000_0000;					inform_R [621][0] <= 8'b0000_0000;					inform_R [622][0] <= 8'b0000_0000;					inform_R [623][0] <= 8'b0000_0000;					inform_R [624][0] <= 8'b0000_0000;					inform_R [625][0] <= 8'b0000_0000;					inform_R [626][0] <= 8'b0000_0000;					inform_R [627][0] <= 8'b0000_0000;					inform_R [628][0] <= 8'b0000_0000;					inform_R [629][0] <= 8'b0000_0000;					inform_R [630][0] <= 8'b0000_0000;					inform_R [631][0] <= 8'b0000_0000;					inform_R [632][0] <= 8'b0000_0000;					inform_R [633][0] <= 8'b0000_0000;					inform_R [634][0] <= 8'b0000_0000;					inform_R [635][0] <= 8'b0000_0000;					inform_R [636][0] <= 8'b0000_0000;					inform_R [637][0] <= 8'b0000_0000;					inform_R [638][0] <= 8'b0000_0000;					inform_R [639][0] <= 8'b0000_0000;					inform_R [640][0] <= 8'b0111_1111;					inform_R [641][0] <= 8'b0111_1111;					inform_R [642][0] <= 8'b0111_1111;					inform_R [643][0] <= 8'b0000_0000;					inform_R [644][0] <= 8'b0111_1111;					inform_R [645][0] <= 8'b0000_0000;					inform_R [646][0] <= 8'b0000_0000;					inform_R [647][0] <= 8'b0000_0000;					inform_R [648][0] <= 8'b0000_0000;					inform_R [649][0] <= 8'b0000_0000;					inform_R [650][0] <= 8'b0000_0000;					inform_R [651][0] <= 8'b0000_0000;					inform_R [652][0] <= 8'b0000_0000;					inform_R [653][0] <= 8'b0000_0000;					inform_R [654][0] <= 8'b0000_0000;					inform_R [655][0] <= 8'b0000_0000;					inform_R [656][0] <= 8'b0000_0000;					inform_R [657][0] <= 8'b0000_0000;					inform_R [658][0] <= 8'b0000_0000;					inform_R [659][0] <= 8'b0000_0000;					inform_R [660][0] <= 8'b0000_0000;					inform_R [661][0] <= 8'b0000_0000;					inform_R [662][0] <= 8'b0000_0000;					inform_R [663][0] <= 8'b0000_0000;					inform_R [664][0] <= 8'b0000_0000;					inform_R [665][0] <= 8'b0000_0000;					inform_R [666][0] <= 8'b0000_0000;					inform_R [667][0] <= 8'b0000_0000;					inform_R [668][0] <= 8'b0000_0000;					inform_R [669][0] <= 8'b0000_0000;					inform_R [670][0] <= 8'b0000_0000;					inform_R [671][0] <= 8'b0000_0000;					inform_R [672][0] <= 8'b0000_0000;					inform_R [673][0] <= 8'b0000_0000;					inform_R [674][0] <= 8'b0000_0000;					inform_R [675][0] <= 8'b0000_0000;					inform_R [676][0] <= 8'b0000_0000;					inform_R [677][0] <= 8'b0000_0000;					inform_R [678][0] <= 8'b0000_0000;					inform_R [679][0] <= 8'b0000_0000;					inform_R [680][0] <= 8'b0000_0000;					inform_R [681][0] <= 8'b0000_0000;					inform_R [682][0] <= 8'b0000_0000;					inform_R [683][0] <= 8'b0000_0000;					inform_R [684][0] <= 8'b0000_0000;					inform_R [685][0] <= 8'b0000_0000;					inform_R [686][0] <= 8'b0000_0000;					inform_R [687][0] <= 8'b0000_0000;					inform_R [688][0] <= 8'b0000_0000;					inform_R [689][0] <= 8'b0000_0000;					inform_R [690][0] <= 8'b0000_0000;					inform_R [691][0] <= 8'b0000_0000;					inform_R [692][0] <= 8'b0000_0000;					inform_R [693][0] <= 8'b0000_0000;					inform_R [694][0] <= 8'b0000_0000;					inform_R [695][0] <= 8'b0000_0000;					inform_R [696][0] <= 8'b0000_0000;					inform_R [697][0] <= 8'b0000_0000;					inform_R [698][0] <= 8'b0000_0000;					inform_R [699][0] <= 8'b0000_0000;					inform_R [700][0] <= 8'b0000_0000;					inform_R [701][0] <= 8'b0000_0000;					inform_R [702][0] <= 8'b0000_0000;					inform_R [703][0] <= 8'b0000_0000;					inform_R [704][0] <= 8'b0000_0000;					inform_R [705][0] <= 8'b0000_0000;					inform_R [706][0] <= 8'b0000_0000;					inform_R [707][0] <= 8'b0000_0000;					inform_R [708][0] <= 8'b0000_0000;					inform_R [709][0] <= 8'b0000_0000;					inform_R [710][0] <= 8'b0000_0000;					inform_R [711][0] <= 8'b0000_0000;					inform_R [712][0] <= 8'b0000_0000;					inform_R [713][0] <= 8'b0000_0000;					inform_R [714][0] <= 8'b0000_0000;					inform_R [715][0] <= 8'b0000_0000;					inform_R [716][0] <= 8'b0000_0000;					inform_R [717][0] <= 8'b0000_0000;					inform_R [718][0] <= 8'b0000_0000;					inform_R [719][0] <= 8'b0000_0000;					inform_R [720][0] <= 8'b0000_0000;					inform_R [721][0] <= 8'b0000_0000;					inform_R [722][0] <= 8'b0000_0000;					inform_R [723][0] <= 8'b0000_0000;					inform_R [724][0] <= 8'b0000_0000;					inform_R [725][0] <= 8'b0000_0000;					inform_R [726][0] <= 8'b0000_0000;					inform_R [727][0] <= 8'b0000_0000;					inform_R [728][0] <= 8'b0000_0000;					inform_R [729][0] <= 8'b0000_0000;					inform_R [730][0] <= 8'b0000_0000;					inform_R [731][0] <= 8'b0000_0000;					inform_R [732][0] <= 8'b0000_0000;					inform_R [733][0] <= 8'b0000_0000;					inform_R [734][0] <= 8'b0000_0000;					inform_R [735][0] <= 8'b0000_0000;					inform_R [736][0] <= 8'b0000_0000;					inform_R [737][0] <= 8'b0000_0000;					inform_R [738][0] <= 8'b0000_0000;					inform_R [739][0] <= 8'b0000_0000;					inform_R [740][0] <= 8'b0000_0000;					inform_R [741][0] <= 8'b0000_0000;					inform_R [742][0] <= 8'b0000_0000;					inform_R [743][0] <= 8'b0000_0000;					inform_R [744][0] <= 8'b0000_0000;					inform_R [745][0] <= 8'b0000_0000;					inform_R [746][0] <= 8'b0000_0000;					inform_R [747][0] <= 8'b0000_0000;					inform_R [748][0] <= 8'b0000_0000;					inform_R [749][0] <= 8'b0000_0000;					inform_R [750][0] <= 8'b0000_0000;					inform_R [751][0] <= 8'b0000_0000;					inform_R [752][0] <= 8'b0000_0000;					inform_R [753][0] <= 8'b0000_0000;					inform_R [754][0] <= 8'b0000_0000;					inform_R [755][0] <= 8'b0000_0000;					inform_R [756][0] <= 8'b0000_0000;					inform_R [757][0] <= 8'b0000_0000;					inform_R [758][0] <= 8'b0000_0000;					inform_R [759][0] <= 8'b0000_0000;					inform_R [760][0] <= 8'b0000_0000;					inform_R [761][0] <= 8'b0000_0000;					inform_R [762][0] <= 8'b0000_0000;					inform_R [763][0] <= 8'b0000_0000;					inform_R [764][0] <= 8'b0000_0000;					inform_R [765][0] <= 8'b0000_0000;					inform_R [766][0] <= 8'b0000_0000;					inform_R [767][0] <= 8'b0000_0000;					inform_R [768][0] <= 8'b0111_1111;					inform_R [769][0] <= 8'b0000_0000;					inform_R [770][0] <= 8'b0000_0000;					inform_R [771][0] <= 8'b0000_0000;					inform_R [772][0] <= 8'b0000_0000;					inform_R [773][0] <= 8'b0000_0000;					inform_R [774][0] <= 8'b0000_0000;					inform_R [775][0] <= 8'b0000_0000;					inform_R [776][0] <= 8'b0000_0000;					inform_R [777][0] <= 8'b0000_0000;					inform_R [778][0] <= 8'b0000_0000;					inform_R [779][0] <= 8'b0000_0000;					inform_R [780][0] <= 8'b0000_0000;					inform_R [781][0] <= 8'b0000_0000;					inform_R [782][0] <= 8'b0000_0000;					inform_R [783][0] <= 8'b0000_0000;					inform_R [784][0] <= 8'b0000_0000;					inform_R [785][0] <= 8'b0000_0000;					inform_R [786][0] <= 8'b0000_0000;					inform_R [787][0] <= 8'b0000_0000;					inform_R [788][0] <= 8'b0000_0000;					inform_R [789][0] <= 8'b0000_0000;					inform_R [790][0] <= 8'b0000_0000;					inform_R [791][0] <= 8'b0000_0000;					inform_R [792][0] <= 8'b0000_0000;					inform_R [793][0] <= 8'b0000_0000;					inform_R [794][0] <= 8'b0000_0000;					inform_R [795][0] <= 8'b0000_0000;					inform_R [796][0] <= 8'b0000_0000;					inform_R [797][0] <= 8'b0000_0000;					inform_R [798][0] <= 8'b0000_0000;					inform_R [799][0] <= 8'b0000_0000;					inform_R [800][0] <= 8'b0000_0000;					inform_R [801][0] <= 8'b0000_0000;					inform_R [802][0] <= 8'b0000_0000;					inform_R [803][0] <= 8'b0000_0000;					inform_R [804][0] <= 8'b0000_0000;					inform_R [805][0] <= 8'b0000_0000;					inform_R [806][0] <= 8'b0000_0000;					inform_R [807][0] <= 8'b0000_0000;					inform_R [808][0] <= 8'b0000_0000;					inform_R [809][0] <= 8'b0000_0000;					inform_R [810][0] <= 8'b0000_0000;					inform_R [811][0] <= 8'b0000_0000;					inform_R [812][0] <= 8'b0000_0000;					inform_R [813][0] <= 8'b0000_0000;					inform_R [814][0] <= 8'b0000_0000;					inform_R [815][0] <= 8'b0000_0000;					inform_R [816][0] <= 8'b0000_0000;					inform_R [817][0] <= 8'b0000_0000;					inform_R [818][0] <= 8'b0000_0000;					inform_R [819][0] <= 8'b0000_0000;					inform_R [820][0] <= 8'b0000_0000;					inform_R [821][0] <= 8'b0000_0000;					inform_R [822][0] <= 8'b0000_0000;					inform_R [823][0] <= 8'b0000_0000;					inform_R [824][0] <= 8'b0000_0000;					inform_R [825][0] <= 8'b0000_0000;					inform_R [826][0] <= 8'b0000_0000;					inform_R [827][0] <= 8'b0000_0000;					inform_R [828][0] <= 8'b0000_0000;					inform_R [829][0] <= 8'b0000_0000;					inform_R [830][0] <= 8'b0000_0000;					inform_R [831][0] <= 8'b0000_0000;					inform_R [832][0] <= 8'b0000_0000;					inform_R [833][0] <= 8'b0000_0000;					inform_R [834][0] <= 8'b0000_0000;					inform_R [835][0] <= 8'b0000_0000;					inform_R [836][0] <= 8'b0000_0000;					inform_R [837][0] <= 8'b0000_0000;					inform_R [838][0] <= 8'b0000_0000;					inform_R [839][0] <= 8'b0000_0000;					inform_R [840][0] <= 8'b0000_0000;					inform_R [841][0] <= 8'b0000_0000;					inform_R [842][0] <= 8'b0000_0000;					inform_R [843][0] <= 8'b0000_0000;					inform_R [844][0] <= 8'b0000_0000;					inform_R [845][0] <= 8'b0000_0000;					inform_R [846][0] <= 8'b0000_0000;					inform_R [847][0] <= 8'b0000_0000;					inform_R [848][0] <= 8'b0000_0000;					inform_R [849][0] <= 8'b0000_0000;					inform_R [850][0] <= 8'b0000_0000;					inform_R [851][0] <= 8'b0000_0000;					inform_R [852][0] <= 8'b0000_0000;					inform_R [853][0] <= 8'b0000_0000;					inform_R [854][0] <= 8'b0000_0000;					inform_R [855][0] <= 8'b0000_0000;					inform_R [856][0] <= 8'b0000_0000;					inform_R [857][0] <= 8'b0000_0000;					inform_R [858][0] <= 8'b0000_0000;					inform_R [859][0] <= 8'b0000_0000;					inform_R [860][0] <= 8'b0000_0000;					inform_R [861][0] <= 8'b0000_0000;					inform_R [862][0] <= 8'b0000_0000;					inform_R [863][0] <= 8'b0000_0000;					inform_R [864][0] <= 8'b0000_0000;					inform_R [865][0] <= 8'b0000_0000;					inform_R [866][0] <= 8'b0000_0000;					inform_R [867][0] <= 8'b0000_0000;					inform_R [868][0] <= 8'b0000_0000;					inform_R [869][0] <= 8'b0000_0000;					inform_R [870][0] <= 8'b0000_0000;					inform_R [871][0] <= 8'b0000_0000;					inform_R [872][0] <= 8'b0000_0000;					inform_R [873][0] <= 8'b0000_0000;					inform_R [874][0] <= 8'b0000_0000;					inform_R [875][0] <= 8'b0000_0000;					inform_R [876][0] <= 8'b0000_0000;					inform_R [877][0] <= 8'b0000_0000;					inform_R [878][0] <= 8'b0000_0000;					inform_R [879][0] <= 8'b0000_0000;					inform_R [880][0] <= 8'b0000_0000;					inform_R [881][0] <= 8'b0000_0000;					inform_R [882][0] <= 8'b0000_0000;					inform_R [883][0] <= 8'b0000_0000;					inform_R [884][0] <= 8'b0000_0000;					inform_R [885][0] <= 8'b0000_0000;					inform_R [886][0] <= 8'b0000_0000;					inform_R [887][0] <= 8'b0000_0000;					inform_R [888][0] <= 8'b0000_0000;					inform_R [889][0] <= 8'b0000_0000;					inform_R [890][0] <= 8'b0000_0000;					inform_R [891][0] <= 8'b0000_0000;					inform_R [892][0] <= 8'b0000_0000;					inform_R [893][0] <= 8'b0000_0000;					inform_R [894][0] <= 8'b0000_0000;					inform_R [895][0] <= 8'b0000_0000;					inform_R [896][0] <= 8'b0000_0000;					inform_R [897][0] <= 8'b0000_0000;					inform_R [898][0] <= 8'b0000_0000;					inform_R [899][0] <= 8'b0000_0000;					inform_R [900][0] <= 8'b0000_0000;					inform_R [901][0] <= 8'b0000_0000;					inform_R [902][0] <= 8'b0000_0000;					inform_R [903][0] <= 8'b0000_0000;					inform_R [904][0] <= 8'b0000_0000;					inform_R [905][0] <= 8'b0000_0000;					inform_R [906][0] <= 8'b0000_0000;					inform_R [907][0] <= 8'b0000_0000;					inform_R [908][0] <= 8'b0000_0000;					inform_R [909][0] <= 8'b0000_0000;					inform_R [910][0] <= 8'b0000_0000;					inform_R [911][0] <= 8'b0000_0000;					inform_R [912][0] <= 8'b0000_0000;					inform_R [913][0] <= 8'b0000_0000;					inform_R [914][0] <= 8'b0000_0000;					inform_R [915][0] <= 8'b0000_0000;					inform_R [916][0] <= 8'b0000_0000;					inform_R [917][0] <= 8'b0000_0000;					inform_R [918][0] <= 8'b0000_0000;					inform_R [919][0] <= 8'b0000_0000;					inform_R [920][0] <= 8'b0000_0000;					inform_R [921][0] <= 8'b0000_0000;					inform_R [922][0] <= 8'b0000_0000;					inform_R [923][0] <= 8'b0000_0000;					inform_R [924][0] <= 8'b0000_0000;					inform_R [925][0] <= 8'b0000_0000;					inform_R [926][0] <= 8'b0000_0000;					inform_R [927][0] <= 8'b0000_0000;					inform_R [928][0] <= 8'b0000_0000;					inform_R [929][0] <= 8'b0000_0000;					inform_R [930][0] <= 8'b0000_0000;					inform_R [931][0] <= 8'b0000_0000;					inform_R [932][0] <= 8'b0000_0000;					inform_R [933][0] <= 8'b0000_0000;					inform_R [934][0] <= 8'b0000_0000;					inform_R [935][0] <= 8'b0000_0000;					inform_R [936][0] <= 8'b0000_0000;					inform_R [937][0] <= 8'b0000_0000;					inform_R [938][0] <= 8'b0000_0000;					inform_R [939][0] <= 8'b0000_0000;					inform_R [940][0] <= 8'b0000_0000;					inform_R [941][0] <= 8'b0000_0000;					inform_R [942][0] <= 8'b0000_0000;					inform_R [943][0] <= 8'b0000_0000;					inform_R [944][0] <= 8'b0000_0000;					inform_R [945][0] <= 8'b0000_0000;					inform_R [946][0] <= 8'b0000_0000;					inform_R [947][0] <= 8'b0000_0000;					inform_R [948][0] <= 8'b0000_0000;					inform_R [949][0] <= 8'b0000_0000;					inform_R [950][0] <= 8'b0000_0000;					inform_R [951][0] <= 8'b0000_0000;					inform_R [952][0] <= 8'b0000_0000;					inform_R [953][0] <= 8'b0000_0000;					inform_R [954][0] <= 8'b0000_0000;					inform_R [955][0] <= 8'b0000_0000;					inform_R [956][0] <= 8'b0000_0000;					inform_R [957][0] <= 8'b0000_0000;					inform_R [958][0] <= 8'b0000_0000;					inform_R [959][0] <= 8'b0000_0000;					inform_R [960][0] <= 8'b0000_0000;					inform_R [961][0] <= 8'b0000_0000;					inform_R [962][0] <= 8'b0000_0000;					inform_R [963][0] <= 8'b0000_0000;					inform_R [964][0] <= 8'b0000_0000;					inform_R [965][0] <= 8'b0000_0000;					inform_R [966][0] <= 8'b0000_0000;					inform_R [967][0] <= 8'b0000_0000;					inform_R [968][0] <= 8'b0000_0000;					inform_R [969][0] <= 8'b0000_0000;					inform_R [970][0] <= 8'b0000_0000;					inform_R [971][0] <= 8'b0000_0000;					inform_R [972][0] <= 8'b0000_0000;					inform_R [973][0] <= 8'b0000_0000;					inform_R [974][0] <= 8'b0000_0000;					inform_R [975][0] <= 8'b0000_0000;					inform_R [976][0] <= 8'b0000_0000;					inform_R [977][0] <= 8'b0000_0000;					inform_R [978][0] <= 8'b0000_0000;					inform_R [979][0] <= 8'b0000_0000;					inform_R [980][0] <= 8'b0000_0000;					inform_R [981][0] <= 8'b0000_0000;					inform_R [982][0] <= 8'b0000_0000;					inform_R [983][0] <= 8'b0000_0000;					inform_R [984][0] <= 8'b0000_0000;					inform_R [985][0] <= 8'b0000_0000;					inform_R [986][0] <= 8'b0000_0000;					inform_R [987][0] <= 8'b0000_0000;					inform_R [988][0] <= 8'b0000_0000;					inform_R [989][0] <= 8'b0000_0000;					inform_R [990][0] <= 8'b0000_0000;					inform_R [991][0] <= 8'b0000_0000;					inform_R [992][0] <= 8'b0000_0000;					inform_R [993][0] <= 8'b0000_0000;					inform_R [994][0] <= 8'b0000_0000;					inform_R [995][0] <= 8'b0000_0000;					inform_R [996][0] <= 8'b0000_0000;					inform_R [997][0] <= 8'b0000_0000;					inform_R [998][0] <= 8'b0000_0000;					inform_R [999][0] <= 8'b0000_0000;					inform_R [1000][0] <= 8'b0000_0000;					inform_R [1001][0] <= 8'b0000_0000;					inform_R [1002][0] <= 8'b0000_0000;					inform_R [1003][0] <= 8'b0000_0000;					inform_R [1004][0] <= 8'b0000_0000;					inform_R [1005][0] <= 8'b0000_0000;					inform_R [1006][0] <= 8'b0000_0000;					inform_R [1007][0] <= 8'b0000_0000;					inform_R [1008][0] <= 8'b0000_0000;					inform_R [1009][0] <= 8'b0000_0000;					inform_R [1010][0] <= 8'b0000_0000;					inform_R [1011][0] <= 8'b0000_0000;					inform_R [1012][0] <= 8'b0000_0000;					inform_R [1013][0] <= 8'b0000_0000;					inform_R [1014][0] <= 8'b0000_0000;					inform_R [1015][0] <= 8'b0000_0000;					inform_R [1016][0] <= 8'b0000_0000;					inform_R [1017][0] <= 8'b0000_0000;					inform_R [1018][0] <= 8'b0000_0000;					inform_R [1019][0] <= 8'b0000_0000;					inform_R [1020][0] <= 8'b0000_0000;					inform_R [1021][0] <= 8'b0000_0000;					inform_R [1022][0] <= 8'b0000_0000;					inform_R [1023][0] <= 8'b0000_0000;					inform_L [0][10] <= LLR_1;					inform_L [1][10] <= LLR_2;					inform_L [2][10] <= LLR_3;					inform_L [3][10] <= LLR_4;					inform_L [4][10] <= LLR_5;					inform_L [5][10] <= LLR_6;					inform_L [6][10] <= LLR_7;					inform_L [7][10] <= LLR_8;					inform_L [8][10] <= LLR_9;					inform_L [9][10] <= LLR_10;					inform_L [10][10] <= LLR_11;					inform_L [11][10] <= LLR_12;					inform_L [12][10] <= LLR_13;					inform_L [13][10] <= LLR_14;					inform_L [14][10] <= LLR_15;					inform_L [15][10] <= LLR_16;					inform_L [16][10] <= LLR_17;					inform_L [17][10] <= LLR_18;					inform_L [18][10] <= LLR_19;					inform_L [19][10] <= LLR_20;					inform_L [20][10] <= LLR_21;					inform_L [21][10] <= LLR_22;					inform_L [22][10] <= LLR_23;					inform_L [23][10] <= LLR_24;					inform_L [24][10] <= LLR_25;					inform_L [25][10] <= LLR_26;					inform_L [26][10] <= LLR_27;					inform_L [27][10] <= LLR_28;					inform_L [28][10] <= LLR_29;					inform_L [29][10] <= LLR_30;					inform_L [30][10] <= LLR_31;					inform_L [31][10] <= LLR_32;					inform_L [32][10] <= LLR_33;					inform_L [33][10] <= LLR_34;					inform_L [34][10] <= LLR_35;					inform_L [35][10] <= LLR_36;					inform_L [36][10] <= LLR_37;					inform_L [37][10] <= LLR_38;					inform_L [38][10] <= LLR_39;					inform_L [39][10] <= LLR_40;					inform_L [40][10] <= LLR_41;					inform_L [41][10] <= LLR_42;					inform_L [42][10] <= LLR_43;					inform_L [43][10] <= LLR_44;					inform_L [44][10] <= LLR_45;					inform_L [45][10] <= LLR_46;					inform_L [46][10] <= LLR_47;					inform_L [47][10] <= LLR_48;					inform_L [48][10] <= LLR_49;					inform_L [49][10] <= LLR_50;					inform_L [50][10] <= LLR_51;					inform_L [51][10] <= LLR_52;					inform_L [52][10] <= LLR_53;					inform_L [53][10] <= LLR_54;					inform_L [54][10] <= LLR_55;					inform_L [55][10] <= LLR_56;					inform_L [56][10] <= LLR_57;					inform_L [57][10] <= LLR_58;					inform_L [58][10] <= LLR_59;					inform_L [59][10] <= LLR_60;					inform_L [60][10] <= LLR_61;					inform_L [61][10] <= LLR_62;					inform_L [62][10] <= LLR_63;					inform_L [63][10] <= LLR_64;					inform_L [64][10] <= LLR_65;					inform_L [65][10] <= LLR_66;					inform_L [66][10] <= LLR_67;					inform_L [67][10] <= LLR_68;					inform_L [68][10] <= LLR_69;					inform_L [69][10] <= LLR_70;					inform_L [70][10] <= LLR_71;					inform_L [71][10] <= LLR_72;					inform_L [72][10] <= LLR_73;					inform_L [73][10] <= LLR_74;					inform_L [74][10] <= LLR_75;					inform_L [75][10] <= LLR_76;					inform_L [76][10] <= LLR_77;					inform_L [77][10] <= LLR_78;					inform_L [78][10] <= LLR_79;					inform_L [79][10] <= LLR_80;					inform_L [80][10] <= LLR_81;					inform_L [81][10] <= LLR_82;					inform_L [82][10] <= LLR_83;					inform_L [83][10] <= LLR_84;					inform_L [84][10] <= LLR_85;					inform_L [85][10] <= LLR_86;					inform_L [86][10] <= LLR_87;					inform_L [87][10] <= LLR_88;					inform_L [88][10] <= LLR_89;					inform_L [89][10] <= LLR_90;					inform_L [90][10] <= LLR_91;					inform_L [91][10] <= LLR_92;					inform_L [92][10] <= LLR_93;					inform_L [93][10] <= LLR_94;					inform_L [94][10] <= LLR_95;					inform_L [95][10] <= LLR_96;					inform_L [96][10] <= LLR_97;					inform_L [97][10] <= LLR_98;					inform_L [98][10] <= LLR_99;					inform_L [99][10] <= LLR_100;					inform_L [100][10] <= LLR_101;					inform_L [101][10] <= LLR_102;					inform_L [102][10] <= LLR_103;					inform_L [103][10] <= LLR_104;					inform_L [104][10] <= LLR_105;					inform_L [105][10] <= LLR_106;					inform_L [106][10] <= LLR_107;					inform_L [107][10] <= LLR_108;					inform_L [108][10] <= LLR_109;					inform_L [109][10] <= LLR_110;					inform_L [110][10] <= LLR_111;					inform_L [111][10] <= LLR_112;					inform_L [112][10] <= LLR_113;					inform_L [113][10] <= LLR_114;					inform_L [114][10] <= LLR_115;					inform_L [115][10] <= LLR_116;					inform_L [116][10] <= LLR_117;					inform_L [117][10] <= LLR_118;					inform_L [118][10] <= LLR_119;					inform_L [119][10] <= LLR_120;					inform_L [120][10] <= LLR_121;					inform_L [121][10] <= LLR_122;					inform_L [122][10] <= LLR_123;					inform_L [123][10] <= LLR_124;					inform_L [124][10] <= LLR_125;					inform_L [125][10] <= LLR_126;					inform_L [126][10] <= LLR_127;					inform_L [127][10] <= LLR_128;					inform_L [128][10] <= LLR_129;					inform_L [129][10] <= LLR_130;					inform_L [130][10] <= LLR_131;					inform_L [131][10] <= LLR_132;					inform_L [132][10] <= LLR_133;					inform_L [133][10] <= LLR_134;					inform_L [134][10] <= LLR_135;					inform_L [135][10] <= LLR_136;					inform_L [136][10] <= LLR_137;					inform_L [137][10] <= LLR_138;					inform_L [138][10] <= LLR_139;					inform_L [139][10] <= LLR_140;					inform_L [140][10] <= LLR_141;					inform_L [141][10] <= LLR_142;					inform_L [142][10] <= LLR_143;					inform_L [143][10] <= LLR_144;					inform_L [144][10] <= LLR_145;					inform_L [145][10] <= LLR_146;					inform_L [146][10] <= LLR_147;					inform_L [147][10] <= LLR_148;					inform_L [148][10] <= LLR_149;					inform_L [149][10] <= LLR_150;					inform_L [150][10] <= LLR_151;					inform_L [151][10] <= LLR_152;					inform_L [152][10] <= LLR_153;					inform_L [153][10] <= LLR_154;					inform_L [154][10] <= LLR_155;					inform_L [155][10] <= LLR_156;					inform_L [156][10] <= LLR_157;					inform_L [157][10] <= LLR_158;					inform_L [158][10] <= LLR_159;					inform_L [159][10] <= LLR_160;					inform_L [160][10] <= LLR_161;					inform_L [161][10] <= LLR_162;					inform_L [162][10] <= LLR_163;					inform_L [163][10] <= LLR_164;					inform_L [164][10] <= LLR_165;					inform_L [165][10] <= LLR_166;					inform_L [166][10] <= LLR_167;					inform_L [167][10] <= LLR_168;					inform_L [168][10] <= LLR_169;					inform_L [169][10] <= LLR_170;					inform_L [170][10] <= LLR_171;					inform_L [171][10] <= LLR_172;					inform_L [172][10] <= LLR_173;					inform_L [173][10] <= LLR_174;					inform_L [174][10] <= LLR_175;					inform_L [175][10] <= LLR_176;					inform_L [176][10] <= LLR_177;					inform_L [177][10] <= LLR_178;					inform_L [178][10] <= LLR_179;					inform_L [179][10] <= LLR_180;					inform_L [180][10] <= LLR_181;					inform_L [181][10] <= LLR_182;					inform_L [182][10] <= LLR_183;					inform_L [183][10] <= LLR_184;					inform_L [184][10] <= LLR_185;					inform_L [185][10] <= LLR_186;					inform_L [186][10] <= LLR_187;					inform_L [187][10] <= LLR_188;					inform_L [188][10] <= LLR_189;					inform_L [189][10] <= LLR_190;					inform_L [190][10] <= LLR_191;					inform_L [191][10] <= LLR_192;					inform_L [192][10] <= LLR_193;					inform_L [193][10] <= LLR_194;					inform_L [194][10] <= LLR_195;					inform_L [195][10] <= LLR_196;					inform_L [196][10] <= LLR_197;					inform_L [197][10] <= LLR_198;					inform_L [198][10] <= LLR_199;					inform_L [199][10] <= LLR_200;					inform_L [200][10] <= LLR_201;					inform_L [201][10] <= LLR_202;					inform_L [202][10] <= LLR_203;					inform_L [203][10] <= LLR_204;					inform_L [204][10] <= LLR_205;					inform_L [205][10] <= LLR_206;					inform_L [206][10] <= LLR_207;					inform_L [207][10] <= LLR_208;					inform_L [208][10] <= LLR_209;					inform_L [209][10] <= LLR_210;					inform_L [210][10] <= LLR_211;					inform_L [211][10] <= LLR_212;					inform_L [212][10] <= LLR_213;					inform_L [213][10] <= LLR_214;					inform_L [214][10] <= LLR_215;					inform_L [215][10] <= LLR_216;					inform_L [216][10] <= LLR_217;					inform_L [217][10] <= LLR_218;					inform_L [218][10] <= LLR_219;					inform_L [219][10] <= LLR_220;					inform_L [220][10] <= LLR_221;					inform_L [221][10] <= LLR_222;					inform_L [222][10] <= LLR_223;					inform_L [223][10] <= LLR_224;					inform_L [224][10] <= LLR_225;					inform_L [225][10] <= LLR_226;					inform_L [226][10] <= LLR_227;					inform_L [227][10] <= LLR_228;					inform_L [228][10] <= LLR_229;					inform_L [229][10] <= LLR_230;					inform_L [230][10] <= LLR_231;					inform_L [231][10] <= LLR_232;					inform_L [232][10] <= LLR_233;					inform_L [233][10] <= LLR_234;					inform_L [234][10] <= LLR_235;					inform_L [235][10] <= LLR_236;					inform_L [236][10] <= LLR_237;					inform_L [237][10] <= LLR_238;					inform_L [238][10] <= LLR_239;					inform_L [239][10] <= LLR_240;					inform_L [240][10] <= LLR_241;					inform_L [241][10] <= LLR_242;					inform_L [242][10] <= LLR_243;					inform_L [243][10] <= LLR_244;					inform_L [244][10] <= LLR_245;					inform_L [245][10] <= LLR_246;					inform_L [246][10] <= LLR_247;					inform_L [247][10] <= LLR_248;					inform_L [248][10] <= LLR_249;					inform_L [249][10] <= LLR_250;					inform_L [250][10] <= LLR_251;					inform_L [251][10] <= LLR_252;					inform_L [252][10] <= LLR_253;					inform_L [253][10] <= LLR_254;					inform_L [254][10] <= LLR_255;					inform_L [255][10] <= LLR_256;					inform_L [256][10] <= LLR_257;					inform_L [257][10] <= LLR_258;					inform_L [258][10] <= LLR_259;					inform_L [259][10] <= LLR_260;					inform_L [260][10] <= LLR_261;					inform_L [261][10] <= LLR_262;					inform_L [262][10] <= LLR_263;					inform_L [263][10] <= LLR_264;					inform_L [264][10] <= LLR_265;					inform_L [265][10] <= LLR_266;					inform_L [266][10] <= LLR_267;					inform_L [267][10] <= LLR_268;					inform_L [268][10] <= LLR_269;					inform_L [269][10] <= LLR_270;					inform_L [270][10] <= LLR_271;					inform_L [271][10] <= LLR_272;					inform_L [272][10] <= LLR_273;					inform_L [273][10] <= LLR_274;					inform_L [274][10] <= LLR_275;					inform_L [275][10] <= LLR_276;					inform_L [276][10] <= LLR_277;					inform_L [277][10] <= LLR_278;					inform_L [278][10] <= LLR_279;					inform_L [279][10] <= LLR_280;					inform_L [280][10] <= LLR_281;					inform_L [281][10] <= LLR_282;					inform_L [282][10] <= LLR_283;					inform_L [283][10] <= LLR_284;					inform_L [284][10] <= LLR_285;					inform_L [285][10] <= LLR_286;					inform_L [286][10] <= LLR_287;					inform_L [287][10] <= LLR_288;					inform_L [288][10] <= LLR_289;					inform_L [289][10] <= LLR_290;					inform_L [290][10] <= LLR_291;					inform_L [291][10] <= LLR_292;					inform_L [292][10] <= LLR_293;					inform_L [293][10] <= LLR_294;					inform_L [294][10] <= LLR_295;					inform_L [295][10] <= LLR_296;					inform_L [296][10] <= LLR_297;					inform_L [297][10] <= LLR_298;					inform_L [298][10] <= LLR_299;					inform_L [299][10] <= LLR_300;					inform_L [300][10] <= LLR_301;					inform_L [301][10] <= LLR_302;					inform_L [302][10] <= LLR_303;					inform_L [303][10] <= LLR_304;					inform_L [304][10] <= LLR_305;					inform_L [305][10] <= LLR_306;					inform_L [306][10] <= LLR_307;					inform_L [307][10] <= LLR_308;					inform_L [308][10] <= LLR_309;					inform_L [309][10] <= LLR_310;					inform_L [310][10] <= LLR_311;					inform_L [311][10] <= LLR_312;					inform_L [312][10] <= LLR_313;					inform_L [313][10] <= LLR_314;					inform_L [314][10] <= LLR_315;					inform_L [315][10] <= LLR_316;					inform_L [316][10] <= LLR_317;					inform_L [317][10] <= LLR_318;					inform_L [318][10] <= LLR_319;					inform_L [319][10] <= LLR_320;					inform_L [320][10] <= LLR_321;					inform_L [321][10] <= LLR_322;					inform_L [322][10] <= LLR_323;					inform_L [323][10] <= LLR_324;					inform_L [324][10] <= LLR_325;					inform_L [325][10] <= LLR_326;					inform_L [326][10] <= LLR_327;					inform_L [327][10] <= LLR_328;					inform_L [328][10] <= LLR_329;					inform_L [329][10] <= LLR_330;					inform_L [330][10] <= LLR_331;					inform_L [331][10] <= LLR_332;					inform_L [332][10] <= LLR_333;					inform_L [333][10] <= LLR_334;					inform_L [334][10] <= LLR_335;					inform_L [335][10] <= LLR_336;					inform_L [336][10] <= LLR_337;					inform_L [337][10] <= LLR_338;					inform_L [338][10] <= LLR_339;					inform_L [339][10] <= LLR_340;					inform_L [340][10] <= LLR_341;					inform_L [341][10] <= LLR_342;					inform_L [342][10] <= LLR_343;					inform_L [343][10] <= LLR_344;					inform_L [344][10] <= LLR_345;					inform_L [345][10] <= LLR_346;					inform_L [346][10] <= LLR_347;					inform_L [347][10] <= LLR_348;					inform_L [348][10] <= LLR_349;					inform_L [349][10] <= LLR_350;					inform_L [350][10] <= LLR_351;					inform_L [351][10] <= LLR_352;					inform_L [352][10] <= LLR_353;					inform_L [353][10] <= LLR_354;					inform_L [354][10] <= LLR_355;					inform_L [355][10] <= LLR_356;					inform_L [356][10] <= LLR_357;					inform_L [357][10] <= LLR_358;					inform_L [358][10] <= LLR_359;					inform_L [359][10] <= LLR_360;					inform_L [360][10] <= LLR_361;					inform_L [361][10] <= LLR_362;					inform_L [362][10] <= LLR_363;					inform_L [363][10] <= LLR_364;					inform_L [364][10] <= LLR_365;					inform_L [365][10] <= LLR_366;					inform_L [366][10] <= LLR_367;					inform_L [367][10] <= LLR_368;					inform_L [368][10] <= LLR_369;					inform_L [369][10] <= LLR_370;					inform_L [370][10] <= LLR_371;					inform_L [371][10] <= LLR_372;					inform_L [372][10] <= LLR_373;					inform_L [373][10] <= LLR_374;					inform_L [374][10] <= LLR_375;					inform_L [375][10] <= LLR_376;					inform_L [376][10] <= LLR_377;					inform_L [377][10] <= LLR_378;					inform_L [378][10] <= LLR_379;					inform_L [379][10] <= LLR_380;					inform_L [380][10] <= LLR_381;					inform_L [381][10] <= LLR_382;					inform_L [382][10] <= LLR_383;					inform_L [383][10] <= LLR_384;					inform_L [384][10] <= LLR_385;					inform_L [385][10] <= LLR_386;					inform_L [386][10] <= LLR_387;					inform_L [387][10] <= LLR_388;					inform_L [388][10] <= LLR_389;					inform_L [389][10] <= LLR_390;					inform_L [390][10] <= LLR_391;					inform_L [391][10] <= LLR_392;					inform_L [392][10] <= LLR_393;					inform_L [393][10] <= LLR_394;					inform_L [394][10] <= LLR_395;					inform_L [395][10] <= LLR_396;					inform_L [396][10] <= LLR_397;					inform_L [397][10] <= LLR_398;					inform_L [398][10] <= LLR_399;					inform_L [399][10] <= LLR_400;					inform_L [400][10] <= LLR_401;					inform_L [401][10] <= LLR_402;					inform_L [402][10] <= LLR_403;					inform_L [403][10] <= LLR_404;					inform_L [404][10] <= LLR_405;					inform_L [405][10] <= LLR_406;					inform_L [406][10] <= LLR_407;					inform_L [407][10] <= LLR_408;					inform_L [408][10] <= LLR_409;					inform_L [409][10] <= LLR_410;					inform_L [410][10] <= LLR_411;					inform_L [411][10] <= LLR_412;					inform_L [412][10] <= LLR_413;					inform_L [413][10] <= LLR_414;					inform_L [414][10] <= LLR_415;					inform_L [415][10] <= LLR_416;					inform_L [416][10] <= LLR_417;					inform_L [417][10] <= LLR_418;					inform_L [418][10] <= LLR_419;					inform_L [419][10] <= LLR_420;					inform_L [420][10] <= LLR_421;					inform_L [421][10] <= LLR_422;					inform_L [422][10] <= LLR_423;					inform_L [423][10] <= LLR_424;					inform_L [424][10] <= LLR_425;					inform_L [425][10] <= LLR_426;					inform_L [426][10] <= LLR_427;					inform_L [427][10] <= LLR_428;					inform_L [428][10] <= LLR_429;					inform_L [429][10] <= LLR_430;					inform_L [430][10] <= LLR_431;					inform_L [431][10] <= LLR_432;					inform_L [432][10] <= LLR_433;					inform_L [433][10] <= LLR_434;					inform_L [434][10] <= LLR_435;					inform_L [435][10] <= LLR_436;					inform_L [436][10] <= LLR_437;					inform_L [437][10] <= LLR_438;					inform_L [438][10] <= LLR_439;					inform_L [439][10] <= LLR_440;					inform_L [440][10] <= LLR_441;					inform_L [441][10] <= LLR_442;					inform_L [442][10] <= LLR_443;					inform_L [443][10] <= LLR_444;					inform_L [444][10] <= LLR_445;					inform_L [445][10] <= LLR_446;					inform_L [446][10] <= LLR_447;					inform_L [447][10] <= LLR_448;					inform_L [448][10] <= LLR_449;					inform_L [449][10] <= LLR_450;					inform_L [450][10] <= LLR_451;					inform_L [451][10] <= LLR_452;					inform_L [452][10] <= LLR_453;					inform_L [453][10] <= LLR_454;					inform_L [454][10] <= LLR_455;					inform_L [455][10] <= LLR_456;					inform_L [456][10] <= LLR_457;					inform_L [457][10] <= LLR_458;					inform_L [458][10] <= LLR_459;					inform_L [459][10] <= LLR_460;					inform_L [460][10] <= LLR_461;					inform_L [461][10] <= LLR_462;					inform_L [462][10] <= LLR_463;					inform_L [463][10] <= LLR_464;					inform_L [464][10] <= LLR_465;					inform_L [465][10] <= LLR_466;					inform_L [466][10] <= LLR_467;					inform_L [467][10] <= LLR_468;					inform_L [468][10] <= LLR_469;					inform_L [469][10] <= LLR_470;					inform_L [470][10] <= LLR_471;					inform_L [471][10] <= LLR_472;					inform_L [472][10] <= LLR_473;					inform_L [473][10] <= LLR_474;					inform_L [474][10] <= LLR_475;					inform_L [475][10] <= LLR_476;					inform_L [476][10] <= LLR_477;					inform_L [477][10] <= LLR_478;					inform_L [478][10] <= LLR_479;					inform_L [479][10] <= LLR_480;					inform_L [480][10] <= LLR_481;					inform_L [481][10] <= LLR_482;					inform_L [482][10] <= LLR_483;					inform_L [483][10] <= LLR_484;					inform_L [484][10] <= LLR_485;					inform_L [485][10] <= LLR_486;					inform_L [486][10] <= LLR_487;					inform_L [487][10] <= LLR_488;					inform_L [488][10] <= LLR_489;					inform_L [489][10] <= LLR_490;					inform_L [490][10] <= LLR_491;					inform_L [491][10] <= LLR_492;					inform_L [492][10] <= LLR_493;					inform_L [493][10] <= LLR_494;					inform_L [494][10] <= LLR_495;					inform_L [495][10] <= LLR_496;					inform_L [496][10] <= LLR_497;					inform_L [497][10] <= LLR_498;					inform_L [498][10] <= LLR_499;					inform_L [499][10] <= LLR_500;					inform_L [500][10] <= LLR_501;					inform_L [501][10] <= LLR_502;					inform_L [502][10] <= LLR_503;					inform_L [503][10] <= LLR_504;					inform_L [504][10] <= LLR_505;					inform_L [505][10] <= LLR_506;					inform_L [506][10] <= LLR_507;					inform_L [507][10] <= LLR_508;					inform_L [508][10] <= LLR_509;					inform_L [509][10] <= LLR_510;					inform_L [510][10] <= LLR_511;					inform_L [511][10] <= LLR_512;					inform_L [512][10] <= LLR_513;					inform_L [513][10] <= LLR_514;					inform_L [514][10] <= LLR_515;					inform_L [515][10] <= LLR_516;					inform_L [516][10] <= LLR_517;					inform_L [517][10] <= LLR_518;					inform_L [518][10] <= LLR_519;					inform_L [519][10] <= LLR_520;					inform_L [520][10] <= LLR_521;					inform_L [521][10] <= LLR_522;					inform_L [522][10] <= LLR_523;					inform_L [523][10] <= LLR_524;					inform_L [524][10] <= LLR_525;					inform_L [525][10] <= LLR_526;					inform_L [526][10] <= LLR_527;					inform_L [527][10] <= LLR_528;					inform_L [528][10] <= LLR_529;					inform_L [529][10] <= LLR_530;					inform_L [530][10] <= LLR_531;					inform_L [531][10] <= LLR_532;					inform_L [532][10] <= LLR_533;					inform_L [533][10] <= LLR_534;					inform_L [534][10] <= LLR_535;					inform_L [535][10] <= LLR_536;					inform_L [536][10] <= LLR_537;					inform_L [537][10] <= LLR_538;					inform_L [538][10] <= LLR_539;					inform_L [539][10] <= LLR_540;					inform_L [540][10] <= LLR_541;					inform_L [541][10] <= LLR_542;					inform_L [542][10] <= LLR_543;					inform_L [543][10] <= LLR_544;					inform_L [544][10] <= LLR_545;					inform_L [545][10] <= LLR_546;					inform_L [546][10] <= LLR_547;					inform_L [547][10] <= LLR_548;					inform_L [548][10] <= LLR_549;					inform_L [549][10] <= LLR_550;					inform_L [550][10] <= LLR_551;					inform_L [551][10] <= LLR_552;					inform_L [552][10] <= LLR_553;					inform_L [553][10] <= LLR_554;					inform_L [554][10] <= LLR_555;					inform_L [555][10] <= LLR_556;					inform_L [556][10] <= LLR_557;					inform_L [557][10] <= LLR_558;					inform_L [558][10] <= LLR_559;					inform_L [559][10] <= LLR_560;					inform_L [560][10] <= LLR_561;					inform_L [561][10] <= LLR_562;					inform_L [562][10] <= LLR_563;					inform_L [563][10] <= LLR_564;					inform_L [564][10] <= LLR_565;					inform_L [565][10] <= LLR_566;					inform_L [566][10] <= LLR_567;					inform_L [567][10] <= LLR_568;					inform_L [568][10] <= LLR_569;					inform_L [569][10] <= LLR_570;					inform_L [570][10] <= LLR_571;					inform_L [571][10] <= LLR_572;					inform_L [572][10] <= LLR_573;					inform_L [573][10] <= LLR_574;					inform_L [574][10] <= LLR_575;					inform_L [575][10] <= LLR_576;					inform_L [576][10] <= LLR_577;					inform_L [577][10] <= LLR_578;					inform_L [578][10] <= LLR_579;					inform_L [579][10] <= LLR_580;					inform_L [580][10] <= LLR_581;					inform_L [581][10] <= LLR_582;					inform_L [582][10] <= LLR_583;					inform_L [583][10] <= LLR_584;					inform_L [584][10] <= LLR_585;					inform_L [585][10] <= LLR_586;					inform_L [586][10] <= LLR_587;					inform_L [587][10] <= LLR_588;					inform_L [588][10] <= LLR_589;					inform_L [589][10] <= LLR_590;					inform_L [590][10] <= LLR_591;					inform_L [591][10] <= LLR_592;					inform_L [592][10] <= LLR_593;					inform_L [593][10] <= LLR_594;					inform_L [594][10] <= LLR_595;					inform_L [595][10] <= LLR_596;					inform_L [596][10] <= LLR_597;					inform_L [597][10] <= LLR_598;					inform_L [598][10] <= LLR_599;					inform_L [599][10] <= LLR_600;					inform_L [600][10] <= LLR_601;					inform_L [601][10] <= LLR_602;					inform_L [602][10] <= LLR_603;					inform_L [603][10] <= LLR_604;					inform_L [604][10] <= LLR_605;					inform_L [605][10] <= LLR_606;					inform_L [606][10] <= LLR_607;					inform_L [607][10] <= LLR_608;					inform_L [608][10] <= LLR_609;					inform_L [609][10] <= LLR_610;					inform_L [610][10] <= LLR_611;					inform_L [611][10] <= LLR_612;					inform_L [612][10] <= LLR_613;					inform_L [613][10] <= LLR_614;					inform_L [614][10] <= LLR_615;					inform_L [615][10] <= LLR_616;					inform_L [616][10] <= LLR_617;					inform_L [617][10] <= LLR_618;					inform_L [618][10] <= LLR_619;					inform_L [619][10] <= LLR_620;					inform_L [620][10] <= LLR_621;					inform_L [621][10] <= LLR_622;					inform_L [622][10] <= LLR_623;					inform_L [623][10] <= LLR_624;					inform_L [624][10] <= LLR_625;					inform_L [625][10] <= LLR_626;					inform_L [626][10] <= LLR_627;					inform_L [627][10] <= LLR_628;					inform_L [628][10] <= LLR_629;					inform_L [629][10] <= LLR_630;					inform_L [630][10] <= LLR_631;					inform_L [631][10] <= LLR_632;					inform_L [632][10] <= LLR_633;					inform_L [633][10] <= LLR_634;					inform_L [634][10] <= LLR_635;					inform_L [635][10] <= LLR_636;					inform_L [636][10] <= LLR_637;					inform_L [637][10] <= LLR_638;					inform_L [638][10] <= LLR_639;					inform_L [639][10] <= LLR_640;					inform_L [640][10] <= LLR_641;					inform_L [641][10] <= LLR_642;					inform_L [642][10] <= LLR_643;					inform_L [643][10] <= LLR_644;					inform_L [644][10] <= LLR_645;					inform_L [645][10] <= LLR_646;					inform_L [646][10] <= LLR_647;					inform_L [647][10] <= LLR_648;					inform_L [648][10] <= LLR_649;					inform_L [649][10] <= LLR_650;					inform_L [650][10] <= LLR_651;					inform_L [651][10] <= LLR_652;					inform_L [652][10] <= LLR_653;					inform_L [653][10] <= LLR_654;					inform_L [654][10] <= LLR_655;					inform_L [655][10] <= LLR_656;					inform_L [656][10] <= LLR_657;					inform_L [657][10] <= LLR_658;					inform_L [658][10] <= LLR_659;					inform_L [659][10] <= LLR_660;					inform_L [660][10] <= LLR_661;					inform_L [661][10] <= LLR_662;					inform_L [662][10] <= LLR_663;					inform_L [663][10] <= LLR_664;					inform_L [664][10] <= LLR_665;					inform_L [665][10] <= LLR_666;					inform_L [666][10] <= LLR_667;					inform_L [667][10] <= LLR_668;					inform_L [668][10] <= LLR_669;					inform_L [669][10] <= LLR_670;					inform_L [670][10] <= LLR_671;					inform_L [671][10] <= LLR_672;					inform_L [672][10] <= LLR_673;					inform_L [673][10] <= LLR_674;					inform_L [674][10] <= LLR_675;					inform_L [675][10] <= LLR_676;					inform_L [676][10] <= LLR_677;					inform_L [677][10] <= LLR_678;					inform_L [678][10] <= LLR_679;					inform_L [679][10] <= LLR_680;					inform_L [680][10] <= LLR_681;					inform_L [681][10] <= LLR_682;					inform_L [682][10] <= LLR_683;					inform_L [683][10] <= LLR_684;					inform_L [684][10] <= LLR_685;					inform_L [685][10] <= LLR_686;					inform_L [686][10] <= LLR_687;					inform_L [687][10] <= LLR_688;					inform_L [688][10] <= LLR_689;					inform_L [689][10] <= LLR_690;					inform_L [690][10] <= LLR_691;					inform_L [691][10] <= LLR_692;					inform_L [692][10] <= LLR_693;					inform_L [693][10] <= LLR_694;					inform_L [694][10] <= LLR_695;					inform_L [695][10] <= LLR_696;					inform_L [696][10] <= LLR_697;					inform_L [697][10] <= LLR_698;					inform_L [698][10] <= LLR_699;					inform_L [699][10] <= LLR_700;					inform_L [700][10] <= LLR_701;					inform_L [701][10] <= LLR_702;					inform_L [702][10] <= LLR_703;					inform_L [703][10] <= LLR_704;					inform_L [704][10] <= LLR_705;					inform_L [705][10] <= LLR_706;					inform_L [706][10] <= LLR_707;					inform_L [707][10] <= LLR_708;					inform_L [708][10] <= LLR_709;					inform_L [709][10] <= LLR_710;					inform_L [710][10] <= LLR_711;					inform_L [711][10] <= LLR_712;					inform_L [712][10] <= LLR_713;					inform_L [713][10] <= LLR_714;					inform_L [714][10] <= LLR_715;					inform_L [715][10] <= LLR_716;					inform_L [716][10] <= LLR_717;					inform_L [717][10] <= LLR_718;					inform_L [718][10] <= LLR_719;					inform_L [719][10] <= LLR_720;					inform_L [720][10] <= LLR_721;					inform_L [721][10] <= LLR_722;					inform_L [722][10] <= LLR_723;					inform_L [723][10] <= LLR_724;					inform_L [724][10] <= LLR_725;					inform_L [725][10] <= LLR_726;					inform_L [726][10] <= LLR_727;					inform_L [727][10] <= LLR_728;					inform_L [728][10] <= LLR_729;					inform_L [729][10] <= LLR_730;					inform_L [730][10] <= LLR_731;					inform_L [731][10] <= LLR_732;					inform_L [732][10] <= LLR_733;					inform_L [733][10] <= LLR_734;					inform_L [734][10] <= LLR_735;					inform_L [735][10] <= LLR_736;					inform_L [736][10] <= LLR_737;					inform_L [737][10] <= LLR_738;					inform_L [738][10] <= LLR_739;					inform_L [739][10] <= LLR_740;					inform_L [740][10] <= LLR_741;					inform_L [741][10] <= LLR_742;					inform_L [742][10] <= LLR_743;					inform_L [743][10] <= LLR_744;					inform_L [744][10] <= LLR_745;					inform_L [745][10] <= LLR_746;					inform_L [746][10] <= LLR_747;					inform_L [747][10] <= LLR_748;					inform_L [748][10] <= LLR_749;					inform_L [749][10] <= LLR_750;					inform_L [750][10] <= LLR_751;					inform_L [751][10] <= LLR_752;					inform_L [752][10] <= LLR_753;					inform_L [753][10] <= LLR_754;					inform_L [754][10] <= LLR_755;					inform_L [755][10] <= LLR_756;					inform_L [756][10] <= LLR_757;					inform_L [757][10] <= LLR_758;					inform_L [758][10] <= LLR_759;					inform_L [759][10] <= LLR_760;					inform_L [760][10] <= LLR_761;					inform_L [761][10] <= LLR_762;					inform_L [762][10] <= LLR_763;					inform_L [763][10] <= LLR_764;					inform_L [764][10] <= LLR_765;					inform_L [765][10] <= LLR_766;					inform_L [766][10] <= LLR_767;					inform_L [767][10] <= LLR_768;					inform_L [768][10] <= LLR_769;					inform_L [769][10] <= LLR_770;					inform_L [770][10] <= LLR_771;					inform_L [771][10] <= LLR_772;					inform_L [772][10] <= LLR_773;					inform_L [773][10] <= LLR_774;					inform_L [774][10] <= LLR_775;					inform_L [775][10] <= LLR_776;					inform_L [776][10] <= LLR_777;					inform_L [777][10] <= LLR_778;					inform_L [778][10] <= LLR_779;					inform_L [779][10] <= LLR_780;					inform_L [780][10] <= LLR_781;					inform_L [781][10] <= LLR_782;					inform_L [782][10] <= LLR_783;					inform_L [783][10] <= LLR_784;					inform_L [784][10] <= LLR_785;					inform_L [785][10] <= LLR_786;					inform_L [786][10] <= LLR_787;					inform_L [787][10] <= LLR_788;					inform_L [788][10] <= LLR_789;					inform_L [789][10] <= LLR_790;					inform_L [790][10] <= LLR_791;					inform_L [791][10] <= LLR_792;					inform_L [792][10] <= LLR_793;					inform_L [793][10] <= LLR_794;					inform_L [794][10] <= LLR_795;					inform_L [795][10] <= LLR_796;					inform_L [796][10] <= LLR_797;					inform_L [797][10] <= LLR_798;					inform_L [798][10] <= LLR_799;					inform_L [799][10] <= LLR_800;					inform_L [800][10] <= LLR_801;					inform_L [801][10] <= LLR_802;					inform_L [802][10] <= LLR_803;					inform_L [803][10] <= LLR_804;					inform_L [804][10] <= LLR_805;					inform_L [805][10] <= LLR_806;					inform_L [806][10] <= LLR_807;					inform_L [807][10] <= LLR_808;					inform_L [808][10] <= LLR_809;					inform_L [809][10] <= LLR_810;					inform_L [810][10] <= LLR_811;					inform_L [811][10] <= LLR_812;					inform_L [812][10] <= LLR_813;					inform_L [813][10] <= LLR_814;					inform_L [814][10] <= LLR_815;					inform_L [815][10] <= LLR_816;					inform_L [816][10] <= LLR_817;					inform_L [817][10] <= LLR_818;					inform_L [818][10] <= LLR_819;					inform_L [819][10] <= LLR_820;					inform_L [820][10] <= LLR_821;					inform_L [821][10] <= LLR_822;					inform_L [822][10] <= LLR_823;					inform_L [823][10] <= LLR_824;					inform_L [824][10] <= LLR_825;					inform_L [825][10] <= LLR_826;					inform_L [826][10] <= LLR_827;					inform_L [827][10] <= LLR_828;					inform_L [828][10] <= LLR_829;					inform_L [829][10] <= LLR_830;					inform_L [830][10] <= LLR_831;					inform_L [831][10] <= LLR_832;					inform_L [832][10] <= LLR_833;					inform_L [833][10] <= LLR_834;					inform_L [834][10] <= LLR_835;					inform_L [835][10] <= LLR_836;					inform_L [836][10] <= LLR_837;					inform_L [837][10] <= LLR_838;					inform_L [838][10] <= LLR_839;					inform_L [839][10] <= LLR_840;					inform_L [840][10] <= LLR_841;					inform_L [841][10] <= LLR_842;					inform_L [842][10] <= LLR_843;					inform_L [843][10] <= LLR_844;					inform_L [844][10] <= LLR_845;					inform_L [845][10] <= LLR_846;					inform_L [846][10] <= LLR_847;					inform_L [847][10] <= LLR_848;					inform_L [848][10] <= LLR_849;					inform_L [849][10] <= LLR_850;					inform_L [850][10] <= LLR_851;					inform_L [851][10] <= LLR_852;					inform_L [852][10] <= LLR_853;					inform_L [853][10] <= LLR_854;					inform_L [854][10] <= LLR_855;					inform_L [855][10] <= LLR_856;					inform_L [856][10] <= LLR_857;					inform_L [857][10] <= LLR_858;					inform_L [858][10] <= LLR_859;					inform_L [859][10] <= LLR_860;					inform_L [860][10] <= LLR_861;					inform_L [861][10] <= LLR_862;					inform_L [862][10] <= LLR_863;					inform_L [863][10] <= LLR_864;					inform_L [864][10] <= LLR_865;					inform_L [865][10] <= LLR_866;					inform_L [866][10] <= LLR_867;					inform_L [867][10] <= LLR_868;					inform_L [868][10] <= LLR_869;					inform_L [869][10] <= LLR_870;					inform_L [870][10] <= LLR_871;					inform_L [871][10] <= LLR_872;					inform_L [872][10] <= LLR_873;					inform_L [873][10] <= LLR_874;					inform_L [874][10] <= LLR_875;					inform_L [875][10] <= LLR_876;					inform_L [876][10] <= LLR_877;					inform_L [877][10] <= LLR_878;					inform_L [878][10] <= LLR_879;					inform_L [879][10] <= LLR_880;					inform_L [880][10] <= LLR_881;					inform_L [881][10] <= LLR_882;					inform_L [882][10] <= LLR_883;					inform_L [883][10] <= LLR_884;					inform_L [884][10] <= LLR_885;					inform_L [885][10] <= LLR_886;					inform_L [886][10] <= LLR_887;					inform_L [887][10] <= LLR_888;					inform_L [888][10] <= LLR_889;					inform_L [889][10] <= LLR_890;					inform_L [890][10] <= LLR_891;					inform_L [891][10] <= LLR_892;					inform_L [892][10] <= LLR_893;					inform_L [893][10] <= LLR_894;					inform_L [894][10] <= LLR_895;					inform_L [895][10] <= LLR_896;					inform_L [896][10] <= LLR_897;					inform_L [897][10] <= LLR_898;					inform_L [898][10] <= LLR_899;					inform_L [899][10] <= LLR_900;					inform_L [900][10] <= LLR_901;					inform_L [901][10] <= LLR_902;					inform_L [902][10] <= LLR_903;					inform_L [903][10] <= LLR_904;					inform_L [904][10] <= LLR_905;					inform_L [905][10] <= LLR_906;					inform_L [906][10] <= LLR_907;					inform_L [907][10] <= LLR_908;					inform_L [908][10] <= LLR_909;					inform_L [909][10] <= LLR_910;					inform_L [910][10] <= LLR_911;					inform_L [911][10] <= LLR_912;					inform_L [912][10] <= LLR_913;					inform_L [913][10] <= LLR_914;					inform_L [914][10] <= LLR_915;					inform_L [915][10] <= LLR_916;					inform_L [916][10] <= LLR_917;					inform_L [917][10] <= LLR_918;					inform_L [918][10] <= LLR_919;					inform_L [919][10] <= LLR_920;					inform_L [920][10] <= LLR_921;					inform_L [921][10] <= LLR_922;					inform_L [922][10] <= LLR_923;					inform_L [923][10] <= LLR_924;					inform_L [924][10] <= LLR_925;					inform_L [925][10] <= LLR_926;					inform_L [926][10] <= LLR_927;					inform_L [927][10] <= LLR_928;					inform_L [928][10] <= LLR_929;					inform_L [929][10] <= LLR_930;					inform_L [930][10] <= LLR_931;					inform_L [931][10] <= LLR_932;					inform_L [932][10] <= LLR_933;					inform_L [933][10] <= LLR_934;					inform_L [934][10] <= LLR_935;					inform_L [935][10] <= LLR_936;					inform_L [936][10] <= LLR_937;					inform_L [937][10] <= LLR_938;					inform_L [938][10] <= LLR_939;					inform_L [939][10] <= LLR_940;					inform_L [940][10] <= LLR_941;					inform_L [941][10] <= LLR_942;					inform_L [942][10] <= LLR_943;					inform_L [943][10] <= LLR_944;					inform_L [944][10] <= LLR_945;					inform_L [945][10] <= LLR_946;					inform_L [946][10] <= LLR_947;					inform_L [947][10] <= LLR_948;					inform_L [948][10] <= LLR_949;					inform_L [949][10] <= LLR_950;					inform_L [950][10] <= LLR_951;					inform_L [951][10] <= LLR_952;					inform_L [952][10] <= LLR_953;					inform_L [953][10] <= LLR_954;					inform_L [954][10] <= LLR_955;					inform_L [955][10] <= LLR_956;					inform_L [956][10] <= LLR_957;					inform_L [957][10] <= LLR_958;					inform_L [958][10] <= LLR_959;					inform_L [959][10] <= LLR_960;					inform_L [960][10] <= LLR_961;					inform_L [961][10] <= LLR_962;					inform_L [962][10] <= LLR_963;					inform_L [963][10] <= LLR_964;					inform_L [964][10] <= LLR_965;					inform_L [965][10] <= LLR_966;					inform_L [966][10] <= LLR_967;					inform_L [967][10] <= LLR_968;					inform_L [968][10] <= LLR_969;					inform_L [969][10] <= LLR_970;					inform_L [970][10] <= LLR_971;					inform_L [971][10] <= LLR_972;					inform_L [972][10] <= LLR_973;					inform_L [973][10] <= LLR_974;					inform_L [974][10] <= LLR_975;					inform_L [975][10] <= LLR_976;					inform_L [976][10] <= LLR_977;					inform_L [977][10] <= LLR_978;					inform_L [978][10] <= LLR_979;					inform_L [979][10] <= LLR_980;					inform_L [980][10] <= LLR_981;					inform_L [981][10] <= LLR_982;					inform_L [982][10] <= LLR_983;					inform_L [983][10] <= LLR_984;					inform_L [984][10] <= LLR_985;					inform_L [985][10] <= LLR_986;					inform_L [986][10] <= LLR_987;					inform_L [987][10] <= LLR_988;					inform_L [988][10] <= LLR_989;					inform_L [989][10] <= LLR_990;					inform_L [990][10] <= LLR_991;					inform_L [991][10] <= LLR_992;					inform_L [992][10] <= LLR_993;					inform_L [993][10] <= LLR_994;					inform_L [994][10] <= LLR_995;					inform_L [995][10] <= LLR_996;					inform_L [996][10] <= LLR_997;					inform_L [997][10] <= LLR_998;					inform_L [998][10] <= LLR_999;					inform_L [999][10] <= LLR_1000;					inform_L [1000][10] <= LLR_1001;					inform_L [1001][10] <= LLR_1002;					inform_L [1002][10] <= LLR_1003;					inform_L [1003][10] <= LLR_1004;					inform_L [1004][10] <= LLR_1005;					inform_L [1005][10] <= LLR_1006;					inform_L [1006][10] <= LLR_1007;					inform_L [1007][10] <= LLR_1008;					inform_L [1008][10] <= LLR_1009;					inform_L [1009][10] <= LLR_1010;					inform_L [1010][10] <= LLR_1011;					inform_L [1011][10] <= LLR_1012;					inform_L [1012][10] <= LLR_1013;					inform_L [1013][10] <= LLR_1014;					inform_L [1014][10] <= LLR_1015;					inform_L [1015][10] <= LLR_1016;					inform_L [1016][10] <= LLR_1017;					inform_L [1017][10] <= LLR_1018;					inform_L [1018][10] <= LLR_1019;					inform_L [1019][10] <= LLR_1020;					inform_L [1020][10] <= LLR_1021;					inform_L [1021][10] <= LLR_1022;					inform_L [1022][10] <= LLR_1023;					inform_L [1023][10] <= LLR_1024;				end				for (x = 0; x < 1024; x = x + 1)					for (y = 0; y < 10; y = y + 1)					begin						inform_R[x][y+1] <= 8'd0;						inform_L[x][y] <= 8'd0;					end			end
		endcase	end
	assign bp_over_flag = (itera_time == `iteration_times + 1) ? 1 : 0;
	always @(*)	begin		case (w2r)			1:			begin				r_cell_reg[0] = inform_R[0][0];				r_cell_reg[1] = inform_R[1][0];				r_cell_reg[2] = inform_R[2][0];				r_cell_reg[3] = inform_R[3][0];				r_cell_reg[4] = inform_R[4][0];				r_cell_reg[5] = inform_R[5][0];				r_cell_reg[6] = inform_R[6][0];				r_cell_reg[7] = inform_R[7][0];				r_cell_reg[8] = inform_R[8][0];				r_cell_reg[9] = inform_R[9][0];				r_cell_reg[10] = inform_R[10][0];				r_cell_reg[11] = inform_R[11][0];				r_cell_reg[12] = inform_R[12][0];				r_cell_reg[13] = inform_R[13][0];				r_cell_reg[14] = inform_R[14][0];				r_cell_reg[15] = inform_R[15][0];				r_cell_reg[16] = inform_R[16][0];				r_cell_reg[17] = inform_R[17][0];				r_cell_reg[18] = inform_R[18][0];				r_cell_reg[19] = inform_R[19][0];				r_cell_reg[20] = inform_R[20][0];				r_cell_reg[21] = inform_R[21][0];				r_cell_reg[22] = inform_R[22][0];				r_cell_reg[23] = inform_R[23][0];				r_cell_reg[24] = inform_R[24][0];				r_cell_reg[25] = inform_R[25][0];				r_cell_reg[26] = inform_R[26][0];				r_cell_reg[27] = inform_R[27][0];				r_cell_reg[28] = inform_R[28][0];				r_cell_reg[29] = inform_R[29][0];				r_cell_reg[30] = inform_R[30][0];				r_cell_reg[31] = inform_R[31][0];				r_cell_reg[32] = inform_R[32][0];				r_cell_reg[33] = inform_R[33][0];				r_cell_reg[34] = inform_R[34][0];				r_cell_reg[35] = inform_R[35][0];				r_cell_reg[36] = inform_R[36][0];				r_cell_reg[37] = inform_R[37][0];				r_cell_reg[38] = inform_R[38][0];				r_cell_reg[39] = inform_R[39][0];				r_cell_reg[40] = inform_R[40][0];				r_cell_reg[41] = inform_R[41][0];				r_cell_reg[42] = inform_R[42][0];				r_cell_reg[43] = inform_R[43][0];				r_cell_reg[44] = inform_R[44][0];				r_cell_reg[45] = inform_R[45][0];				r_cell_reg[46] = inform_R[46][0];				r_cell_reg[47] = inform_R[47][0];				r_cell_reg[48] = inform_R[48][0];				r_cell_reg[49] = inform_R[49][0];				r_cell_reg[50] = inform_R[50][0];				r_cell_reg[51] = inform_R[51][0];				r_cell_reg[52] = inform_R[52][0];				r_cell_reg[53] = inform_R[53][0];				r_cell_reg[54] = inform_R[54][0];				r_cell_reg[55] = inform_R[55][0];				r_cell_reg[56] = inform_R[56][0];				r_cell_reg[57] = inform_R[57][0];				r_cell_reg[58] = inform_R[58][0];				r_cell_reg[59] = inform_R[59][0];				r_cell_reg[60] = inform_R[60][0];				r_cell_reg[61] = inform_R[61][0];				r_cell_reg[62] = inform_R[62][0];				r_cell_reg[63] = inform_R[63][0];				r_cell_reg[64] = inform_R[64][0];				r_cell_reg[65] = inform_R[65][0];				r_cell_reg[66] = inform_R[66][0];				r_cell_reg[67] = inform_R[67][0];				r_cell_reg[68] = inform_R[68][0];				r_cell_reg[69] = inform_R[69][0];				r_cell_reg[70] = inform_R[70][0];				r_cell_reg[71] = inform_R[71][0];				r_cell_reg[72] = inform_R[72][0];				r_cell_reg[73] = inform_R[73][0];				r_cell_reg[74] = inform_R[74][0];				r_cell_reg[75] = inform_R[75][0];				r_cell_reg[76] = inform_R[76][0];				r_cell_reg[77] = inform_R[77][0];				r_cell_reg[78] = inform_R[78][0];				r_cell_reg[79] = inform_R[79][0];				r_cell_reg[80] = inform_R[80][0];				r_cell_reg[81] = inform_R[81][0];				r_cell_reg[82] = inform_R[82][0];				r_cell_reg[83] = inform_R[83][0];				r_cell_reg[84] = inform_R[84][0];				r_cell_reg[85] = inform_R[85][0];				r_cell_reg[86] = inform_R[86][0];				r_cell_reg[87] = inform_R[87][0];				r_cell_reg[88] = inform_R[88][0];				r_cell_reg[89] = inform_R[89][0];				r_cell_reg[90] = inform_R[90][0];				r_cell_reg[91] = inform_R[91][0];				r_cell_reg[92] = inform_R[92][0];				r_cell_reg[93] = inform_R[93][0];				r_cell_reg[94] = inform_R[94][0];				r_cell_reg[95] = inform_R[95][0];				r_cell_reg[96] = inform_R[96][0];				r_cell_reg[97] = inform_R[97][0];				r_cell_reg[98] = inform_R[98][0];				r_cell_reg[99] = inform_R[99][0];				r_cell_reg[100] = inform_R[100][0];				r_cell_reg[101] = inform_R[101][0];				r_cell_reg[102] = inform_R[102][0];				r_cell_reg[103] = inform_R[103][0];				r_cell_reg[104] = inform_R[104][0];				r_cell_reg[105] = inform_R[105][0];				r_cell_reg[106] = inform_R[106][0];				r_cell_reg[107] = inform_R[107][0];				r_cell_reg[108] = inform_R[108][0];				r_cell_reg[109] = inform_R[109][0];				r_cell_reg[110] = inform_R[110][0];				r_cell_reg[111] = inform_R[111][0];				r_cell_reg[112] = inform_R[112][0];				r_cell_reg[113] = inform_R[113][0];				r_cell_reg[114] = inform_R[114][0];				r_cell_reg[115] = inform_R[115][0];				r_cell_reg[116] = inform_R[116][0];				r_cell_reg[117] = inform_R[117][0];				r_cell_reg[118] = inform_R[118][0];				r_cell_reg[119] = inform_R[119][0];				r_cell_reg[120] = inform_R[120][0];				r_cell_reg[121] = inform_R[121][0];				r_cell_reg[122] = inform_R[122][0];				r_cell_reg[123] = inform_R[123][0];				r_cell_reg[124] = inform_R[124][0];				r_cell_reg[125] = inform_R[125][0];				r_cell_reg[126] = inform_R[126][0];				r_cell_reg[127] = inform_R[127][0];				r_cell_reg[128] = inform_R[128][0];				r_cell_reg[129] = inform_R[129][0];				r_cell_reg[130] = inform_R[130][0];				r_cell_reg[131] = inform_R[131][0];				r_cell_reg[132] = inform_R[132][0];				r_cell_reg[133] = inform_R[133][0];				r_cell_reg[134] = inform_R[134][0];				r_cell_reg[135] = inform_R[135][0];				r_cell_reg[136] = inform_R[136][0];				r_cell_reg[137] = inform_R[137][0];				r_cell_reg[138] = inform_R[138][0];				r_cell_reg[139] = inform_R[139][0];				r_cell_reg[140] = inform_R[140][0];				r_cell_reg[141] = inform_R[141][0];				r_cell_reg[142] = inform_R[142][0];				r_cell_reg[143] = inform_R[143][0];				r_cell_reg[144] = inform_R[144][0];				r_cell_reg[145] = inform_R[145][0];				r_cell_reg[146] = inform_R[146][0];				r_cell_reg[147] = inform_R[147][0];				r_cell_reg[148] = inform_R[148][0];				r_cell_reg[149] = inform_R[149][0];				r_cell_reg[150] = inform_R[150][0];				r_cell_reg[151] = inform_R[151][0];				r_cell_reg[152] = inform_R[152][0];				r_cell_reg[153] = inform_R[153][0];				r_cell_reg[154] = inform_R[154][0];				r_cell_reg[155] = inform_R[155][0];				r_cell_reg[156] = inform_R[156][0];				r_cell_reg[157] = inform_R[157][0];				r_cell_reg[158] = inform_R[158][0];				r_cell_reg[159] = inform_R[159][0];				r_cell_reg[160] = inform_R[160][0];				r_cell_reg[161] = inform_R[161][0];				r_cell_reg[162] = inform_R[162][0];				r_cell_reg[163] = inform_R[163][0];				r_cell_reg[164] = inform_R[164][0];				r_cell_reg[165] = inform_R[165][0];				r_cell_reg[166] = inform_R[166][0];				r_cell_reg[167] = inform_R[167][0];				r_cell_reg[168] = inform_R[168][0];				r_cell_reg[169] = inform_R[169][0];				r_cell_reg[170] = inform_R[170][0];				r_cell_reg[171] = inform_R[171][0];				r_cell_reg[172] = inform_R[172][0];				r_cell_reg[173] = inform_R[173][0];				r_cell_reg[174] = inform_R[174][0];				r_cell_reg[175] = inform_R[175][0];				r_cell_reg[176] = inform_R[176][0];				r_cell_reg[177] = inform_R[177][0];				r_cell_reg[178] = inform_R[178][0];				r_cell_reg[179] = inform_R[179][0];				r_cell_reg[180] = inform_R[180][0];				r_cell_reg[181] = inform_R[181][0];				r_cell_reg[182] = inform_R[182][0];				r_cell_reg[183] = inform_R[183][0];				r_cell_reg[184] = inform_R[184][0];				r_cell_reg[185] = inform_R[185][0];				r_cell_reg[186] = inform_R[186][0];				r_cell_reg[187] = inform_R[187][0];				r_cell_reg[188] = inform_R[188][0];				r_cell_reg[189] = inform_R[189][0];				r_cell_reg[190] = inform_R[190][0];				r_cell_reg[191] = inform_R[191][0];				r_cell_reg[192] = inform_R[192][0];				r_cell_reg[193] = inform_R[193][0];				r_cell_reg[194] = inform_R[194][0];				r_cell_reg[195] = inform_R[195][0];				r_cell_reg[196] = inform_R[196][0];				r_cell_reg[197] = inform_R[197][0];				r_cell_reg[198] = inform_R[198][0];				r_cell_reg[199] = inform_R[199][0];				r_cell_reg[200] = inform_R[200][0];				r_cell_reg[201] = inform_R[201][0];				r_cell_reg[202] = inform_R[202][0];				r_cell_reg[203] = inform_R[203][0];				r_cell_reg[204] = inform_R[204][0];				r_cell_reg[205] = inform_R[205][0];				r_cell_reg[206] = inform_R[206][0];				r_cell_reg[207] = inform_R[207][0];				r_cell_reg[208] = inform_R[208][0];				r_cell_reg[209] = inform_R[209][0];				r_cell_reg[210] = inform_R[210][0];				r_cell_reg[211] = inform_R[211][0];				r_cell_reg[212] = inform_R[212][0];				r_cell_reg[213] = inform_R[213][0];				r_cell_reg[214] = inform_R[214][0];				r_cell_reg[215] = inform_R[215][0];				r_cell_reg[216] = inform_R[216][0];				r_cell_reg[217] = inform_R[217][0];				r_cell_reg[218] = inform_R[218][0];				r_cell_reg[219] = inform_R[219][0];				r_cell_reg[220] = inform_R[220][0];				r_cell_reg[221] = inform_R[221][0];				r_cell_reg[222] = inform_R[222][0];				r_cell_reg[223] = inform_R[223][0];				r_cell_reg[224] = inform_R[224][0];				r_cell_reg[225] = inform_R[225][0];				r_cell_reg[226] = inform_R[226][0];				r_cell_reg[227] = inform_R[227][0];				r_cell_reg[228] = inform_R[228][0];				r_cell_reg[229] = inform_R[229][0];				r_cell_reg[230] = inform_R[230][0];				r_cell_reg[231] = inform_R[231][0];				r_cell_reg[232] = inform_R[232][0];				r_cell_reg[233] = inform_R[233][0];				r_cell_reg[234] = inform_R[234][0];				r_cell_reg[235] = inform_R[235][0];				r_cell_reg[236] = inform_R[236][0];				r_cell_reg[237] = inform_R[237][0];				r_cell_reg[238] = inform_R[238][0];				r_cell_reg[239] = inform_R[239][0];				r_cell_reg[240] = inform_R[240][0];				r_cell_reg[241] = inform_R[241][0];				r_cell_reg[242] = inform_R[242][0];				r_cell_reg[243] = inform_R[243][0];				r_cell_reg[244] = inform_R[244][0];				r_cell_reg[245] = inform_R[245][0];				r_cell_reg[246] = inform_R[246][0];				r_cell_reg[247] = inform_R[247][0];				r_cell_reg[248] = inform_R[248][0];				r_cell_reg[249] = inform_R[249][0];				r_cell_reg[250] = inform_R[250][0];				r_cell_reg[251] = inform_R[251][0];				r_cell_reg[252] = inform_R[252][0];				r_cell_reg[253] = inform_R[253][0];				r_cell_reg[254] = inform_R[254][0];				r_cell_reg[255] = inform_R[255][0];				r_cell_reg[256] = inform_R[256][0];				r_cell_reg[257] = inform_R[257][0];				r_cell_reg[258] = inform_R[258][0];				r_cell_reg[259] = inform_R[259][0];				r_cell_reg[260] = inform_R[260][0];				r_cell_reg[261] = inform_R[261][0];				r_cell_reg[262] = inform_R[262][0];				r_cell_reg[263] = inform_R[263][0];				r_cell_reg[264] = inform_R[264][0];				r_cell_reg[265] = inform_R[265][0];				r_cell_reg[266] = inform_R[266][0];				r_cell_reg[267] = inform_R[267][0];				r_cell_reg[268] = inform_R[268][0];				r_cell_reg[269] = inform_R[269][0];				r_cell_reg[270] = inform_R[270][0];				r_cell_reg[271] = inform_R[271][0];				r_cell_reg[272] = inform_R[272][0];				r_cell_reg[273] = inform_R[273][0];				r_cell_reg[274] = inform_R[274][0];				r_cell_reg[275] = inform_R[275][0];				r_cell_reg[276] = inform_R[276][0];				r_cell_reg[277] = inform_R[277][0];				r_cell_reg[278] = inform_R[278][0];				r_cell_reg[279] = inform_R[279][0];				r_cell_reg[280] = inform_R[280][0];				r_cell_reg[281] = inform_R[281][0];				r_cell_reg[282] = inform_R[282][0];				r_cell_reg[283] = inform_R[283][0];				r_cell_reg[284] = inform_R[284][0];				r_cell_reg[285] = inform_R[285][0];				r_cell_reg[286] = inform_R[286][0];				r_cell_reg[287] = inform_R[287][0];				r_cell_reg[288] = inform_R[288][0];				r_cell_reg[289] = inform_R[289][0];				r_cell_reg[290] = inform_R[290][0];				r_cell_reg[291] = inform_R[291][0];				r_cell_reg[292] = inform_R[292][0];				r_cell_reg[293] = inform_R[293][0];				r_cell_reg[294] = inform_R[294][0];				r_cell_reg[295] = inform_R[295][0];				r_cell_reg[296] = inform_R[296][0];				r_cell_reg[297] = inform_R[297][0];				r_cell_reg[298] = inform_R[298][0];				r_cell_reg[299] = inform_R[299][0];				r_cell_reg[300] = inform_R[300][0];				r_cell_reg[301] = inform_R[301][0];				r_cell_reg[302] = inform_R[302][0];				r_cell_reg[303] = inform_R[303][0];				r_cell_reg[304] = inform_R[304][0];				r_cell_reg[305] = inform_R[305][0];				r_cell_reg[306] = inform_R[306][0];				r_cell_reg[307] = inform_R[307][0];				r_cell_reg[308] = inform_R[308][0];				r_cell_reg[309] = inform_R[309][0];				r_cell_reg[310] = inform_R[310][0];				r_cell_reg[311] = inform_R[311][0];				r_cell_reg[312] = inform_R[312][0];				r_cell_reg[313] = inform_R[313][0];				r_cell_reg[314] = inform_R[314][0];				r_cell_reg[315] = inform_R[315][0];				r_cell_reg[316] = inform_R[316][0];				r_cell_reg[317] = inform_R[317][0];				r_cell_reg[318] = inform_R[318][0];				r_cell_reg[319] = inform_R[319][0];				r_cell_reg[320] = inform_R[320][0];				r_cell_reg[321] = inform_R[321][0];				r_cell_reg[322] = inform_R[322][0];				r_cell_reg[323] = inform_R[323][0];				r_cell_reg[324] = inform_R[324][0];				r_cell_reg[325] = inform_R[325][0];				r_cell_reg[326] = inform_R[326][0];				r_cell_reg[327] = inform_R[327][0];				r_cell_reg[328] = inform_R[328][0];				r_cell_reg[329] = inform_R[329][0];				r_cell_reg[330] = inform_R[330][0];				r_cell_reg[331] = inform_R[331][0];				r_cell_reg[332] = inform_R[332][0];				r_cell_reg[333] = inform_R[333][0];				r_cell_reg[334] = inform_R[334][0];				r_cell_reg[335] = inform_R[335][0];				r_cell_reg[336] = inform_R[336][0];				r_cell_reg[337] = inform_R[337][0];				r_cell_reg[338] = inform_R[338][0];				r_cell_reg[339] = inform_R[339][0];				r_cell_reg[340] = inform_R[340][0];				r_cell_reg[341] = inform_R[341][0];				r_cell_reg[342] = inform_R[342][0];				r_cell_reg[343] = inform_R[343][0];				r_cell_reg[344] = inform_R[344][0];				r_cell_reg[345] = inform_R[345][0];				r_cell_reg[346] = inform_R[346][0];				r_cell_reg[347] = inform_R[347][0];				r_cell_reg[348] = inform_R[348][0];				r_cell_reg[349] = inform_R[349][0];				r_cell_reg[350] = inform_R[350][0];				r_cell_reg[351] = inform_R[351][0];				r_cell_reg[352] = inform_R[352][0];				r_cell_reg[353] = inform_R[353][0];				r_cell_reg[354] = inform_R[354][0];				r_cell_reg[355] = inform_R[355][0];				r_cell_reg[356] = inform_R[356][0];				r_cell_reg[357] = inform_R[357][0];				r_cell_reg[358] = inform_R[358][0];				r_cell_reg[359] = inform_R[359][0];				r_cell_reg[360] = inform_R[360][0];				r_cell_reg[361] = inform_R[361][0];				r_cell_reg[362] = inform_R[362][0];				r_cell_reg[363] = inform_R[363][0];				r_cell_reg[364] = inform_R[364][0];				r_cell_reg[365] = inform_R[365][0];				r_cell_reg[366] = inform_R[366][0];				r_cell_reg[367] = inform_R[367][0];				r_cell_reg[368] = inform_R[368][0];				r_cell_reg[369] = inform_R[369][0];				r_cell_reg[370] = inform_R[370][0];				r_cell_reg[371] = inform_R[371][0];				r_cell_reg[372] = inform_R[372][0];				r_cell_reg[373] = inform_R[373][0];				r_cell_reg[374] = inform_R[374][0];				r_cell_reg[375] = inform_R[375][0];				r_cell_reg[376] = inform_R[376][0];				r_cell_reg[377] = inform_R[377][0];				r_cell_reg[378] = inform_R[378][0];				r_cell_reg[379] = inform_R[379][0];				r_cell_reg[380] = inform_R[380][0];				r_cell_reg[381] = inform_R[381][0];				r_cell_reg[382] = inform_R[382][0];				r_cell_reg[383] = inform_R[383][0];				r_cell_reg[384] = inform_R[384][0];				r_cell_reg[385] = inform_R[385][0];				r_cell_reg[386] = inform_R[386][0];				r_cell_reg[387] = inform_R[387][0];				r_cell_reg[388] = inform_R[388][0];				r_cell_reg[389] = inform_R[389][0];				r_cell_reg[390] = inform_R[390][0];				r_cell_reg[391] = inform_R[391][0];				r_cell_reg[392] = inform_R[392][0];				r_cell_reg[393] = inform_R[393][0];				r_cell_reg[394] = inform_R[394][0];				r_cell_reg[395] = inform_R[395][0];				r_cell_reg[396] = inform_R[396][0];				r_cell_reg[397] = inform_R[397][0];				r_cell_reg[398] = inform_R[398][0];				r_cell_reg[399] = inform_R[399][0];				r_cell_reg[400] = inform_R[400][0];				r_cell_reg[401] = inform_R[401][0];				r_cell_reg[402] = inform_R[402][0];				r_cell_reg[403] = inform_R[403][0];				r_cell_reg[404] = inform_R[404][0];				r_cell_reg[405] = inform_R[405][0];				r_cell_reg[406] = inform_R[406][0];				r_cell_reg[407] = inform_R[407][0];				r_cell_reg[408] = inform_R[408][0];				r_cell_reg[409] = inform_R[409][0];				r_cell_reg[410] = inform_R[410][0];				r_cell_reg[411] = inform_R[411][0];				r_cell_reg[412] = inform_R[412][0];				r_cell_reg[413] = inform_R[413][0];				r_cell_reg[414] = inform_R[414][0];				r_cell_reg[415] = inform_R[415][0];				r_cell_reg[416] = inform_R[416][0];				r_cell_reg[417] = inform_R[417][0];				r_cell_reg[418] = inform_R[418][0];				r_cell_reg[419] = inform_R[419][0];				r_cell_reg[420] = inform_R[420][0];				r_cell_reg[421] = inform_R[421][0];				r_cell_reg[422] = inform_R[422][0];				r_cell_reg[423] = inform_R[423][0];				r_cell_reg[424] = inform_R[424][0];				r_cell_reg[425] = inform_R[425][0];				r_cell_reg[426] = inform_R[426][0];				r_cell_reg[427] = inform_R[427][0];				r_cell_reg[428] = inform_R[428][0];				r_cell_reg[429] = inform_R[429][0];				r_cell_reg[430] = inform_R[430][0];				r_cell_reg[431] = inform_R[431][0];				r_cell_reg[432] = inform_R[432][0];				r_cell_reg[433] = inform_R[433][0];				r_cell_reg[434] = inform_R[434][0];				r_cell_reg[435] = inform_R[435][0];				r_cell_reg[436] = inform_R[436][0];				r_cell_reg[437] = inform_R[437][0];				r_cell_reg[438] = inform_R[438][0];				r_cell_reg[439] = inform_R[439][0];				r_cell_reg[440] = inform_R[440][0];				r_cell_reg[441] = inform_R[441][0];				r_cell_reg[442] = inform_R[442][0];				r_cell_reg[443] = inform_R[443][0];				r_cell_reg[444] = inform_R[444][0];				r_cell_reg[445] = inform_R[445][0];				r_cell_reg[446] = inform_R[446][0];				r_cell_reg[447] = inform_R[447][0];				r_cell_reg[448] = inform_R[448][0];				r_cell_reg[449] = inform_R[449][0];				r_cell_reg[450] = inform_R[450][0];				r_cell_reg[451] = inform_R[451][0];				r_cell_reg[452] = inform_R[452][0];				r_cell_reg[453] = inform_R[453][0];				r_cell_reg[454] = inform_R[454][0];				r_cell_reg[455] = inform_R[455][0];				r_cell_reg[456] = inform_R[456][0];				r_cell_reg[457] = inform_R[457][0];				r_cell_reg[458] = inform_R[458][0];				r_cell_reg[459] = inform_R[459][0];				r_cell_reg[460] = inform_R[460][0];				r_cell_reg[461] = inform_R[461][0];				r_cell_reg[462] = inform_R[462][0];				r_cell_reg[463] = inform_R[463][0];				r_cell_reg[464] = inform_R[464][0];				r_cell_reg[465] = inform_R[465][0];				r_cell_reg[466] = inform_R[466][0];				r_cell_reg[467] = inform_R[467][0];				r_cell_reg[468] = inform_R[468][0];				r_cell_reg[469] = inform_R[469][0];				r_cell_reg[470] = inform_R[470][0];				r_cell_reg[471] = inform_R[471][0];				r_cell_reg[472] = inform_R[472][0];				r_cell_reg[473] = inform_R[473][0];				r_cell_reg[474] = inform_R[474][0];				r_cell_reg[475] = inform_R[475][0];				r_cell_reg[476] = inform_R[476][0];				r_cell_reg[477] = inform_R[477][0];				r_cell_reg[478] = inform_R[478][0];				r_cell_reg[479] = inform_R[479][0];				r_cell_reg[480] = inform_R[480][0];				r_cell_reg[481] = inform_R[481][0];				r_cell_reg[482] = inform_R[482][0];				r_cell_reg[483] = inform_R[483][0];				r_cell_reg[484] = inform_R[484][0];				r_cell_reg[485] = inform_R[485][0];				r_cell_reg[486] = inform_R[486][0];				r_cell_reg[487] = inform_R[487][0];				r_cell_reg[488] = inform_R[488][0];				r_cell_reg[489] = inform_R[489][0];				r_cell_reg[490] = inform_R[490][0];				r_cell_reg[491] = inform_R[491][0];				r_cell_reg[492] = inform_R[492][0];				r_cell_reg[493] = inform_R[493][0];				r_cell_reg[494] = inform_R[494][0];				r_cell_reg[495] = inform_R[495][0];				r_cell_reg[496] = inform_R[496][0];				r_cell_reg[497] = inform_R[497][0];				r_cell_reg[498] = inform_R[498][0];				r_cell_reg[499] = inform_R[499][0];				r_cell_reg[500] = inform_R[500][0];				r_cell_reg[501] = inform_R[501][0];				r_cell_reg[502] = inform_R[502][0];				r_cell_reg[503] = inform_R[503][0];				r_cell_reg[504] = inform_R[504][0];				r_cell_reg[505] = inform_R[505][0];				r_cell_reg[506] = inform_R[506][0];				r_cell_reg[507] = inform_R[507][0];				r_cell_reg[508] = inform_R[508][0];				r_cell_reg[509] = inform_R[509][0];				r_cell_reg[510] = inform_R[510][0];				r_cell_reg[511] = inform_R[511][0];				r_cell_reg[512] = inform_R[512][0];				r_cell_reg[513] = inform_R[513][0];				r_cell_reg[514] = inform_R[514][0];				r_cell_reg[515] = inform_R[515][0];				r_cell_reg[516] = inform_R[516][0];				r_cell_reg[517] = inform_R[517][0];				r_cell_reg[518] = inform_R[518][0];				r_cell_reg[519] = inform_R[519][0];				r_cell_reg[520] = inform_R[520][0];				r_cell_reg[521] = inform_R[521][0];				r_cell_reg[522] = inform_R[522][0];				r_cell_reg[523] = inform_R[523][0];				r_cell_reg[524] = inform_R[524][0];				r_cell_reg[525] = inform_R[525][0];				r_cell_reg[526] = inform_R[526][0];				r_cell_reg[527] = inform_R[527][0];				r_cell_reg[528] = inform_R[528][0];				r_cell_reg[529] = inform_R[529][0];				r_cell_reg[530] = inform_R[530][0];				r_cell_reg[531] = inform_R[531][0];				r_cell_reg[532] = inform_R[532][0];				r_cell_reg[533] = inform_R[533][0];				r_cell_reg[534] = inform_R[534][0];				r_cell_reg[535] = inform_R[535][0];				r_cell_reg[536] = inform_R[536][0];				r_cell_reg[537] = inform_R[537][0];				r_cell_reg[538] = inform_R[538][0];				r_cell_reg[539] = inform_R[539][0];				r_cell_reg[540] = inform_R[540][0];				r_cell_reg[541] = inform_R[541][0];				r_cell_reg[542] = inform_R[542][0];				r_cell_reg[543] = inform_R[543][0];				r_cell_reg[544] = inform_R[544][0];				r_cell_reg[545] = inform_R[545][0];				r_cell_reg[546] = inform_R[546][0];				r_cell_reg[547] = inform_R[547][0];				r_cell_reg[548] = inform_R[548][0];				r_cell_reg[549] = inform_R[549][0];				r_cell_reg[550] = inform_R[550][0];				r_cell_reg[551] = inform_R[551][0];				r_cell_reg[552] = inform_R[552][0];				r_cell_reg[553] = inform_R[553][0];				r_cell_reg[554] = inform_R[554][0];				r_cell_reg[555] = inform_R[555][0];				r_cell_reg[556] = inform_R[556][0];				r_cell_reg[557] = inform_R[557][0];				r_cell_reg[558] = inform_R[558][0];				r_cell_reg[559] = inform_R[559][0];				r_cell_reg[560] = inform_R[560][0];				r_cell_reg[561] = inform_R[561][0];				r_cell_reg[562] = inform_R[562][0];				r_cell_reg[563] = inform_R[563][0];				r_cell_reg[564] = inform_R[564][0];				r_cell_reg[565] = inform_R[565][0];				r_cell_reg[566] = inform_R[566][0];				r_cell_reg[567] = inform_R[567][0];				r_cell_reg[568] = inform_R[568][0];				r_cell_reg[569] = inform_R[569][0];				r_cell_reg[570] = inform_R[570][0];				r_cell_reg[571] = inform_R[571][0];				r_cell_reg[572] = inform_R[572][0];				r_cell_reg[573] = inform_R[573][0];				r_cell_reg[574] = inform_R[574][0];				r_cell_reg[575] = inform_R[575][0];				r_cell_reg[576] = inform_R[576][0];				r_cell_reg[577] = inform_R[577][0];				r_cell_reg[578] = inform_R[578][0];				r_cell_reg[579] = inform_R[579][0];				r_cell_reg[580] = inform_R[580][0];				r_cell_reg[581] = inform_R[581][0];				r_cell_reg[582] = inform_R[582][0];				r_cell_reg[583] = inform_R[583][0];				r_cell_reg[584] = inform_R[584][0];				r_cell_reg[585] = inform_R[585][0];				r_cell_reg[586] = inform_R[586][0];				r_cell_reg[587] = inform_R[587][0];				r_cell_reg[588] = inform_R[588][0];				r_cell_reg[589] = inform_R[589][0];				r_cell_reg[590] = inform_R[590][0];				r_cell_reg[591] = inform_R[591][0];				r_cell_reg[592] = inform_R[592][0];				r_cell_reg[593] = inform_R[593][0];				r_cell_reg[594] = inform_R[594][0];				r_cell_reg[595] = inform_R[595][0];				r_cell_reg[596] = inform_R[596][0];				r_cell_reg[597] = inform_R[597][0];				r_cell_reg[598] = inform_R[598][0];				r_cell_reg[599] = inform_R[599][0];				r_cell_reg[600] = inform_R[600][0];				r_cell_reg[601] = inform_R[601][0];				r_cell_reg[602] = inform_R[602][0];				r_cell_reg[603] = inform_R[603][0];				r_cell_reg[604] = inform_R[604][0];				r_cell_reg[605] = inform_R[605][0];				r_cell_reg[606] = inform_R[606][0];				r_cell_reg[607] = inform_R[607][0];				r_cell_reg[608] = inform_R[608][0];				r_cell_reg[609] = inform_R[609][0];				r_cell_reg[610] = inform_R[610][0];				r_cell_reg[611] = inform_R[611][0];				r_cell_reg[612] = inform_R[612][0];				r_cell_reg[613] = inform_R[613][0];				r_cell_reg[614] = inform_R[614][0];				r_cell_reg[615] = inform_R[615][0];				r_cell_reg[616] = inform_R[616][0];				r_cell_reg[617] = inform_R[617][0];				r_cell_reg[618] = inform_R[618][0];				r_cell_reg[619] = inform_R[619][0];				r_cell_reg[620] = inform_R[620][0];				r_cell_reg[621] = inform_R[621][0];				r_cell_reg[622] = inform_R[622][0];				r_cell_reg[623] = inform_R[623][0];				r_cell_reg[624] = inform_R[624][0];				r_cell_reg[625] = inform_R[625][0];				r_cell_reg[626] = inform_R[626][0];				r_cell_reg[627] = inform_R[627][0];				r_cell_reg[628] = inform_R[628][0];				r_cell_reg[629] = inform_R[629][0];				r_cell_reg[630] = inform_R[630][0];				r_cell_reg[631] = inform_R[631][0];				r_cell_reg[632] = inform_R[632][0];				r_cell_reg[633] = inform_R[633][0];				r_cell_reg[634] = inform_R[634][0];				r_cell_reg[635] = inform_R[635][0];				r_cell_reg[636] = inform_R[636][0];				r_cell_reg[637] = inform_R[637][0];				r_cell_reg[638] = inform_R[638][0];				r_cell_reg[639] = inform_R[639][0];				r_cell_reg[640] = inform_R[640][0];				r_cell_reg[641] = inform_R[641][0];				r_cell_reg[642] = inform_R[642][0];				r_cell_reg[643] = inform_R[643][0];				r_cell_reg[644] = inform_R[644][0];				r_cell_reg[645] = inform_R[645][0];				r_cell_reg[646] = inform_R[646][0];				r_cell_reg[647] = inform_R[647][0];				r_cell_reg[648] = inform_R[648][0];				r_cell_reg[649] = inform_R[649][0];				r_cell_reg[650] = inform_R[650][0];				r_cell_reg[651] = inform_R[651][0];				r_cell_reg[652] = inform_R[652][0];				r_cell_reg[653] = inform_R[653][0];				r_cell_reg[654] = inform_R[654][0];				r_cell_reg[655] = inform_R[655][0];				r_cell_reg[656] = inform_R[656][0];				r_cell_reg[657] = inform_R[657][0];				r_cell_reg[658] = inform_R[658][0];				r_cell_reg[659] = inform_R[659][0];				r_cell_reg[660] = inform_R[660][0];				r_cell_reg[661] = inform_R[661][0];				r_cell_reg[662] = inform_R[662][0];				r_cell_reg[663] = inform_R[663][0];				r_cell_reg[664] = inform_R[664][0];				r_cell_reg[665] = inform_R[665][0];				r_cell_reg[666] = inform_R[666][0];				r_cell_reg[667] = inform_R[667][0];				r_cell_reg[668] = inform_R[668][0];				r_cell_reg[669] = inform_R[669][0];				r_cell_reg[670] = inform_R[670][0];				r_cell_reg[671] = inform_R[671][0];				r_cell_reg[672] = inform_R[672][0];				r_cell_reg[673] = inform_R[673][0];				r_cell_reg[674] = inform_R[674][0];				r_cell_reg[675] = inform_R[675][0];				r_cell_reg[676] = inform_R[676][0];				r_cell_reg[677] = inform_R[677][0];				r_cell_reg[678] = inform_R[678][0];				r_cell_reg[679] = inform_R[679][0];				r_cell_reg[680] = inform_R[680][0];				r_cell_reg[681] = inform_R[681][0];				r_cell_reg[682] = inform_R[682][0];				r_cell_reg[683] = inform_R[683][0];				r_cell_reg[684] = inform_R[684][0];				r_cell_reg[685] = inform_R[685][0];				r_cell_reg[686] = inform_R[686][0];				r_cell_reg[687] = inform_R[687][0];				r_cell_reg[688] = inform_R[688][0];				r_cell_reg[689] = inform_R[689][0];				r_cell_reg[690] = inform_R[690][0];				r_cell_reg[691] = inform_R[691][0];				r_cell_reg[692] = inform_R[692][0];				r_cell_reg[693] = inform_R[693][0];				r_cell_reg[694] = inform_R[694][0];				r_cell_reg[695] = inform_R[695][0];				r_cell_reg[696] = inform_R[696][0];				r_cell_reg[697] = inform_R[697][0];				r_cell_reg[698] = inform_R[698][0];				r_cell_reg[699] = inform_R[699][0];				r_cell_reg[700] = inform_R[700][0];				r_cell_reg[701] = inform_R[701][0];				r_cell_reg[702] = inform_R[702][0];				r_cell_reg[703] = inform_R[703][0];				r_cell_reg[704] = inform_R[704][0];				r_cell_reg[705] = inform_R[705][0];				r_cell_reg[706] = inform_R[706][0];				r_cell_reg[707] = inform_R[707][0];				r_cell_reg[708] = inform_R[708][0];				r_cell_reg[709] = inform_R[709][0];				r_cell_reg[710] = inform_R[710][0];				r_cell_reg[711] = inform_R[711][0];				r_cell_reg[712] = inform_R[712][0];				r_cell_reg[713] = inform_R[713][0];				r_cell_reg[714] = inform_R[714][0];				r_cell_reg[715] = inform_R[715][0];				r_cell_reg[716] = inform_R[716][0];				r_cell_reg[717] = inform_R[717][0];				r_cell_reg[718] = inform_R[718][0];				r_cell_reg[719] = inform_R[719][0];				r_cell_reg[720] = inform_R[720][0];				r_cell_reg[721] = inform_R[721][0];				r_cell_reg[722] = inform_R[722][0];				r_cell_reg[723] = inform_R[723][0];				r_cell_reg[724] = inform_R[724][0];				r_cell_reg[725] = inform_R[725][0];				r_cell_reg[726] = inform_R[726][0];				r_cell_reg[727] = inform_R[727][0];				r_cell_reg[728] = inform_R[728][0];				r_cell_reg[729] = inform_R[729][0];				r_cell_reg[730] = inform_R[730][0];				r_cell_reg[731] = inform_R[731][0];				r_cell_reg[732] = inform_R[732][0];				r_cell_reg[733] = inform_R[733][0];				r_cell_reg[734] = inform_R[734][0];				r_cell_reg[735] = inform_R[735][0];				r_cell_reg[736] = inform_R[736][0];				r_cell_reg[737] = inform_R[737][0];				r_cell_reg[738] = inform_R[738][0];				r_cell_reg[739] = inform_R[739][0];				r_cell_reg[740] = inform_R[740][0];				r_cell_reg[741] = inform_R[741][0];				r_cell_reg[742] = inform_R[742][0];				r_cell_reg[743] = inform_R[743][0];				r_cell_reg[744] = inform_R[744][0];				r_cell_reg[745] = inform_R[745][0];				r_cell_reg[746] = inform_R[746][0];				r_cell_reg[747] = inform_R[747][0];				r_cell_reg[748] = inform_R[748][0];				r_cell_reg[749] = inform_R[749][0];				r_cell_reg[750] = inform_R[750][0];				r_cell_reg[751] = inform_R[751][0];				r_cell_reg[752] = inform_R[752][0];				r_cell_reg[753] = inform_R[753][0];				r_cell_reg[754] = inform_R[754][0];				r_cell_reg[755] = inform_R[755][0];				r_cell_reg[756] = inform_R[756][0];				r_cell_reg[757] = inform_R[757][0];				r_cell_reg[758] = inform_R[758][0];				r_cell_reg[759] = inform_R[759][0];				r_cell_reg[760] = inform_R[760][0];				r_cell_reg[761] = inform_R[761][0];				r_cell_reg[762] = inform_R[762][0];				r_cell_reg[763] = inform_R[763][0];				r_cell_reg[764] = inform_R[764][0];				r_cell_reg[765] = inform_R[765][0];				r_cell_reg[766] = inform_R[766][0];				r_cell_reg[767] = inform_R[767][0];				r_cell_reg[768] = inform_R[768][0];				r_cell_reg[769] = inform_R[769][0];				r_cell_reg[770] = inform_R[770][0];				r_cell_reg[771] = inform_R[771][0];				r_cell_reg[772] = inform_R[772][0];				r_cell_reg[773] = inform_R[773][0];				r_cell_reg[774] = inform_R[774][0];				r_cell_reg[775] = inform_R[775][0];				r_cell_reg[776] = inform_R[776][0];				r_cell_reg[777] = inform_R[777][0];				r_cell_reg[778] = inform_R[778][0];				r_cell_reg[779] = inform_R[779][0];				r_cell_reg[780] = inform_R[780][0];				r_cell_reg[781] = inform_R[781][0];				r_cell_reg[782] = inform_R[782][0];				r_cell_reg[783] = inform_R[783][0];				r_cell_reg[784] = inform_R[784][0];				r_cell_reg[785] = inform_R[785][0];				r_cell_reg[786] = inform_R[786][0];				r_cell_reg[787] = inform_R[787][0];				r_cell_reg[788] = inform_R[788][0];				r_cell_reg[789] = inform_R[789][0];				r_cell_reg[790] = inform_R[790][0];				r_cell_reg[791] = inform_R[791][0];				r_cell_reg[792] = inform_R[792][0];				r_cell_reg[793] = inform_R[793][0];				r_cell_reg[794] = inform_R[794][0];				r_cell_reg[795] = inform_R[795][0];				r_cell_reg[796] = inform_R[796][0];				r_cell_reg[797] = inform_R[797][0];				r_cell_reg[798] = inform_R[798][0];				r_cell_reg[799] = inform_R[799][0];				r_cell_reg[800] = inform_R[800][0];				r_cell_reg[801] = inform_R[801][0];				r_cell_reg[802] = inform_R[802][0];				r_cell_reg[803] = inform_R[803][0];				r_cell_reg[804] = inform_R[804][0];				r_cell_reg[805] = inform_R[805][0];				r_cell_reg[806] = inform_R[806][0];				r_cell_reg[807] = inform_R[807][0];				r_cell_reg[808] = inform_R[808][0];				r_cell_reg[809] = inform_R[809][0];				r_cell_reg[810] = inform_R[810][0];				r_cell_reg[811] = inform_R[811][0];				r_cell_reg[812] = inform_R[812][0];				r_cell_reg[813] = inform_R[813][0];				r_cell_reg[814] = inform_R[814][0];				r_cell_reg[815] = inform_R[815][0];				r_cell_reg[816] = inform_R[816][0];				r_cell_reg[817] = inform_R[817][0];				r_cell_reg[818] = inform_R[818][0];				r_cell_reg[819] = inform_R[819][0];				r_cell_reg[820] = inform_R[820][0];				r_cell_reg[821] = inform_R[821][0];				r_cell_reg[822] = inform_R[822][0];				r_cell_reg[823] = inform_R[823][0];				r_cell_reg[824] = inform_R[824][0];				r_cell_reg[825] = inform_R[825][0];				r_cell_reg[826] = inform_R[826][0];				r_cell_reg[827] = inform_R[827][0];				r_cell_reg[828] = inform_R[828][0];				r_cell_reg[829] = inform_R[829][0];				r_cell_reg[830] = inform_R[830][0];				r_cell_reg[831] = inform_R[831][0];				r_cell_reg[832] = inform_R[832][0];				r_cell_reg[833] = inform_R[833][0];				r_cell_reg[834] = inform_R[834][0];				r_cell_reg[835] = inform_R[835][0];				r_cell_reg[836] = inform_R[836][0];				r_cell_reg[837] = inform_R[837][0];				r_cell_reg[838] = inform_R[838][0];				r_cell_reg[839] = inform_R[839][0];				r_cell_reg[840] = inform_R[840][0];				r_cell_reg[841] = inform_R[841][0];				r_cell_reg[842] = inform_R[842][0];				r_cell_reg[843] = inform_R[843][0];				r_cell_reg[844] = inform_R[844][0];				r_cell_reg[845] = inform_R[845][0];				r_cell_reg[846] = inform_R[846][0];				r_cell_reg[847] = inform_R[847][0];				r_cell_reg[848] = inform_R[848][0];				r_cell_reg[849] = inform_R[849][0];				r_cell_reg[850] = inform_R[850][0];				r_cell_reg[851] = inform_R[851][0];				r_cell_reg[852] = inform_R[852][0];				r_cell_reg[853] = inform_R[853][0];				r_cell_reg[854] = inform_R[854][0];				r_cell_reg[855] = inform_R[855][0];				r_cell_reg[856] = inform_R[856][0];				r_cell_reg[857] = inform_R[857][0];				r_cell_reg[858] = inform_R[858][0];				r_cell_reg[859] = inform_R[859][0];				r_cell_reg[860] = inform_R[860][0];				r_cell_reg[861] = inform_R[861][0];				r_cell_reg[862] = inform_R[862][0];				r_cell_reg[863] = inform_R[863][0];				r_cell_reg[864] = inform_R[864][0];				r_cell_reg[865] = inform_R[865][0];				r_cell_reg[866] = inform_R[866][0];				r_cell_reg[867] = inform_R[867][0];				r_cell_reg[868] = inform_R[868][0];				r_cell_reg[869] = inform_R[869][0];				r_cell_reg[870] = inform_R[870][0];				r_cell_reg[871] = inform_R[871][0];				r_cell_reg[872] = inform_R[872][0];				r_cell_reg[873] = inform_R[873][0];				r_cell_reg[874] = inform_R[874][0];				r_cell_reg[875] = inform_R[875][0];				r_cell_reg[876] = inform_R[876][0];				r_cell_reg[877] = inform_R[877][0];				r_cell_reg[878] = inform_R[878][0];				r_cell_reg[879] = inform_R[879][0];				r_cell_reg[880] = inform_R[880][0];				r_cell_reg[881] = inform_R[881][0];				r_cell_reg[882] = inform_R[882][0];				r_cell_reg[883] = inform_R[883][0];				r_cell_reg[884] = inform_R[884][0];				r_cell_reg[885] = inform_R[885][0];				r_cell_reg[886] = inform_R[886][0];				r_cell_reg[887] = inform_R[887][0];				r_cell_reg[888] = inform_R[888][0];				r_cell_reg[889] = inform_R[889][0];				r_cell_reg[890] = inform_R[890][0];				r_cell_reg[891] = inform_R[891][0];				r_cell_reg[892] = inform_R[892][0];				r_cell_reg[893] = inform_R[893][0];				r_cell_reg[894] = inform_R[894][0];				r_cell_reg[895] = inform_R[895][0];				r_cell_reg[896] = inform_R[896][0];				r_cell_reg[897] = inform_R[897][0];				r_cell_reg[898] = inform_R[898][0];				r_cell_reg[899] = inform_R[899][0];				r_cell_reg[900] = inform_R[900][0];				r_cell_reg[901] = inform_R[901][0];				r_cell_reg[902] = inform_R[902][0];				r_cell_reg[903] = inform_R[903][0];				r_cell_reg[904] = inform_R[904][0];				r_cell_reg[905] = inform_R[905][0];				r_cell_reg[906] = inform_R[906][0];				r_cell_reg[907] = inform_R[907][0];				r_cell_reg[908] = inform_R[908][0];				r_cell_reg[909] = inform_R[909][0];				r_cell_reg[910] = inform_R[910][0];				r_cell_reg[911] = inform_R[911][0];				r_cell_reg[912] = inform_R[912][0];				r_cell_reg[913] = inform_R[913][0];				r_cell_reg[914] = inform_R[914][0];				r_cell_reg[915] = inform_R[915][0];				r_cell_reg[916] = inform_R[916][0];				r_cell_reg[917] = inform_R[917][0];				r_cell_reg[918] = inform_R[918][0];				r_cell_reg[919] = inform_R[919][0];				r_cell_reg[920] = inform_R[920][0];				r_cell_reg[921] = inform_R[921][0];				r_cell_reg[922] = inform_R[922][0];				r_cell_reg[923] = inform_R[923][0];				r_cell_reg[924] = inform_R[924][0];				r_cell_reg[925] = inform_R[925][0];				r_cell_reg[926] = inform_R[926][0];				r_cell_reg[927] = inform_R[927][0];				r_cell_reg[928] = inform_R[928][0];				r_cell_reg[929] = inform_R[929][0];				r_cell_reg[930] = inform_R[930][0];				r_cell_reg[931] = inform_R[931][0];				r_cell_reg[932] = inform_R[932][0];				r_cell_reg[933] = inform_R[933][0];				r_cell_reg[934] = inform_R[934][0];				r_cell_reg[935] = inform_R[935][0];				r_cell_reg[936] = inform_R[936][0];				r_cell_reg[937] = inform_R[937][0];				r_cell_reg[938] = inform_R[938][0];				r_cell_reg[939] = inform_R[939][0];				r_cell_reg[940] = inform_R[940][0];				r_cell_reg[941] = inform_R[941][0];				r_cell_reg[942] = inform_R[942][0];				r_cell_reg[943] = inform_R[943][0];				r_cell_reg[944] = inform_R[944][0];				r_cell_reg[945] = inform_R[945][0];				r_cell_reg[946] = inform_R[946][0];				r_cell_reg[947] = inform_R[947][0];				r_cell_reg[948] = inform_R[948][0];				r_cell_reg[949] = inform_R[949][0];				r_cell_reg[950] = inform_R[950][0];				r_cell_reg[951] = inform_R[951][0];				r_cell_reg[952] = inform_R[952][0];				r_cell_reg[953] = inform_R[953][0];				r_cell_reg[954] = inform_R[954][0];				r_cell_reg[955] = inform_R[955][0];				r_cell_reg[956] = inform_R[956][0];				r_cell_reg[957] = inform_R[957][0];				r_cell_reg[958] = inform_R[958][0];				r_cell_reg[959] = inform_R[959][0];				r_cell_reg[960] = inform_R[960][0];				r_cell_reg[961] = inform_R[961][0];				r_cell_reg[962] = inform_R[962][0];				r_cell_reg[963] = inform_R[963][0];				r_cell_reg[964] = inform_R[964][0];				r_cell_reg[965] = inform_R[965][0];				r_cell_reg[966] = inform_R[966][0];				r_cell_reg[967] = inform_R[967][0];				r_cell_reg[968] = inform_R[968][0];				r_cell_reg[969] = inform_R[969][0];				r_cell_reg[970] = inform_R[970][0];				r_cell_reg[971] = inform_R[971][0];				r_cell_reg[972] = inform_R[972][0];				r_cell_reg[973] = inform_R[973][0];				r_cell_reg[974] = inform_R[974][0];				r_cell_reg[975] = inform_R[975][0];				r_cell_reg[976] = inform_R[976][0];				r_cell_reg[977] = inform_R[977][0];				r_cell_reg[978] = inform_R[978][0];				r_cell_reg[979] = inform_R[979][0];				r_cell_reg[980] = inform_R[980][0];				r_cell_reg[981] = inform_R[981][0];				r_cell_reg[982] = inform_R[982][0];				r_cell_reg[983] = inform_R[983][0];				r_cell_reg[984] = inform_R[984][0];				r_cell_reg[985] = inform_R[985][0];				r_cell_reg[986] = inform_R[986][0];				r_cell_reg[987] = inform_R[987][0];				r_cell_reg[988] = inform_R[988][0];				r_cell_reg[989] = inform_R[989][0];				r_cell_reg[990] = inform_R[990][0];				r_cell_reg[991] = inform_R[991][0];				r_cell_reg[992] = inform_R[992][0];				r_cell_reg[993] = inform_R[993][0];				r_cell_reg[994] = inform_R[994][0];				r_cell_reg[995] = inform_R[995][0];				r_cell_reg[996] = inform_R[996][0];				r_cell_reg[997] = inform_R[997][0];				r_cell_reg[998] = inform_R[998][0];				r_cell_reg[999] = inform_R[999][0];				r_cell_reg[1000] = inform_R[1000][0];				r_cell_reg[1001] = inform_R[1001][0];				r_cell_reg[1002] = inform_R[1002][0];				r_cell_reg[1003] = inform_R[1003][0];				r_cell_reg[1004] = inform_R[1004][0];				r_cell_reg[1005] = inform_R[1005][0];				r_cell_reg[1006] = inform_R[1006][0];				r_cell_reg[1007] = inform_R[1007][0];				r_cell_reg[1008] = inform_R[1008][0];				r_cell_reg[1009] = inform_R[1009][0];				r_cell_reg[1010] = inform_R[1010][0];				r_cell_reg[1011] = inform_R[1011][0];				r_cell_reg[1012] = inform_R[1012][0];				r_cell_reg[1013] = inform_R[1013][0];				r_cell_reg[1014] = inform_R[1014][0];				r_cell_reg[1015] = inform_R[1015][0];				r_cell_reg[1016] = inform_R[1016][0];				r_cell_reg[1017] = inform_R[1017][0];				r_cell_reg[1018] = inform_R[1018][0];				r_cell_reg[1019] = inform_R[1019][0];				r_cell_reg[1020] = inform_R[1020][0];				r_cell_reg[1021] = inform_R[1021][0];				r_cell_reg[1022] = inform_R[1022][0];				r_cell_reg[1023] = inform_R[1023][0];				l_cell_reg[0] = inform_L[0][1];				l_cell_reg[1] = inform_L[1][1];				l_cell_reg[2] = inform_L[2][1];				l_cell_reg[3] = inform_L[3][1];				l_cell_reg[4] = inform_L[4][1];				l_cell_reg[5] = inform_L[5][1];				l_cell_reg[6] = inform_L[6][1];				l_cell_reg[7] = inform_L[7][1];				l_cell_reg[8] = inform_L[8][1];				l_cell_reg[9] = inform_L[9][1];				l_cell_reg[10] = inform_L[10][1];				l_cell_reg[11] = inform_L[11][1];				l_cell_reg[12] = inform_L[12][1];				l_cell_reg[13] = inform_L[13][1];				l_cell_reg[14] = inform_L[14][1];				l_cell_reg[15] = inform_L[15][1];				l_cell_reg[16] = inform_L[16][1];				l_cell_reg[17] = inform_L[17][1];				l_cell_reg[18] = inform_L[18][1];				l_cell_reg[19] = inform_L[19][1];				l_cell_reg[20] = inform_L[20][1];				l_cell_reg[21] = inform_L[21][1];				l_cell_reg[22] = inform_L[22][1];				l_cell_reg[23] = inform_L[23][1];				l_cell_reg[24] = inform_L[24][1];				l_cell_reg[25] = inform_L[25][1];				l_cell_reg[26] = inform_L[26][1];				l_cell_reg[27] = inform_L[27][1];				l_cell_reg[28] = inform_L[28][1];				l_cell_reg[29] = inform_L[29][1];				l_cell_reg[30] = inform_L[30][1];				l_cell_reg[31] = inform_L[31][1];				l_cell_reg[32] = inform_L[32][1];				l_cell_reg[33] = inform_L[33][1];				l_cell_reg[34] = inform_L[34][1];				l_cell_reg[35] = inform_L[35][1];				l_cell_reg[36] = inform_L[36][1];				l_cell_reg[37] = inform_L[37][1];				l_cell_reg[38] = inform_L[38][1];				l_cell_reg[39] = inform_L[39][1];				l_cell_reg[40] = inform_L[40][1];				l_cell_reg[41] = inform_L[41][1];				l_cell_reg[42] = inform_L[42][1];				l_cell_reg[43] = inform_L[43][1];				l_cell_reg[44] = inform_L[44][1];				l_cell_reg[45] = inform_L[45][1];				l_cell_reg[46] = inform_L[46][1];				l_cell_reg[47] = inform_L[47][1];				l_cell_reg[48] = inform_L[48][1];				l_cell_reg[49] = inform_L[49][1];				l_cell_reg[50] = inform_L[50][1];				l_cell_reg[51] = inform_L[51][1];				l_cell_reg[52] = inform_L[52][1];				l_cell_reg[53] = inform_L[53][1];				l_cell_reg[54] = inform_L[54][1];				l_cell_reg[55] = inform_L[55][1];				l_cell_reg[56] = inform_L[56][1];				l_cell_reg[57] = inform_L[57][1];				l_cell_reg[58] = inform_L[58][1];				l_cell_reg[59] = inform_L[59][1];				l_cell_reg[60] = inform_L[60][1];				l_cell_reg[61] = inform_L[61][1];				l_cell_reg[62] = inform_L[62][1];				l_cell_reg[63] = inform_L[63][1];				l_cell_reg[64] = inform_L[64][1];				l_cell_reg[65] = inform_L[65][1];				l_cell_reg[66] = inform_L[66][1];				l_cell_reg[67] = inform_L[67][1];				l_cell_reg[68] = inform_L[68][1];				l_cell_reg[69] = inform_L[69][1];				l_cell_reg[70] = inform_L[70][1];				l_cell_reg[71] = inform_L[71][1];				l_cell_reg[72] = inform_L[72][1];				l_cell_reg[73] = inform_L[73][1];				l_cell_reg[74] = inform_L[74][1];				l_cell_reg[75] = inform_L[75][1];				l_cell_reg[76] = inform_L[76][1];				l_cell_reg[77] = inform_L[77][1];				l_cell_reg[78] = inform_L[78][1];				l_cell_reg[79] = inform_L[79][1];				l_cell_reg[80] = inform_L[80][1];				l_cell_reg[81] = inform_L[81][1];				l_cell_reg[82] = inform_L[82][1];				l_cell_reg[83] = inform_L[83][1];				l_cell_reg[84] = inform_L[84][1];				l_cell_reg[85] = inform_L[85][1];				l_cell_reg[86] = inform_L[86][1];				l_cell_reg[87] = inform_L[87][1];				l_cell_reg[88] = inform_L[88][1];				l_cell_reg[89] = inform_L[89][1];				l_cell_reg[90] = inform_L[90][1];				l_cell_reg[91] = inform_L[91][1];				l_cell_reg[92] = inform_L[92][1];				l_cell_reg[93] = inform_L[93][1];				l_cell_reg[94] = inform_L[94][1];				l_cell_reg[95] = inform_L[95][1];				l_cell_reg[96] = inform_L[96][1];				l_cell_reg[97] = inform_L[97][1];				l_cell_reg[98] = inform_L[98][1];				l_cell_reg[99] = inform_L[99][1];				l_cell_reg[100] = inform_L[100][1];				l_cell_reg[101] = inform_L[101][1];				l_cell_reg[102] = inform_L[102][1];				l_cell_reg[103] = inform_L[103][1];				l_cell_reg[104] = inform_L[104][1];				l_cell_reg[105] = inform_L[105][1];				l_cell_reg[106] = inform_L[106][1];				l_cell_reg[107] = inform_L[107][1];				l_cell_reg[108] = inform_L[108][1];				l_cell_reg[109] = inform_L[109][1];				l_cell_reg[110] = inform_L[110][1];				l_cell_reg[111] = inform_L[111][1];				l_cell_reg[112] = inform_L[112][1];				l_cell_reg[113] = inform_L[113][1];				l_cell_reg[114] = inform_L[114][1];				l_cell_reg[115] = inform_L[115][1];				l_cell_reg[116] = inform_L[116][1];				l_cell_reg[117] = inform_L[117][1];				l_cell_reg[118] = inform_L[118][1];				l_cell_reg[119] = inform_L[119][1];				l_cell_reg[120] = inform_L[120][1];				l_cell_reg[121] = inform_L[121][1];				l_cell_reg[122] = inform_L[122][1];				l_cell_reg[123] = inform_L[123][1];				l_cell_reg[124] = inform_L[124][1];				l_cell_reg[125] = inform_L[125][1];				l_cell_reg[126] = inform_L[126][1];				l_cell_reg[127] = inform_L[127][1];				l_cell_reg[128] = inform_L[128][1];				l_cell_reg[129] = inform_L[129][1];				l_cell_reg[130] = inform_L[130][1];				l_cell_reg[131] = inform_L[131][1];				l_cell_reg[132] = inform_L[132][1];				l_cell_reg[133] = inform_L[133][1];				l_cell_reg[134] = inform_L[134][1];				l_cell_reg[135] = inform_L[135][1];				l_cell_reg[136] = inform_L[136][1];				l_cell_reg[137] = inform_L[137][1];				l_cell_reg[138] = inform_L[138][1];				l_cell_reg[139] = inform_L[139][1];				l_cell_reg[140] = inform_L[140][1];				l_cell_reg[141] = inform_L[141][1];				l_cell_reg[142] = inform_L[142][1];				l_cell_reg[143] = inform_L[143][1];				l_cell_reg[144] = inform_L[144][1];				l_cell_reg[145] = inform_L[145][1];				l_cell_reg[146] = inform_L[146][1];				l_cell_reg[147] = inform_L[147][1];				l_cell_reg[148] = inform_L[148][1];				l_cell_reg[149] = inform_L[149][1];				l_cell_reg[150] = inform_L[150][1];				l_cell_reg[151] = inform_L[151][1];				l_cell_reg[152] = inform_L[152][1];				l_cell_reg[153] = inform_L[153][1];				l_cell_reg[154] = inform_L[154][1];				l_cell_reg[155] = inform_L[155][1];				l_cell_reg[156] = inform_L[156][1];				l_cell_reg[157] = inform_L[157][1];				l_cell_reg[158] = inform_L[158][1];				l_cell_reg[159] = inform_L[159][1];				l_cell_reg[160] = inform_L[160][1];				l_cell_reg[161] = inform_L[161][1];				l_cell_reg[162] = inform_L[162][1];				l_cell_reg[163] = inform_L[163][1];				l_cell_reg[164] = inform_L[164][1];				l_cell_reg[165] = inform_L[165][1];				l_cell_reg[166] = inform_L[166][1];				l_cell_reg[167] = inform_L[167][1];				l_cell_reg[168] = inform_L[168][1];				l_cell_reg[169] = inform_L[169][1];				l_cell_reg[170] = inform_L[170][1];				l_cell_reg[171] = inform_L[171][1];				l_cell_reg[172] = inform_L[172][1];				l_cell_reg[173] = inform_L[173][1];				l_cell_reg[174] = inform_L[174][1];				l_cell_reg[175] = inform_L[175][1];				l_cell_reg[176] = inform_L[176][1];				l_cell_reg[177] = inform_L[177][1];				l_cell_reg[178] = inform_L[178][1];				l_cell_reg[179] = inform_L[179][1];				l_cell_reg[180] = inform_L[180][1];				l_cell_reg[181] = inform_L[181][1];				l_cell_reg[182] = inform_L[182][1];				l_cell_reg[183] = inform_L[183][1];				l_cell_reg[184] = inform_L[184][1];				l_cell_reg[185] = inform_L[185][1];				l_cell_reg[186] = inform_L[186][1];				l_cell_reg[187] = inform_L[187][1];				l_cell_reg[188] = inform_L[188][1];				l_cell_reg[189] = inform_L[189][1];				l_cell_reg[190] = inform_L[190][1];				l_cell_reg[191] = inform_L[191][1];				l_cell_reg[192] = inform_L[192][1];				l_cell_reg[193] = inform_L[193][1];				l_cell_reg[194] = inform_L[194][1];				l_cell_reg[195] = inform_L[195][1];				l_cell_reg[196] = inform_L[196][1];				l_cell_reg[197] = inform_L[197][1];				l_cell_reg[198] = inform_L[198][1];				l_cell_reg[199] = inform_L[199][1];				l_cell_reg[200] = inform_L[200][1];				l_cell_reg[201] = inform_L[201][1];				l_cell_reg[202] = inform_L[202][1];				l_cell_reg[203] = inform_L[203][1];				l_cell_reg[204] = inform_L[204][1];				l_cell_reg[205] = inform_L[205][1];				l_cell_reg[206] = inform_L[206][1];				l_cell_reg[207] = inform_L[207][1];				l_cell_reg[208] = inform_L[208][1];				l_cell_reg[209] = inform_L[209][1];				l_cell_reg[210] = inform_L[210][1];				l_cell_reg[211] = inform_L[211][1];				l_cell_reg[212] = inform_L[212][1];				l_cell_reg[213] = inform_L[213][1];				l_cell_reg[214] = inform_L[214][1];				l_cell_reg[215] = inform_L[215][1];				l_cell_reg[216] = inform_L[216][1];				l_cell_reg[217] = inform_L[217][1];				l_cell_reg[218] = inform_L[218][1];				l_cell_reg[219] = inform_L[219][1];				l_cell_reg[220] = inform_L[220][1];				l_cell_reg[221] = inform_L[221][1];				l_cell_reg[222] = inform_L[222][1];				l_cell_reg[223] = inform_L[223][1];				l_cell_reg[224] = inform_L[224][1];				l_cell_reg[225] = inform_L[225][1];				l_cell_reg[226] = inform_L[226][1];				l_cell_reg[227] = inform_L[227][1];				l_cell_reg[228] = inform_L[228][1];				l_cell_reg[229] = inform_L[229][1];				l_cell_reg[230] = inform_L[230][1];				l_cell_reg[231] = inform_L[231][1];				l_cell_reg[232] = inform_L[232][1];				l_cell_reg[233] = inform_L[233][1];				l_cell_reg[234] = inform_L[234][1];				l_cell_reg[235] = inform_L[235][1];				l_cell_reg[236] = inform_L[236][1];				l_cell_reg[237] = inform_L[237][1];				l_cell_reg[238] = inform_L[238][1];				l_cell_reg[239] = inform_L[239][1];				l_cell_reg[240] = inform_L[240][1];				l_cell_reg[241] = inform_L[241][1];				l_cell_reg[242] = inform_L[242][1];				l_cell_reg[243] = inform_L[243][1];				l_cell_reg[244] = inform_L[244][1];				l_cell_reg[245] = inform_L[245][1];				l_cell_reg[246] = inform_L[246][1];				l_cell_reg[247] = inform_L[247][1];				l_cell_reg[248] = inform_L[248][1];				l_cell_reg[249] = inform_L[249][1];				l_cell_reg[250] = inform_L[250][1];				l_cell_reg[251] = inform_L[251][1];				l_cell_reg[252] = inform_L[252][1];				l_cell_reg[253] = inform_L[253][1];				l_cell_reg[254] = inform_L[254][1];				l_cell_reg[255] = inform_L[255][1];				l_cell_reg[256] = inform_L[256][1];				l_cell_reg[257] = inform_L[257][1];				l_cell_reg[258] = inform_L[258][1];				l_cell_reg[259] = inform_L[259][1];				l_cell_reg[260] = inform_L[260][1];				l_cell_reg[261] = inform_L[261][1];				l_cell_reg[262] = inform_L[262][1];				l_cell_reg[263] = inform_L[263][1];				l_cell_reg[264] = inform_L[264][1];				l_cell_reg[265] = inform_L[265][1];				l_cell_reg[266] = inform_L[266][1];				l_cell_reg[267] = inform_L[267][1];				l_cell_reg[268] = inform_L[268][1];				l_cell_reg[269] = inform_L[269][1];				l_cell_reg[270] = inform_L[270][1];				l_cell_reg[271] = inform_L[271][1];				l_cell_reg[272] = inform_L[272][1];				l_cell_reg[273] = inform_L[273][1];				l_cell_reg[274] = inform_L[274][1];				l_cell_reg[275] = inform_L[275][1];				l_cell_reg[276] = inform_L[276][1];				l_cell_reg[277] = inform_L[277][1];				l_cell_reg[278] = inform_L[278][1];				l_cell_reg[279] = inform_L[279][1];				l_cell_reg[280] = inform_L[280][1];				l_cell_reg[281] = inform_L[281][1];				l_cell_reg[282] = inform_L[282][1];				l_cell_reg[283] = inform_L[283][1];				l_cell_reg[284] = inform_L[284][1];				l_cell_reg[285] = inform_L[285][1];				l_cell_reg[286] = inform_L[286][1];				l_cell_reg[287] = inform_L[287][1];				l_cell_reg[288] = inform_L[288][1];				l_cell_reg[289] = inform_L[289][1];				l_cell_reg[290] = inform_L[290][1];				l_cell_reg[291] = inform_L[291][1];				l_cell_reg[292] = inform_L[292][1];				l_cell_reg[293] = inform_L[293][1];				l_cell_reg[294] = inform_L[294][1];				l_cell_reg[295] = inform_L[295][1];				l_cell_reg[296] = inform_L[296][1];				l_cell_reg[297] = inform_L[297][1];				l_cell_reg[298] = inform_L[298][1];				l_cell_reg[299] = inform_L[299][1];				l_cell_reg[300] = inform_L[300][1];				l_cell_reg[301] = inform_L[301][1];				l_cell_reg[302] = inform_L[302][1];				l_cell_reg[303] = inform_L[303][1];				l_cell_reg[304] = inform_L[304][1];				l_cell_reg[305] = inform_L[305][1];				l_cell_reg[306] = inform_L[306][1];				l_cell_reg[307] = inform_L[307][1];				l_cell_reg[308] = inform_L[308][1];				l_cell_reg[309] = inform_L[309][1];				l_cell_reg[310] = inform_L[310][1];				l_cell_reg[311] = inform_L[311][1];				l_cell_reg[312] = inform_L[312][1];				l_cell_reg[313] = inform_L[313][1];				l_cell_reg[314] = inform_L[314][1];				l_cell_reg[315] = inform_L[315][1];				l_cell_reg[316] = inform_L[316][1];				l_cell_reg[317] = inform_L[317][1];				l_cell_reg[318] = inform_L[318][1];				l_cell_reg[319] = inform_L[319][1];				l_cell_reg[320] = inform_L[320][1];				l_cell_reg[321] = inform_L[321][1];				l_cell_reg[322] = inform_L[322][1];				l_cell_reg[323] = inform_L[323][1];				l_cell_reg[324] = inform_L[324][1];				l_cell_reg[325] = inform_L[325][1];				l_cell_reg[326] = inform_L[326][1];				l_cell_reg[327] = inform_L[327][1];				l_cell_reg[328] = inform_L[328][1];				l_cell_reg[329] = inform_L[329][1];				l_cell_reg[330] = inform_L[330][1];				l_cell_reg[331] = inform_L[331][1];				l_cell_reg[332] = inform_L[332][1];				l_cell_reg[333] = inform_L[333][1];				l_cell_reg[334] = inform_L[334][1];				l_cell_reg[335] = inform_L[335][1];				l_cell_reg[336] = inform_L[336][1];				l_cell_reg[337] = inform_L[337][1];				l_cell_reg[338] = inform_L[338][1];				l_cell_reg[339] = inform_L[339][1];				l_cell_reg[340] = inform_L[340][1];				l_cell_reg[341] = inform_L[341][1];				l_cell_reg[342] = inform_L[342][1];				l_cell_reg[343] = inform_L[343][1];				l_cell_reg[344] = inform_L[344][1];				l_cell_reg[345] = inform_L[345][1];				l_cell_reg[346] = inform_L[346][1];				l_cell_reg[347] = inform_L[347][1];				l_cell_reg[348] = inform_L[348][1];				l_cell_reg[349] = inform_L[349][1];				l_cell_reg[350] = inform_L[350][1];				l_cell_reg[351] = inform_L[351][1];				l_cell_reg[352] = inform_L[352][1];				l_cell_reg[353] = inform_L[353][1];				l_cell_reg[354] = inform_L[354][1];				l_cell_reg[355] = inform_L[355][1];				l_cell_reg[356] = inform_L[356][1];				l_cell_reg[357] = inform_L[357][1];				l_cell_reg[358] = inform_L[358][1];				l_cell_reg[359] = inform_L[359][1];				l_cell_reg[360] = inform_L[360][1];				l_cell_reg[361] = inform_L[361][1];				l_cell_reg[362] = inform_L[362][1];				l_cell_reg[363] = inform_L[363][1];				l_cell_reg[364] = inform_L[364][1];				l_cell_reg[365] = inform_L[365][1];				l_cell_reg[366] = inform_L[366][1];				l_cell_reg[367] = inform_L[367][1];				l_cell_reg[368] = inform_L[368][1];				l_cell_reg[369] = inform_L[369][1];				l_cell_reg[370] = inform_L[370][1];				l_cell_reg[371] = inform_L[371][1];				l_cell_reg[372] = inform_L[372][1];				l_cell_reg[373] = inform_L[373][1];				l_cell_reg[374] = inform_L[374][1];				l_cell_reg[375] = inform_L[375][1];				l_cell_reg[376] = inform_L[376][1];				l_cell_reg[377] = inform_L[377][1];				l_cell_reg[378] = inform_L[378][1];				l_cell_reg[379] = inform_L[379][1];				l_cell_reg[380] = inform_L[380][1];				l_cell_reg[381] = inform_L[381][1];				l_cell_reg[382] = inform_L[382][1];				l_cell_reg[383] = inform_L[383][1];				l_cell_reg[384] = inform_L[384][1];				l_cell_reg[385] = inform_L[385][1];				l_cell_reg[386] = inform_L[386][1];				l_cell_reg[387] = inform_L[387][1];				l_cell_reg[388] = inform_L[388][1];				l_cell_reg[389] = inform_L[389][1];				l_cell_reg[390] = inform_L[390][1];				l_cell_reg[391] = inform_L[391][1];				l_cell_reg[392] = inform_L[392][1];				l_cell_reg[393] = inform_L[393][1];				l_cell_reg[394] = inform_L[394][1];				l_cell_reg[395] = inform_L[395][1];				l_cell_reg[396] = inform_L[396][1];				l_cell_reg[397] = inform_L[397][1];				l_cell_reg[398] = inform_L[398][1];				l_cell_reg[399] = inform_L[399][1];				l_cell_reg[400] = inform_L[400][1];				l_cell_reg[401] = inform_L[401][1];				l_cell_reg[402] = inform_L[402][1];				l_cell_reg[403] = inform_L[403][1];				l_cell_reg[404] = inform_L[404][1];				l_cell_reg[405] = inform_L[405][1];				l_cell_reg[406] = inform_L[406][1];				l_cell_reg[407] = inform_L[407][1];				l_cell_reg[408] = inform_L[408][1];				l_cell_reg[409] = inform_L[409][1];				l_cell_reg[410] = inform_L[410][1];				l_cell_reg[411] = inform_L[411][1];				l_cell_reg[412] = inform_L[412][1];				l_cell_reg[413] = inform_L[413][1];				l_cell_reg[414] = inform_L[414][1];				l_cell_reg[415] = inform_L[415][1];				l_cell_reg[416] = inform_L[416][1];				l_cell_reg[417] = inform_L[417][1];				l_cell_reg[418] = inform_L[418][1];				l_cell_reg[419] = inform_L[419][1];				l_cell_reg[420] = inform_L[420][1];				l_cell_reg[421] = inform_L[421][1];				l_cell_reg[422] = inform_L[422][1];				l_cell_reg[423] = inform_L[423][1];				l_cell_reg[424] = inform_L[424][1];				l_cell_reg[425] = inform_L[425][1];				l_cell_reg[426] = inform_L[426][1];				l_cell_reg[427] = inform_L[427][1];				l_cell_reg[428] = inform_L[428][1];				l_cell_reg[429] = inform_L[429][1];				l_cell_reg[430] = inform_L[430][1];				l_cell_reg[431] = inform_L[431][1];				l_cell_reg[432] = inform_L[432][1];				l_cell_reg[433] = inform_L[433][1];				l_cell_reg[434] = inform_L[434][1];				l_cell_reg[435] = inform_L[435][1];				l_cell_reg[436] = inform_L[436][1];				l_cell_reg[437] = inform_L[437][1];				l_cell_reg[438] = inform_L[438][1];				l_cell_reg[439] = inform_L[439][1];				l_cell_reg[440] = inform_L[440][1];				l_cell_reg[441] = inform_L[441][1];				l_cell_reg[442] = inform_L[442][1];				l_cell_reg[443] = inform_L[443][1];				l_cell_reg[444] = inform_L[444][1];				l_cell_reg[445] = inform_L[445][1];				l_cell_reg[446] = inform_L[446][1];				l_cell_reg[447] = inform_L[447][1];				l_cell_reg[448] = inform_L[448][1];				l_cell_reg[449] = inform_L[449][1];				l_cell_reg[450] = inform_L[450][1];				l_cell_reg[451] = inform_L[451][1];				l_cell_reg[452] = inform_L[452][1];				l_cell_reg[453] = inform_L[453][1];				l_cell_reg[454] = inform_L[454][1];				l_cell_reg[455] = inform_L[455][1];				l_cell_reg[456] = inform_L[456][1];				l_cell_reg[457] = inform_L[457][1];				l_cell_reg[458] = inform_L[458][1];				l_cell_reg[459] = inform_L[459][1];				l_cell_reg[460] = inform_L[460][1];				l_cell_reg[461] = inform_L[461][1];				l_cell_reg[462] = inform_L[462][1];				l_cell_reg[463] = inform_L[463][1];				l_cell_reg[464] = inform_L[464][1];				l_cell_reg[465] = inform_L[465][1];				l_cell_reg[466] = inform_L[466][1];				l_cell_reg[467] = inform_L[467][1];				l_cell_reg[468] = inform_L[468][1];				l_cell_reg[469] = inform_L[469][1];				l_cell_reg[470] = inform_L[470][1];				l_cell_reg[471] = inform_L[471][1];				l_cell_reg[472] = inform_L[472][1];				l_cell_reg[473] = inform_L[473][1];				l_cell_reg[474] = inform_L[474][1];				l_cell_reg[475] = inform_L[475][1];				l_cell_reg[476] = inform_L[476][1];				l_cell_reg[477] = inform_L[477][1];				l_cell_reg[478] = inform_L[478][1];				l_cell_reg[479] = inform_L[479][1];				l_cell_reg[480] = inform_L[480][1];				l_cell_reg[481] = inform_L[481][1];				l_cell_reg[482] = inform_L[482][1];				l_cell_reg[483] = inform_L[483][1];				l_cell_reg[484] = inform_L[484][1];				l_cell_reg[485] = inform_L[485][1];				l_cell_reg[486] = inform_L[486][1];				l_cell_reg[487] = inform_L[487][1];				l_cell_reg[488] = inform_L[488][1];				l_cell_reg[489] = inform_L[489][1];				l_cell_reg[490] = inform_L[490][1];				l_cell_reg[491] = inform_L[491][1];				l_cell_reg[492] = inform_L[492][1];				l_cell_reg[493] = inform_L[493][1];				l_cell_reg[494] = inform_L[494][1];				l_cell_reg[495] = inform_L[495][1];				l_cell_reg[496] = inform_L[496][1];				l_cell_reg[497] = inform_L[497][1];				l_cell_reg[498] = inform_L[498][1];				l_cell_reg[499] = inform_L[499][1];				l_cell_reg[500] = inform_L[500][1];				l_cell_reg[501] = inform_L[501][1];				l_cell_reg[502] = inform_L[502][1];				l_cell_reg[503] = inform_L[503][1];				l_cell_reg[504] = inform_L[504][1];				l_cell_reg[505] = inform_L[505][1];				l_cell_reg[506] = inform_L[506][1];				l_cell_reg[507] = inform_L[507][1];				l_cell_reg[508] = inform_L[508][1];				l_cell_reg[509] = inform_L[509][1];				l_cell_reg[510] = inform_L[510][1];				l_cell_reg[511] = inform_L[511][1];				l_cell_reg[512] = inform_L[512][1];				l_cell_reg[513] = inform_L[513][1];				l_cell_reg[514] = inform_L[514][1];				l_cell_reg[515] = inform_L[515][1];				l_cell_reg[516] = inform_L[516][1];				l_cell_reg[517] = inform_L[517][1];				l_cell_reg[518] = inform_L[518][1];				l_cell_reg[519] = inform_L[519][1];				l_cell_reg[520] = inform_L[520][1];				l_cell_reg[521] = inform_L[521][1];				l_cell_reg[522] = inform_L[522][1];				l_cell_reg[523] = inform_L[523][1];				l_cell_reg[524] = inform_L[524][1];				l_cell_reg[525] = inform_L[525][1];				l_cell_reg[526] = inform_L[526][1];				l_cell_reg[527] = inform_L[527][1];				l_cell_reg[528] = inform_L[528][1];				l_cell_reg[529] = inform_L[529][1];				l_cell_reg[530] = inform_L[530][1];				l_cell_reg[531] = inform_L[531][1];				l_cell_reg[532] = inform_L[532][1];				l_cell_reg[533] = inform_L[533][1];				l_cell_reg[534] = inform_L[534][1];				l_cell_reg[535] = inform_L[535][1];				l_cell_reg[536] = inform_L[536][1];				l_cell_reg[537] = inform_L[537][1];				l_cell_reg[538] = inform_L[538][1];				l_cell_reg[539] = inform_L[539][1];				l_cell_reg[540] = inform_L[540][1];				l_cell_reg[541] = inform_L[541][1];				l_cell_reg[542] = inform_L[542][1];				l_cell_reg[543] = inform_L[543][1];				l_cell_reg[544] = inform_L[544][1];				l_cell_reg[545] = inform_L[545][1];				l_cell_reg[546] = inform_L[546][1];				l_cell_reg[547] = inform_L[547][1];				l_cell_reg[548] = inform_L[548][1];				l_cell_reg[549] = inform_L[549][1];				l_cell_reg[550] = inform_L[550][1];				l_cell_reg[551] = inform_L[551][1];				l_cell_reg[552] = inform_L[552][1];				l_cell_reg[553] = inform_L[553][1];				l_cell_reg[554] = inform_L[554][1];				l_cell_reg[555] = inform_L[555][1];				l_cell_reg[556] = inform_L[556][1];				l_cell_reg[557] = inform_L[557][1];				l_cell_reg[558] = inform_L[558][1];				l_cell_reg[559] = inform_L[559][1];				l_cell_reg[560] = inform_L[560][1];				l_cell_reg[561] = inform_L[561][1];				l_cell_reg[562] = inform_L[562][1];				l_cell_reg[563] = inform_L[563][1];				l_cell_reg[564] = inform_L[564][1];				l_cell_reg[565] = inform_L[565][1];				l_cell_reg[566] = inform_L[566][1];				l_cell_reg[567] = inform_L[567][1];				l_cell_reg[568] = inform_L[568][1];				l_cell_reg[569] = inform_L[569][1];				l_cell_reg[570] = inform_L[570][1];				l_cell_reg[571] = inform_L[571][1];				l_cell_reg[572] = inform_L[572][1];				l_cell_reg[573] = inform_L[573][1];				l_cell_reg[574] = inform_L[574][1];				l_cell_reg[575] = inform_L[575][1];				l_cell_reg[576] = inform_L[576][1];				l_cell_reg[577] = inform_L[577][1];				l_cell_reg[578] = inform_L[578][1];				l_cell_reg[579] = inform_L[579][1];				l_cell_reg[580] = inform_L[580][1];				l_cell_reg[581] = inform_L[581][1];				l_cell_reg[582] = inform_L[582][1];				l_cell_reg[583] = inform_L[583][1];				l_cell_reg[584] = inform_L[584][1];				l_cell_reg[585] = inform_L[585][1];				l_cell_reg[586] = inform_L[586][1];				l_cell_reg[587] = inform_L[587][1];				l_cell_reg[588] = inform_L[588][1];				l_cell_reg[589] = inform_L[589][1];				l_cell_reg[590] = inform_L[590][1];				l_cell_reg[591] = inform_L[591][1];				l_cell_reg[592] = inform_L[592][1];				l_cell_reg[593] = inform_L[593][1];				l_cell_reg[594] = inform_L[594][1];				l_cell_reg[595] = inform_L[595][1];				l_cell_reg[596] = inform_L[596][1];				l_cell_reg[597] = inform_L[597][1];				l_cell_reg[598] = inform_L[598][1];				l_cell_reg[599] = inform_L[599][1];				l_cell_reg[600] = inform_L[600][1];				l_cell_reg[601] = inform_L[601][1];				l_cell_reg[602] = inform_L[602][1];				l_cell_reg[603] = inform_L[603][1];				l_cell_reg[604] = inform_L[604][1];				l_cell_reg[605] = inform_L[605][1];				l_cell_reg[606] = inform_L[606][1];				l_cell_reg[607] = inform_L[607][1];				l_cell_reg[608] = inform_L[608][1];				l_cell_reg[609] = inform_L[609][1];				l_cell_reg[610] = inform_L[610][1];				l_cell_reg[611] = inform_L[611][1];				l_cell_reg[612] = inform_L[612][1];				l_cell_reg[613] = inform_L[613][1];				l_cell_reg[614] = inform_L[614][1];				l_cell_reg[615] = inform_L[615][1];				l_cell_reg[616] = inform_L[616][1];				l_cell_reg[617] = inform_L[617][1];				l_cell_reg[618] = inform_L[618][1];				l_cell_reg[619] = inform_L[619][1];				l_cell_reg[620] = inform_L[620][1];				l_cell_reg[621] = inform_L[621][1];				l_cell_reg[622] = inform_L[622][1];				l_cell_reg[623] = inform_L[623][1];				l_cell_reg[624] = inform_L[624][1];				l_cell_reg[625] = inform_L[625][1];				l_cell_reg[626] = inform_L[626][1];				l_cell_reg[627] = inform_L[627][1];				l_cell_reg[628] = inform_L[628][1];				l_cell_reg[629] = inform_L[629][1];				l_cell_reg[630] = inform_L[630][1];				l_cell_reg[631] = inform_L[631][1];				l_cell_reg[632] = inform_L[632][1];				l_cell_reg[633] = inform_L[633][1];				l_cell_reg[634] = inform_L[634][1];				l_cell_reg[635] = inform_L[635][1];				l_cell_reg[636] = inform_L[636][1];				l_cell_reg[637] = inform_L[637][1];				l_cell_reg[638] = inform_L[638][1];				l_cell_reg[639] = inform_L[639][1];				l_cell_reg[640] = inform_L[640][1];				l_cell_reg[641] = inform_L[641][1];				l_cell_reg[642] = inform_L[642][1];				l_cell_reg[643] = inform_L[643][1];				l_cell_reg[644] = inform_L[644][1];				l_cell_reg[645] = inform_L[645][1];				l_cell_reg[646] = inform_L[646][1];				l_cell_reg[647] = inform_L[647][1];				l_cell_reg[648] = inform_L[648][1];				l_cell_reg[649] = inform_L[649][1];				l_cell_reg[650] = inform_L[650][1];				l_cell_reg[651] = inform_L[651][1];				l_cell_reg[652] = inform_L[652][1];				l_cell_reg[653] = inform_L[653][1];				l_cell_reg[654] = inform_L[654][1];				l_cell_reg[655] = inform_L[655][1];				l_cell_reg[656] = inform_L[656][1];				l_cell_reg[657] = inform_L[657][1];				l_cell_reg[658] = inform_L[658][1];				l_cell_reg[659] = inform_L[659][1];				l_cell_reg[660] = inform_L[660][1];				l_cell_reg[661] = inform_L[661][1];				l_cell_reg[662] = inform_L[662][1];				l_cell_reg[663] = inform_L[663][1];				l_cell_reg[664] = inform_L[664][1];				l_cell_reg[665] = inform_L[665][1];				l_cell_reg[666] = inform_L[666][1];				l_cell_reg[667] = inform_L[667][1];				l_cell_reg[668] = inform_L[668][1];				l_cell_reg[669] = inform_L[669][1];				l_cell_reg[670] = inform_L[670][1];				l_cell_reg[671] = inform_L[671][1];				l_cell_reg[672] = inform_L[672][1];				l_cell_reg[673] = inform_L[673][1];				l_cell_reg[674] = inform_L[674][1];				l_cell_reg[675] = inform_L[675][1];				l_cell_reg[676] = inform_L[676][1];				l_cell_reg[677] = inform_L[677][1];				l_cell_reg[678] = inform_L[678][1];				l_cell_reg[679] = inform_L[679][1];				l_cell_reg[680] = inform_L[680][1];				l_cell_reg[681] = inform_L[681][1];				l_cell_reg[682] = inform_L[682][1];				l_cell_reg[683] = inform_L[683][1];				l_cell_reg[684] = inform_L[684][1];				l_cell_reg[685] = inform_L[685][1];				l_cell_reg[686] = inform_L[686][1];				l_cell_reg[687] = inform_L[687][1];				l_cell_reg[688] = inform_L[688][1];				l_cell_reg[689] = inform_L[689][1];				l_cell_reg[690] = inform_L[690][1];				l_cell_reg[691] = inform_L[691][1];				l_cell_reg[692] = inform_L[692][1];				l_cell_reg[693] = inform_L[693][1];				l_cell_reg[694] = inform_L[694][1];				l_cell_reg[695] = inform_L[695][1];				l_cell_reg[696] = inform_L[696][1];				l_cell_reg[697] = inform_L[697][1];				l_cell_reg[698] = inform_L[698][1];				l_cell_reg[699] = inform_L[699][1];				l_cell_reg[700] = inform_L[700][1];				l_cell_reg[701] = inform_L[701][1];				l_cell_reg[702] = inform_L[702][1];				l_cell_reg[703] = inform_L[703][1];				l_cell_reg[704] = inform_L[704][1];				l_cell_reg[705] = inform_L[705][1];				l_cell_reg[706] = inform_L[706][1];				l_cell_reg[707] = inform_L[707][1];				l_cell_reg[708] = inform_L[708][1];				l_cell_reg[709] = inform_L[709][1];				l_cell_reg[710] = inform_L[710][1];				l_cell_reg[711] = inform_L[711][1];				l_cell_reg[712] = inform_L[712][1];				l_cell_reg[713] = inform_L[713][1];				l_cell_reg[714] = inform_L[714][1];				l_cell_reg[715] = inform_L[715][1];				l_cell_reg[716] = inform_L[716][1];				l_cell_reg[717] = inform_L[717][1];				l_cell_reg[718] = inform_L[718][1];				l_cell_reg[719] = inform_L[719][1];				l_cell_reg[720] = inform_L[720][1];				l_cell_reg[721] = inform_L[721][1];				l_cell_reg[722] = inform_L[722][1];				l_cell_reg[723] = inform_L[723][1];				l_cell_reg[724] = inform_L[724][1];				l_cell_reg[725] = inform_L[725][1];				l_cell_reg[726] = inform_L[726][1];				l_cell_reg[727] = inform_L[727][1];				l_cell_reg[728] = inform_L[728][1];				l_cell_reg[729] = inform_L[729][1];				l_cell_reg[730] = inform_L[730][1];				l_cell_reg[731] = inform_L[731][1];				l_cell_reg[732] = inform_L[732][1];				l_cell_reg[733] = inform_L[733][1];				l_cell_reg[734] = inform_L[734][1];				l_cell_reg[735] = inform_L[735][1];				l_cell_reg[736] = inform_L[736][1];				l_cell_reg[737] = inform_L[737][1];				l_cell_reg[738] = inform_L[738][1];				l_cell_reg[739] = inform_L[739][1];				l_cell_reg[740] = inform_L[740][1];				l_cell_reg[741] = inform_L[741][1];				l_cell_reg[742] = inform_L[742][1];				l_cell_reg[743] = inform_L[743][1];				l_cell_reg[744] = inform_L[744][1];				l_cell_reg[745] = inform_L[745][1];				l_cell_reg[746] = inform_L[746][1];				l_cell_reg[747] = inform_L[747][1];				l_cell_reg[748] = inform_L[748][1];				l_cell_reg[749] = inform_L[749][1];				l_cell_reg[750] = inform_L[750][1];				l_cell_reg[751] = inform_L[751][1];				l_cell_reg[752] = inform_L[752][1];				l_cell_reg[753] = inform_L[753][1];				l_cell_reg[754] = inform_L[754][1];				l_cell_reg[755] = inform_L[755][1];				l_cell_reg[756] = inform_L[756][1];				l_cell_reg[757] = inform_L[757][1];				l_cell_reg[758] = inform_L[758][1];				l_cell_reg[759] = inform_L[759][1];				l_cell_reg[760] = inform_L[760][1];				l_cell_reg[761] = inform_L[761][1];				l_cell_reg[762] = inform_L[762][1];				l_cell_reg[763] = inform_L[763][1];				l_cell_reg[764] = inform_L[764][1];				l_cell_reg[765] = inform_L[765][1];				l_cell_reg[766] = inform_L[766][1];				l_cell_reg[767] = inform_L[767][1];				l_cell_reg[768] = inform_L[768][1];				l_cell_reg[769] = inform_L[769][1];				l_cell_reg[770] = inform_L[770][1];				l_cell_reg[771] = inform_L[771][1];				l_cell_reg[772] = inform_L[772][1];				l_cell_reg[773] = inform_L[773][1];				l_cell_reg[774] = inform_L[774][1];				l_cell_reg[775] = inform_L[775][1];				l_cell_reg[776] = inform_L[776][1];				l_cell_reg[777] = inform_L[777][1];				l_cell_reg[778] = inform_L[778][1];				l_cell_reg[779] = inform_L[779][1];				l_cell_reg[780] = inform_L[780][1];				l_cell_reg[781] = inform_L[781][1];				l_cell_reg[782] = inform_L[782][1];				l_cell_reg[783] = inform_L[783][1];				l_cell_reg[784] = inform_L[784][1];				l_cell_reg[785] = inform_L[785][1];				l_cell_reg[786] = inform_L[786][1];				l_cell_reg[787] = inform_L[787][1];				l_cell_reg[788] = inform_L[788][1];				l_cell_reg[789] = inform_L[789][1];				l_cell_reg[790] = inform_L[790][1];				l_cell_reg[791] = inform_L[791][1];				l_cell_reg[792] = inform_L[792][1];				l_cell_reg[793] = inform_L[793][1];				l_cell_reg[794] = inform_L[794][1];				l_cell_reg[795] = inform_L[795][1];				l_cell_reg[796] = inform_L[796][1];				l_cell_reg[797] = inform_L[797][1];				l_cell_reg[798] = inform_L[798][1];				l_cell_reg[799] = inform_L[799][1];				l_cell_reg[800] = inform_L[800][1];				l_cell_reg[801] = inform_L[801][1];				l_cell_reg[802] = inform_L[802][1];				l_cell_reg[803] = inform_L[803][1];				l_cell_reg[804] = inform_L[804][1];				l_cell_reg[805] = inform_L[805][1];				l_cell_reg[806] = inform_L[806][1];				l_cell_reg[807] = inform_L[807][1];				l_cell_reg[808] = inform_L[808][1];				l_cell_reg[809] = inform_L[809][1];				l_cell_reg[810] = inform_L[810][1];				l_cell_reg[811] = inform_L[811][1];				l_cell_reg[812] = inform_L[812][1];				l_cell_reg[813] = inform_L[813][1];				l_cell_reg[814] = inform_L[814][1];				l_cell_reg[815] = inform_L[815][1];				l_cell_reg[816] = inform_L[816][1];				l_cell_reg[817] = inform_L[817][1];				l_cell_reg[818] = inform_L[818][1];				l_cell_reg[819] = inform_L[819][1];				l_cell_reg[820] = inform_L[820][1];				l_cell_reg[821] = inform_L[821][1];				l_cell_reg[822] = inform_L[822][1];				l_cell_reg[823] = inform_L[823][1];				l_cell_reg[824] = inform_L[824][1];				l_cell_reg[825] = inform_L[825][1];				l_cell_reg[826] = inform_L[826][1];				l_cell_reg[827] = inform_L[827][1];				l_cell_reg[828] = inform_L[828][1];				l_cell_reg[829] = inform_L[829][1];				l_cell_reg[830] = inform_L[830][1];				l_cell_reg[831] = inform_L[831][1];				l_cell_reg[832] = inform_L[832][1];				l_cell_reg[833] = inform_L[833][1];				l_cell_reg[834] = inform_L[834][1];				l_cell_reg[835] = inform_L[835][1];				l_cell_reg[836] = inform_L[836][1];				l_cell_reg[837] = inform_L[837][1];				l_cell_reg[838] = inform_L[838][1];				l_cell_reg[839] = inform_L[839][1];				l_cell_reg[840] = inform_L[840][1];				l_cell_reg[841] = inform_L[841][1];				l_cell_reg[842] = inform_L[842][1];				l_cell_reg[843] = inform_L[843][1];				l_cell_reg[844] = inform_L[844][1];				l_cell_reg[845] = inform_L[845][1];				l_cell_reg[846] = inform_L[846][1];				l_cell_reg[847] = inform_L[847][1];				l_cell_reg[848] = inform_L[848][1];				l_cell_reg[849] = inform_L[849][1];				l_cell_reg[850] = inform_L[850][1];				l_cell_reg[851] = inform_L[851][1];				l_cell_reg[852] = inform_L[852][1];				l_cell_reg[853] = inform_L[853][1];				l_cell_reg[854] = inform_L[854][1];				l_cell_reg[855] = inform_L[855][1];				l_cell_reg[856] = inform_L[856][1];				l_cell_reg[857] = inform_L[857][1];				l_cell_reg[858] = inform_L[858][1];				l_cell_reg[859] = inform_L[859][1];				l_cell_reg[860] = inform_L[860][1];				l_cell_reg[861] = inform_L[861][1];				l_cell_reg[862] = inform_L[862][1];				l_cell_reg[863] = inform_L[863][1];				l_cell_reg[864] = inform_L[864][1];				l_cell_reg[865] = inform_L[865][1];				l_cell_reg[866] = inform_L[866][1];				l_cell_reg[867] = inform_L[867][1];				l_cell_reg[868] = inform_L[868][1];				l_cell_reg[869] = inform_L[869][1];				l_cell_reg[870] = inform_L[870][1];				l_cell_reg[871] = inform_L[871][1];				l_cell_reg[872] = inform_L[872][1];				l_cell_reg[873] = inform_L[873][1];				l_cell_reg[874] = inform_L[874][1];				l_cell_reg[875] = inform_L[875][1];				l_cell_reg[876] = inform_L[876][1];				l_cell_reg[877] = inform_L[877][1];				l_cell_reg[878] = inform_L[878][1];				l_cell_reg[879] = inform_L[879][1];				l_cell_reg[880] = inform_L[880][1];				l_cell_reg[881] = inform_L[881][1];				l_cell_reg[882] = inform_L[882][1];				l_cell_reg[883] = inform_L[883][1];				l_cell_reg[884] = inform_L[884][1];				l_cell_reg[885] = inform_L[885][1];				l_cell_reg[886] = inform_L[886][1];				l_cell_reg[887] = inform_L[887][1];				l_cell_reg[888] = inform_L[888][1];				l_cell_reg[889] = inform_L[889][1];				l_cell_reg[890] = inform_L[890][1];				l_cell_reg[891] = inform_L[891][1];				l_cell_reg[892] = inform_L[892][1];				l_cell_reg[893] = inform_L[893][1];				l_cell_reg[894] = inform_L[894][1];				l_cell_reg[895] = inform_L[895][1];				l_cell_reg[896] = inform_L[896][1];				l_cell_reg[897] = inform_L[897][1];				l_cell_reg[898] = inform_L[898][1];				l_cell_reg[899] = inform_L[899][1];				l_cell_reg[900] = inform_L[900][1];				l_cell_reg[901] = inform_L[901][1];				l_cell_reg[902] = inform_L[902][1];				l_cell_reg[903] = inform_L[903][1];				l_cell_reg[904] = inform_L[904][1];				l_cell_reg[905] = inform_L[905][1];				l_cell_reg[906] = inform_L[906][1];				l_cell_reg[907] = inform_L[907][1];				l_cell_reg[908] = inform_L[908][1];				l_cell_reg[909] = inform_L[909][1];				l_cell_reg[910] = inform_L[910][1];				l_cell_reg[911] = inform_L[911][1];				l_cell_reg[912] = inform_L[912][1];				l_cell_reg[913] = inform_L[913][1];				l_cell_reg[914] = inform_L[914][1];				l_cell_reg[915] = inform_L[915][1];				l_cell_reg[916] = inform_L[916][1];				l_cell_reg[917] = inform_L[917][1];				l_cell_reg[918] = inform_L[918][1];				l_cell_reg[919] = inform_L[919][1];				l_cell_reg[920] = inform_L[920][1];				l_cell_reg[921] = inform_L[921][1];				l_cell_reg[922] = inform_L[922][1];				l_cell_reg[923] = inform_L[923][1];				l_cell_reg[924] = inform_L[924][1];				l_cell_reg[925] = inform_L[925][1];				l_cell_reg[926] = inform_L[926][1];				l_cell_reg[927] = inform_L[927][1];				l_cell_reg[928] = inform_L[928][1];				l_cell_reg[929] = inform_L[929][1];				l_cell_reg[930] = inform_L[930][1];				l_cell_reg[931] = inform_L[931][1];				l_cell_reg[932] = inform_L[932][1];				l_cell_reg[933] = inform_L[933][1];				l_cell_reg[934] = inform_L[934][1];				l_cell_reg[935] = inform_L[935][1];				l_cell_reg[936] = inform_L[936][1];				l_cell_reg[937] = inform_L[937][1];				l_cell_reg[938] = inform_L[938][1];				l_cell_reg[939] = inform_L[939][1];				l_cell_reg[940] = inform_L[940][1];				l_cell_reg[941] = inform_L[941][1];				l_cell_reg[942] = inform_L[942][1];				l_cell_reg[943] = inform_L[943][1];				l_cell_reg[944] = inform_L[944][1];				l_cell_reg[945] = inform_L[945][1];				l_cell_reg[946] = inform_L[946][1];				l_cell_reg[947] = inform_L[947][1];				l_cell_reg[948] = inform_L[948][1];				l_cell_reg[949] = inform_L[949][1];				l_cell_reg[950] = inform_L[950][1];				l_cell_reg[951] = inform_L[951][1];				l_cell_reg[952] = inform_L[952][1];				l_cell_reg[953] = inform_L[953][1];				l_cell_reg[954] = inform_L[954][1];				l_cell_reg[955] = inform_L[955][1];				l_cell_reg[956] = inform_L[956][1];				l_cell_reg[957] = inform_L[957][1];				l_cell_reg[958] = inform_L[958][1];				l_cell_reg[959] = inform_L[959][1];				l_cell_reg[960] = inform_L[960][1];				l_cell_reg[961] = inform_L[961][1];				l_cell_reg[962] = inform_L[962][1];				l_cell_reg[963] = inform_L[963][1];				l_cell_reg[964] = inform_L[964][1];				l_cell_reg[965] = inform_L[965][1];				l_cell_reg[966] = inform_L[966][1];				l_cell_reg[967] = inform_L[967][1];				l_cell_reg[968] = inform_L[968][1];				l_cell_reg[969] = inform_L[969][1];				l_cell_reg[970] = inform_L[970][1];				l_cell_reg[971] = inform_L[971][1];				l_cell_reg[972] = inform_L[972][1];				l_cell_reg[973] = inform_L[973][1];				l_cell_reg[974] = inform_L[974][1];				l_cell_reg[975] = inform_L[975][1];				l_cell_reg[976] = inform_L[976][1];				l_cell_reg[977] = inform_L[977][1];				l_cell_reg[978] = inform_L[978][1];				l_cell_reg[979] = inform_L[979][1];				l_cell_reg[980] = inform_L[980][1];				l_cell_reg[981] = inform_L[981][1];				l_cell_reg[982] = inform_L[982][1];				l_cell_reg[983] = inform_L[983][1];				l_cell_reg[984] = inform_L[984][1];				l_cell_reg[985] = inform_L[985][1];				l_cell_reg[986] = inform_L[986][1];				l_cell_reg[987] = inform_L[987][1];				l_cell_reg[988] = inform_L[988][1];				l_cell_reg[989] = inform_L[989][1];				l_cell_reg[990] = inform_L[990][1];				l_cell_reg[991] = inform_L[991][1];				l_cell_reg[992] = inform_L[992][1];				l_cell_reg[993] = inform_L[993][1];				l_cell_reg[994] = inform_L[994][1];				l_cell_reg[995] = inform_L[995][1];				l_cell_reg[996] = inform_L[996][1];				l_cell_reg[997] = inform_L[997][1];				l_cell_reg[998] = inform_L[998][1];				l_cell_reg[999] = inform_L[999][1];				l_cell_reg[1000] = inform_L[1000][1];				l_cell_reg[1001] = inform_L[1001][1];				l_cell_reg[1002] = inform_L[1002][1];				l_cell_reg[1003] = inform_L[1003][1];				l_cell_reg[1004] = inform_L[1004][1];				l_cell_reg[1005] = inform_L[1005][1];				l_cell_reg[1006] = inform_L[1006][1];				l_cell_reg[1007] = inform_L[1007][1];				l_cell_reg[1008] = inform_L[1008][1];				l_cell_reg[1009] = inform_L[1009][1];				l_cell_reg[1010] = inform_L[1010][1];				l_cell_reg[1011] = inform_L[1011][1];				l_cell_reg[1012] = inform_L[1012][1];				l_cell_reg[1013] = inform_L[1013][1];				l_cell_reg[1014] = inform_L[1014][1];				l_cell_reg[1015] = inform_L[1015][1];				l_cell_reg[1016] = inform_L[1016][1];				l_cell_reg[1017] = inform_L[1017][1];				l_cell_reg[1018] = inform_L[1018][1];				l_cell_reg[1019] = inform_L[1019][1];				l_cell_reg[1020] = inform_L[1020][1];				l_cell_reg[1021] = inform_L[1021][1];				l_cell_reg[1022] = inform_L[1022][1];				l_cell_reg[1023] = inform_L[1023][1];			end
			2:			begin				r_cell_reg[0] = inform_R[0][1];				r_cell_reg[1] = inform_R[2][1];				r_cell_reg[2] = inform_R[1][1];				r_cell_reg[3] = inform_R[3][1];				r_cell_reg[4] = inform_R[4][1];				r_cell_reg[5] = inform_R[6][1];				r_cell_reg[6] = inform_R[5][1];				r_cell_reg[7] = inform_R[7][1];				r_cell_reg[8] = inform_R[8][1];				r_cell_reg[9] = inform_R[10][1];				r_cell_reg[10] = inform_R[9][1];				r_cell_reg[11] = inform_R[11][1];				r_cell_reg[12] = inform_R[12][1];				r_cell_reg[13] = inform_R[14][1];				r_cell_reg[14] = inform_R[13][1];				r_cell_reg[15] = inform_R[15][1];				r_cell_reg[16] = inform_R[16][1];				r_cell_reg[17] = inform_R[18][1];				r_cell_reg[18] = inform_R[17][1];				r_cell_reg[19] = inform_R[19][1];				r_cell_reg[20] = inform_R[20][1];				r_cell_reg[21] = inform_R[22][1];				r_cell_reg[22] = inform_R[21][1];				r_cell_reg[23] = inform_R[23][1];				r_cell_reg[24] = inform_R[24][1];				r_cell_reg[25] = inform_R[26][1];				r_cell_reg[26] = inform_R[25][1];				r_cell_reg[27] = inform_R[27][1];				r_cell_reg[28] = inform_R[28][1];				r_cell_reg[29] = inform_R[30][1];				r_cell_reg[30] = inform_R[29][1];				r_cell_reg[31] = inform_R[31][1];				r_cell_reg[32] = inform_R[32][1];				r_cell_reg[33] = inform_R[34][1];				r_cell_reg[34] = inform_R[33][1];				r_cell_reg[35] = inform_R[35][1];				r_cell_reg[36] = inform_R[36][1];				r_cell_reg[37] = inform_R[38][1];				r_cell_reg[38] = inform_R[37][1];				r_cell_reg[39] = inform_R[39][1];				r_cell_reg[40] = inform_R[40][1];				r_cell_reg[41] = inform_R[42][1];				r_cell_reg[42] = inform_R[41][1];				r_cell_reg[43] = inform_R[43][1];				r_cell_reg[44] = inform_R[44][1];				r_cell_reg[45] = inform_R[46][1];				r_cell_reg[46] = inform_R[45][1];				r_cell_reg[47] = inform_R[47][1];				r_cell_reg[48] = inform_R[48][1];				r_cell_reg[49] = inform_R[50][1];				r_cell_reg[50] = inform_R[49][1];				r_cell_reg[51] = inform_R[51][1];				r_cell_reg[52] = inform_R[52][1];				r_cell_reg[53] = inform_R[54][1];				r_cell_reg[54] = inform_R[53][1];				r_cell_reg[55] = inform_R[55][1];				r_cell_reg[56] = inform_R[56][1];				r_cell_reg[57] = inform_R[58][1];				r_cell_reg[58] = inform_R[57][1];				r_cell_reg[59] = inform_R[59][1];				r_cell_reg[60] = inform_R[60][1];				r_cell_reg[61] = inform_R[62][1];				r_cell_reg[62] = inform_R[61][1];				r_cell_reg[63] = inform_R[63][1];				r_cell_reg[64] = inform_R[64][1];				r_cell_reg[65] = inform_R[66][1];				r_cell_reg[66] = inform_R[65][1];				r_cell_reg[67] = inform_R[67][1];				r_cell_reg[68] = inform_R[68][1];				r_cell_reg[69] = inform_R[70][1];				r_cell_reg[70] = inform_R[69][1];				r_cell_reg[71] = inform_R[71][1];				r_cell_reg[72] = inform_R[72][1];				r_cell_reg[73] = inform_R[74][1];				r_cell_reg[74] = inform_R[73][1];				r_cell_reg[75] = inform_R[75][1];				r_cell_reg[76] = inform_R[76][1];				r_cell_reg[77] = inform_R[78][1];				r_cell_reg[78] = inform_R[77][1];				r_cell_reg[79] = inform_R[79][1];				r_cell_reg[80] = inform_R[80][1];				r_cell_reg[81] = inform_R[82][1];				r_cell_reg[82] = inform_R[81][1];				r_cell_reg[83] = inform_R[83][1];				r_cell_reg[84] = inform_R[84][1];				r_cell_reg[85] = inform_R[86][1];				r_cell_reg[86] = inform_R[85][1];				r_cell_reg[87] = inform_R[87][1];				r_cell_reg[88] = inform_R[88][1];				r_cell_reg[89] = inform_R[90][1];				r_cell_reg[90] = inform_R[89][1];				r_cell_reg[91] = inform_R[91][1];				r_cell_reg[92] = inform_R[92][1];				r_cell_reg[93] = inform_R[94][1];				r_cell_reg[94] = inform_R[93][1];				r_cell_reg[95] = inform_R[95][1];				r_cell_reg[96] = inform_R[96][1];				r_cell_reg[97] = inform_R[98][1];				r_cell_reg[98] = inform_R[97][1];				r_cell_reg[99] = inform_R[99][1];				r_cell_reg[100] = inform_R[100][1];				r_cell_reg[101] = inform_R[102][1];				r_cell_reg[102] = inform_R[101][1];				r_cell_reg[103] = inform_R[103][1];				r_cell_reg[104] = inform_R[104][1];				r_cell_reg[105] = inform_R[106][1];				r_cell_reg[106] = inform_R[105][1];				r_cell_reg[107] = inform_R[107][1];				r_cell_reg[108] = inform_R[108][1];				r_cell_reg[109] = inform_R[110][1];				r_cell_reg[110] = inform_R[109][1];				r_cell_reg[111] = inform_R[111][1];				r_cell_reg[112] = inform_R[112][1];				r_cell_reg[113] = inform_R[114][1];				r_cell_reg[114] = inform_R[113][1];				r_cell_reg[115] = inform_R[115][1];				r_cell_reg[116] = inform_R[116][1];				r_cell_reg[117] = inform_R[118][1];				r_cell_reg[118] = inform_R[117][1];				r_cell_reg[119] = inform_R[119][1];				r_cell_reg[120] = inform_R[120][1];				r_cell_reg[121] = inform_R[122][1];				r_cell_reg[122] = inform_R[121][1];				r_cell_reg[123] = inform_R[123][1];				r_cell_reg[124] = inform_R[124][1];				r_cell_reg[125] = inform_R[126][1];				r_cell_reg[126] = inform_R[125][1];				r_cell_reg[127] = inform_R[127][1];				r_cell_reg[128] = inform_R[128][1];				r_cell_reg[129] = inform_R[130][1];				r_cell_reg[130] = inform_R[129][1];				r_cell_reg[131] = inform_R[131][1];				r_cell_reg[132] = inform_R[132][1];				r_cell_reg[133] = inform_R[134][1];				r_cell_reg[134] = inform_R[133][1];				r_cell_reg[135] = inform_R[135][1];				r_cell_reg[136] = inform_R[136][1];				r_cell_reg[137] = inform_R[138][1];				r_cell_reg[138] = inform_R[137][1];				r_cell_reg[139] = inform_R[139][1];				r_cell_reg[140] = inform_R[140][1];				r_cell_reg[141] = inform_R[142][1];				r_cell_reg[142] = inform_R[141][1];				r_cell_reg[143] = inform_R[143][1];				r_cell_reg[144] = inform_R[144][1];				r_cell_reg[145] = inform_R[146][1];				r_cell_reg[146] = inform_R[145][1];				r_cell_reg[147] = inform_R[147][1];				r_cell_reg[148] = inform_R[148][1];				r_cell_reg[149] = inform_R[150][1];				r_cell_reg[150] = inform_R[149][1];				r_cell_reg[151] = inform_R[151][1];				r_cell_reg[152] = inform_R[152][1];				r_cell_reg[153] = inform_R[154][1];				r_cell_reg[154] = inform_R[153][1];				r_cell_reg[155] = inform_R[155][1];				r_cell_reg[156] = inform_R[156][1];				r_cell_reg[157] = inform_R[158][1];				r_cell_reg[158] = inform_R[157][1];				r_cell_reg[159] = inform_R[159][1];				r_cell_reg[160] = inform_R[160][1];				r_cell_reg[161] = inform_R[162][1];				r_cell_reg[162] = inform_R[161][1];				r_cell_reg[163] = inform_R[163][1];				r_cell_reg[164] = inform_R[164][1];				r_cell_reg[165] = inform_R[166][1];				r_cell_reg[166] = inform_R[165][1];				r_cell_reg[167] = inform_R[167][1];				r_cell_reg[168] = inform_R[168][1];				r_cell_reg[169] = inform_R[170][1];				r_cell_reg[170] = inform_R[169][1];				r_cell_reg[171] = inform_R[171][1];				r_cell_reg[172] = inform_R[172][1];				r_cell_reg[173] = inform_R[174][1];				r_cell_reg[174] = inform_R[173][1];				r_cell_reg[175] = inform_R[175][1];				r_cell_reg[176] = inform_R[176][1];				r_cell_reg[177] = inform_R[178][1];				r_cell_reg[178] = inform_R[177][1];				r_cell_reg[179] = inform_R[179][1];				r_cell_reg[180] = inform_R[180][1];				r_cell_reg[181] = inform_R[182][1];				r_cell_reg[182] = inform_R[181][1];				r_cell_reg[183] = inform_R[183][1];				r_cell_reg[184] = inform_R[184][1];				r_cell_reg[185] = inform_R[186][1];				r_cell_reg[186] = inform_R[185][1];				r_cell_reg[187] = inform_R[187][1];				r_cell_reg[188] = inform_R[188][1];				r_cell_reg[189] = inform_R[190][1];				r_cell_reg[190] = inform_R[189][1];				r_cell_reg[191] = inform_R[191][1];				r_cell_reg[192] = inform_R[192][1];				r_cell_reg[193] = inform_R[194][1];				r_cell_reg[194] = inform_R[193][1];				r_cell_reg[195] = inform_R[195][1];				r_cell_reg[196] = inform_R[196][1];				r_cell_reg[197] = inform_R[198][1];				r_cell_reg[198] = inform_R[197][1];				r_cell_reg[199] = inform_R[199][1];				r_cell_reg[200] = inform_R[200][1];				r_cell_reg[201] = inform_R[202][1];				r_cell_reg[202] = inform_R[201][1];				r_cell_reg[203] = inform_R[203][1];				r_cell_reg[204] = inform_R[204][1];				r_cell_reg[205] = inform_R[206][1];				r_cell_reg[206] = inform_R[205][1];				r_cell_reg[207] = inform_R[207][1];				r_cell_reg[208] = inform_R[208][1];				r_cell_reg[209] = inform_R[210][1];				r_cell_reg[210] = inform_R[209][1];				r_cell_reg[211] = inform_R[211][1];				r_cell_reg[212] = inform_R[212][1];				r_cell_reg[213] = inform_R[214][1];				r_cell_reg[214] = inform_R[213][1];				r_cell_reg[215] = inform_R[215][1];				r_cell_reg[216] = inform_R[216][1];				r_cell_reg[217] = inform_R[218][1];				r_cell_reg[218] = inform_R[217][1];				r_cell_reg[219] = inform_R[219][1];				r_cell_reg[220] = inform_R[220][1];				r_cell_reg[221] = inform_R[222][1];				r_cell_reg[222] = inform_R[221][1];				r_cell_reg[223] = inform_R[223][1];				r_cell_reg[224] = inform_R[224][1];				r_cell_reg[225] = inform_R[226][1];				r_cell_reg[226] = inform_R[225][1];				r_cell_reg[227] = inform_R[227][1];				r_cell_reg[228] = inform_R[228][1];				r_cell_reg[229] = inform_R[230][1];				r_cell_reg[230] = inform_R[229][1];				r_cell_reg[231] = inform_R[231][1];				r_cell_reg[232] = inform_R[232][1];				r_cell_reg[233] = inform_R[234][1];				r_cell_reg[234] = inform_R[233][1];				r_cell_reg[235] = inform_R[235][1];				r_cell_reg[236] = inform_R[236][1];				r_cell_reg[237] = inform_R[238][1];				r_cell_reg[238] = inform_R[237][1];				r_cell_reg[239] = inform_R[239][1];				r_cell_reg[240] = inform_R[240][1];				r_cell_reg[241] = inform_R[242][1];				r_cell_reg[242] = inform_R[241][1];				r_cell_reg[243] = inform_R[243][1];				r_cell_reg[244] = inform_R[244][1];				r_cell_reg[245] = inform_R[246][1];				r_cell_reg[246] = inform_R[245][1];				r_cell_reg[247] = inform_R[247][1];				r_cell_reg[248] = inform_R[248][1];				r_cell_reg[249] = inform_R[250][1];				r_cell_reg[250] = inform_R[249][1];				r_cell_reg[251] = inform_R[251][1];				r_cell_reg[252] = inform_R[252][1];				r_cell_reg[253] = inform_R[254][1];				r_cell_reg[254] = inform_R[253][1];				r_cell_reg[255] = inform_R[255][1];				r_cell_reg[256] = inform_R[256][1];				r_cell_reg[257] = inform_R[258][1];				r_cell_reg[258] = inform_R[257][1];				r_cell_reg[259] = inform_R[259][1];				r_cell_reg[260] = inform_R[260][1];				r_cell_reg[261] = inform_R[262][1];				r_cell_reg[262] = inform_R[261][1];				r_cell_reg[263] = inform_R[263][1];				r_cell_reg[264] = inform_R[264][1];				r_cell_reg[265] = inform_R[266][1];				r_cell_reg[266] = inform_R[265][1];				r_cell_reg[267] = inform_R[267][1];				r_cell_reg[268] = inform_R[268][1];				r_cell_reg[269] = inform_R[270][1];				r_cell_reg[270] = inform_R[269][1];				r_cell_reg[271] = inform_R[271][1];				r_cell_reg[272] = inform_R[272][1];				r_cell_reg[273] = inform_R[274][1];				r_cell_reg[274] = inform_R[273][1];				r_cell_reg[275] = inform_R[275][1];				r_cell_reg[276] = inform_R[276][1];				r_cell_reg[277] = inform_R[278][1];				r_cell_reg[278] = inform_R[277][1];				r_cell_reg[279] = inform_R[279][1];				r_cell_reg[280] = inform_R[280][1];				r_cell_reg[281] = inform_R[282][1];				r_cell_reg[282] = inform_R[281][1];				r_cell_reg[283] = inform_R[283][1];				r_cell_reg[284] = inform_R[284][1];				r_cell_reg[285] = inform_R[286][1];				r_cell_reg[286] = inform_R[285][1];				r_cell_reg[287] = inform_R[287][1];				r_cell_reg[288] = inform_R[288][1];				r_cell_reg[289] = inform_R[290][1];				r_cell_reg[290] = inform_R[289][1];				r_cell_reg[291] = inform_R[291][1];				r_cell_reg[292] = inform_R[292][1];				r_cell_reg[293] = inform_R[294][1];				r_cell_reg[294] = inform_R[293][1];				r_cell_reg[295] = inform_R[295][1];				r_cell_reg[296] = inform_R[296][1];				r_cell_reg[297] = inform_R[298][1];				r_cell_reg[298] = inform_R[297][1];				r_cell_reg[299] = inform_R[299][1];				r_cell_reg[300] = inform_R[300][1];				r_cell_reg[301] = inform_R[302][1];				r_cell_reg[302] = inform_R[301][1];				r_cell_reg[303] = inform_R[303][1];				r_cell_reg[304] = inform_R[304][1];				r_cell_reg[305] = inform_R[306][1];				r_cell_reg[306] = inform_R[305][1];				r_cell_reg[307] = inform_R[307][1];				r_cell_reg[308] = inform_R[308][1];				r_cell_reg[309] = inform_R[310][1];				r_cell_reg[310] = inform_R[309][1];				r_cell_reg[311] = inform_R[311][1];				r_cell_reg[312] = inform_R[312][1];				r_cell_reg[313] = inform_R[314][1];				r_cell_reg[314] = inform_R[313][1];				r_cell_reg[315] = inform_R[315][1];				r_cell_reg[316] = inform_R[316][1];				r_cell_reg[317] = inform_R[318][1];				r_cell_reg[318] = inform_R[317][1];				r_cell_reg[319] = inform_R[319][1];				r_cell_reg[320] = inform_R[320][1];				r_cell_reg[321] = inform_R[322][1];				r_cell_reg[322] = inform_R[321][1];				r_cell_reg[323] = inform_R[323][1];				r_cell_reg[324] = inform_R[324][1];				r_cell_reg[325] = inform_R[326][1];				r_cell_reg[326] = inform_R[325][1];				r_cell_reg[327] = inform_R[327][1];				r_cell_reg[328] = inform_R[328][1];				r_cell_reg[329] = inform_R[330][1];				r_cell_reg[330] = inform_R[329][1];				r_cell_reg[331] = inform_R[331][1];				r_cell_reg[332] = inform_R[332][1];				r_cell_reg[333] = inform_R[334][1];				r_cell_reg[334] = inform_R[333][1];				r_cell_reg[335] = inform_R[335][1];				r_cell_reg[336] = inform_R[336][1];				r_cell_reg[337] = inform_R[338][1];				r_cell_reg[338] = inform_R[337][1];				r_cell_reg[339] = inform_R[339][1];				r_cell_reg[340] = inform_R[340][1];				r_cell_reg[341] = inform_R[342][1];				r_cell_reg[342] = inform_R[341][1];				r_cell_reg[343] = inform_R[343][1];				r_cell_reg[344] = inform_R[344][1];				r_cell_reg[345] = inform_R[346][1];				r_cell_reg[346] = inform_R[345][1];				r_cell_reg[347] = inform_R[347][1];				r_cell_reg[348] = inform_R[348][1];				r_cell_reg[349] = inform_R[350][1];				r_cell_reg[350] = inform_R[349][1];				r_cell_reg[351] = inform_R[351][1];				r_cell_reg[352] = inform_R[352][1];				r_cell_reg[353] = inform_R[354][1];				r_cell_reg[354] = inform_R[353][1];				r_cell_reg[355] = inform_R[355][1];				r_cell_reg[356] = inform_R[356][1];				r_cell_reg[357] = inform_R[358][1];				r_cell_reg[358] = inform_R[357][1];				r_cell_reg[359] = inform_R[359][1];				r_cell_reg[360] = inform_R[360][1];				r_cell_reg[361] = inform_R[362][1];				r_cell_reg[362] = inform_R[361][1];				r_cell_reg[363] = inform_R[363][1];				r_cell_reg[364] = inform_R[364][1];				r_cell_reg[365] = inform_R[366][1];				r_cell_reg[366] = inform_R[365][1];				r_cell_reg[367] = inform_R[367][1];				r_cell_reg[368] = inform_R[368][1];				r_cell_reg[369] = inform_R[370][1];				r_cell_reg[370] = inform_R[369][1];				r_cell_reg[371] = inform_R[371][1];				r_cell_reg[372] = inform_R[372][1];				r_cell_reg[373] = inform_R[374][1];				r_cell_reg[374] = inform_R[373][1];				r_cell_reg[375] = inform_R[375][1];				r_cell_reg[376] = inform_R[376][1];				r_cell_reg[377] = inform_R[378][1];				r_cell_reg[378] = inform_R[377][1];				r_cell_reg[379] = inform_R[379][1];				r_cell_reg[380] = inform_R[380][1];				r_cell_reg[381] = inform_R[382][1];				r_cell_reg[382] = inform_R[381][1];				r_cell_reg[383] = inform_R[383][1];				r_cell_reg[384] = inform_R[384][1];				r_cell_reg[385] = inform_R[386][1];				r_cell_reg[386] = inform_R[385][1];				r_cell_reg[387] = inform_R[387][1];				r_cell_reg[388] = inform_R[388][1];				r_cell_reg[389] = inform_R[390][1];				r_cell_reg[390] = inform_R[389][1];				r_cell_reg[391] = inform_R[391][1];				r_cell_reg[392] = inform_R[392][1];				r_cell_reg[393] = inform_R[394][1];				r_cell_reg[394] = inform_R[393][1];				r_cell_reg[395] = inform_R[395][1];				r_cell_reg[396] = inform_R[396][1];				r_cell_reg[397] = inform_R[398][1];				r_cell_reg[398] = inform_R[397][1];				r_cell_reg[399] = inform_R[399][1];				r_cell_reg[400] = inform_R[400][1];				r_cell_reg[401] = inform_R[402][1];				r_cell_reg[402] = inform_R[401][1];				r_cell_reg[403] = inform_R[403][1];				r_cell_reg[404] = inform_R[404][1];				r_cell_reg[405] = inform_R[406][1];				r_cell_reg[406] = inform_R[405][1];				r_cell_reg[407] = inform_R[407][1];				r_cell_reg[408] = inform_R[408][1];				r_cell_reg[409] = inform_R[410][1];				r_cell_reg[410] = inform_R[409][1];				r_cell_reg[411] = inform_R[411][1];				r_cell_reg[412] = inform_R[412][1];				r_cell_reg[413] = inform_R[414][1];				r_cell_reg[414] = inform_R[413][1];				r_cell_reg[415] = inform_R[415][1];				r_cell_reg[416] = inform_R[416][1];				r_cell_reg[417] = inform_R[418][1];				r_cell_reg[418] = inform_R[417][1];				r_cell_reg[419] = inform_R[419][1];				r_cell_reg[420] = inform_R[420][1];				r_cell_reg[421] = inform_R[422][1];				r_cell_reg[422] = inform_R[421][1];				r_cell_reg[423] = inform_R[423][1];				r_cell_reg[424] = inform_R[424][1];				r_cell_reg[425] = inform_R[426][1];				r_cell_reg[426] = inform_R[425][1];				r_cell_reg[427] = inform_R[427][1];				r_cell_reg[428] = inform_R[428][1];				r_cell_reg[429] = inform_R[430][1];				r_cell_reg[430] = inform_R[429][1];				r_cell_reg[431] = inform_R[431][1];				r_cell_reg[432] = inform_R[432][1];				r_cell_reg[433] = inform_R[434][1];				r_cell_reg[434] = inform_R[433][1];				r_cell_reg[435] = inform_R[435][1];				r_cell_reg[436] = inform_R[436][1];				r_cell_reg[437] = inform_R[438][1];				r_cell_reg[438] = inform_R[437][1];				r_cell_reg[439] = inform_R[439][1];				r_cell_reg[440] = inform_R[440][1];				r_cell_reg[441] = inform_R[442][1];				r_cell_reg[442] = inform_R[441][1];				r_cell_reg[443] = inform_R[443][1];				r_cell_reg[444] = inform_R[444][1];				r_cell_reg[445] = inform_R[446][1];				r_cell_reg[446] = inform_R[445][1];				r_cell_reg[447] = inform_R[447][1];				r_cell_reg[448] = inform_R[448][1];				r_cell_reg[449] = inform_R[450][1];				r_cell_reg[450] = inform_R[449][1];				r_cell_reg[451] = inform_R[451][1];				r_cell_reg[452] = inform_R[452][1];				r_cell_reg[453] = inform_R[454][1];				r_cell_reg[454] = inform_R[453][1];				r_cell_reg[455] = inform_R[455][1];				r_cell_reg[456] = inform_R[456][1];				r_cell_reg[457] = inform_R[458][1];				r_cell_reg[458] = inform_R[457][1];				r_cell_reg[459] = inform_R[459][1];				r_cell_reg[460] = inform_R[460][1];				r_cell_reg[461] = inform_R[462][1];				r_cell_reg[462] = inform_R[461][1];				r_cell_reg[463] = inform_R[463][1];				r_cell_reg[464] = inform_R[464][1];				r_cell_reg[465] = inform_R[466][1];				r_cell_reg[466] = inform_R[465][1];				r_cell_reg[467] = inform_R[467][1];				r_cell_reg[468] = inform_R[468][1];				r_cell_reg[469] = inform_R[470][1];				r_cell_reg[470] = inform_R[469][1];				r_cell_reg[471] = inform_R[471][1];				r_cell_reg[472] = inform_R[472][1];				r_cell_reg[473] = inform_R[474][1];				r_cell_reg[474] = inform_R[473][1];				r_cell_reg[475] = inform_R[475][1];				r_cell_reg[476] = inform_R[476][1];				r_cell_reg[477] = inform_R[478][1];				r_cell_reg[478] = inform_R[477][1];				r_cell_reg[479] = inform_R[479][1];				r_cell_reg[480] = inform_R[480][1];				r_cell_reg[481] = inform_R[482][1];				r_cell_reg[482] = inform_R[481][1];				r_cell_reg[483] = inform_R[483][1];				r_cell_reg[484] = inform_R[484][1];				r_cell_reg[485] = inform_R[486][1];				r_cell_reg[486] = inform_R[485][1];				r_cell_reg[487] = inform_R[487][1];				r_cell_reg[488] = inform_R[488][1];				r_cell_reg[489] = inform_R[490][1];				r_cell_reg[490] = inform_R[489][1];				r_cell_reg[491] = inform_R[491][1];				r_cell_reg[492] = inform_R[492][1];				r_cell_reg[493] = inform_R[494][1];				r_cell_reg[494] = inform_R[493][1];				r_cell_reg[495] = inform_R[495][1];				r_cell_reg[496] = inform_R[496][1];				r_cell_reg[497] = inform_R[498][1];				r_cell_reg[498] = inform_R[497][1];				r_cell_reg[499] = inform_R[499][1];				r_cell_reg[500] = inform_R[500][1];				r_cell_reg[501] = inform_R[502][1];				r_cell_reg[502] = inform_R[501][1];				r_cell_reg[503] = inform_R[503][1];				r_cell_reg[504] = inform_R[504][1];				r_cell_reg[505] = inform_R[506][1];				r_cell_reg[506] = inform_R[505][1];				r_cell_reg[507] = inform_R[507][1];				r_cell_reg[508] = inform_R[508][1];				r_cell_reg[509] = inform_R[510][1];				r_cell_reg[510] = inform_R[509][1];				r_cell_reg[511] = inform_R[511][1];				r_cell_reg[512] = inform_R[512][1];				r_cell_reg[513] = inform_R[514][1];				r_cell_reg[514] = inform_R[513][1];				r_cell_reg[515] = inform_R[515][1];				r_cell_reg[516] = inform_R[516][1];				r_cell_reg[517] = inform_R[518][1];				r_cell_reg[518] = inform_R[517][1];				r_cell_reg[519] = inform_R[519][1];				r_cell_reg[520] = inform_R[520][1];				r_cell_reg[521] = inform_R[522][1];				r_cell_reg[522] = inform_R[521][1];				r_cell_reg[523] = inform_R[523][1];				r_cell_reg[524] = inform_R[524][1];				r_cell_reg[525] = inform_R[526][1];				r_cell_reg[526] = inform_R[525][1];				r_cell_reg[527] = inform_R[527][1];				r_cell_reg[528] = inform_R[528][1];				r_cell_reg[529] = inform_R[530][1];				r_cell_reg[530] = inform_R[529][1];				r_cell_reg[531] = inform_R[531][1];				r_cell_reg[532] = inform_R[532][1];				r_cell_reg[533] = inform_R[534][1];				r_cell_reg[534] = inform_R[533][1];				r_cell_reg[535] = inform_R[535][1];				r_cell_reg[536] = inform_R[536][1];				r_cell_reg[537] = inform_R[538][1];				r_cell_reg[538] = inform_R[537][1];				r_cell_reg[539] = inform_R[539][1];				r_cell_reg[540] = inform_R[540][1];				r_cell_reg[541] = inform_R[542][1];				r_cell_reg[542] = inform_R[541][1];				r_cell_reg[543] = inform_R[543][1];				r_cell_reg[544] = inform_R[544][1];				r_cell_reg[545] = inform_R[546][1];				r_cell_reg[546] = inform_R[545][1];				r_cell_reg[547] = inform_R[547][1];				r_cell_reg[548] = inform_R[548][1];				r_cell_reg[549] = inform_R[550][1];				r_cell_reg[550] = inform_R[549][1];				r_cell_reg[551] = inform_R[551][1];				r_cell_reg[552] = inform_R[552][1];				r_cell_reg[553] = inform_R[554][1];				r_cell_reg[554] = inform_R[553][1];				r_cell_reg[555] = inform_R[555][1];				r_cell_reg[556] = inform_R[556][1];				r_cell_reg[557] = inform_R[558][1];				r_cell_reg[558] = inform_R[557][1];				r_cell_reg[559] = inform_R[559][1];				r_cell_reg[560] = inform_R[560][1];				r_cell_reg[561] = inform_R[562][1];				r_cell_reg[562] = inform_R[561][1];				r_cell_reg[563] = inform_R[563][1];				r_cell_reg[564] = inform_R[564][1];				r_cell_reg[565] = inform_R[566][1];				r_cell_reg[566] = inform_R[565][1];				r_cell_reg[567] = inform_R[567][1];				r_cell_reg[568] = inform_R[568][1];				r_cell_reg[569] = inform_R[570][1];				r_cell_reg[570] = inform_R[569][1];				r_cell_reg[571] = inform_R[571][1];				r_cell_reg[572] = inform_R[572][1];				r_cell_reg[573] = inform_R[574][1];				r_cell_reg[574] = inform_R[573][1];				r_cell_reg[575] = inform_R[575][1];				r_cell_reg[576] = inform_R[576][1];				r_cell_reg[577] = inform_R[578][1];				r_cell_reg[578] = inform_R[577][1];				r_cell_reg[579] = inform_R[579][1];				r_cell_reg[580] = inform_R[580][1];				r_cell_reg[581] = inform_R[582][1];				r_cell_reg[582] = inform_R[581][1];				r_cell_reg[583] = inform_R[583][1];				r_cell_reg[584] = inform_R[584][1];				r_cell_reg[585] = inform_R[586][1];				r_cell_reg[586] = inform_R[585][1];				r_cell_reg[587] = inform_R[587][1];				r_cell_reg[588] = inform_R[588][1];				r_cell_reg[589] = inform_R[590][1];				r_cell_reg[590] = inform_R[589][1];				r_cell_reg[591] = inform_R[591][1];				r_cell_reg[592] = inform_R[592][1];				r_cell_reg[593] = inform_R[594][1];				r_cell_reg[594] = inform_R[593][1];				r_cell_reg[595] = inform_R[595][1];				r_cell_reg[596] = inform_R[596][1];				r_cell_reg[597] = inform_R[598][1];				r_cell_reg[598] = inform_R[597][1];				r_cell_reg[599] = inform_R[599][1];				r_cell_reg[600] = inform_R[600][1];				r_cell_reg[601] = inform_R[602][1];				r_cell_reg[602] = inform_R[601][1];				r_cell_reg[603] = inform_R[603][1];				r_cell_reg[604] = inform_R[604][1];				r_cell_reg[605] = inform_R[606][1];				r_cell_reg[606] = inform_R[605][1];				r_cell_reg[607] = inform_R[607][1];				r_cell_reg[608] = inform_R[608][1];				r_cell_reg[609] = inform_R[610][1];				r_cell_reg[610] = inform_R[609][1];				r_cell_reg[611] = inform_R[611][1];				r_cell_reg[612] = inform_R[612][1];				r_cell_reg[613] = inform_R[614][1];				r_cell_reg[614] = inform_R[613][1];				r_cell_reg[615] = inform_R[615][1];				r_cell_reg[616] = inform_R[616][1];				r_cell_reg[617] = inform_R[618][1];				r_cell_reg[618] = inform_R[617][1];				r_cell_reg[619] = inform_R[619][1];				r_cell_reg[620] = inform_R[620][1];				r_cell_reg[621] = inform_R[622][1];				r_cell_reg[622] = inform_R[621][1];				r_cell_reg[623] = inform_R[623][1];				r_cell_reg[624] = inform_R[624][1];				r_cell_reg[625] = inform_R[626][1];				r_cell_reg[626] = inform_R[625][1];				r_cell_reg[627] = inform_R[627][1];				r_cell_reg[628] = inform_R[628][1];				r_cell_reg[629] = inform_R[630][1];				r_cell_reg[630] = inform_R[629][1];				r_cell_reg[631] = inform_R[631][1];				r_cell_reg[632] = inform_R[632][1];				r_cell_reg[633] = inform_R[634][1];				r_cell_reg[634] = inform_R[633][1];				r_cell_reg[635] = inform_R[635][1];				r_cell_reg[636] = inform_R[636][1];				r_cell_reg[637] = inform_R[638][1];				r_cell_reg[638] = inform_R[637][1];				r_cell_reg[639] = inform_R[639][1];				r_cell_reg[640] = inform_R[640][1];				r_cell_reg[641] = inform_R[642][1];				r_cell_reg[642] = inform_R[641][1];				r_cell_reg[643] = inform_R[643][1];				r_cell_reg[644] = inform_R[644][1];				r_cell_reg[645] = inform_R[646][1];				r_cell_reg[646] = inform_R[645][1];				r_cell_reg[647] = inform_R[647][1];				r_cell_reg[648] = inform_R[648][1];				r_cell_reg[649] = inform_R[650][1];				r_cell_reg[650] = inform_R[649][1];				r_cell_reg[651] = inform_R[651][1];				r_cell_reg[652] = inform_R[652][1];				r_cell_reg[653] = inform_R[654][1];				r_cell_reg[654] = inform_R[653][1];				r_cell_reg[655] = inform_R[655][1];				r_cell_reg[656] = inform_R[656][1];				r_cell_reg[657] = inform_R[658][1];				r_cell_reg[658] = inform_R[657][1];				r_cell_reg[659] = inform_R[659][1];				r_cell_reg[660] = inform_R[660][1];				r_cell_reg[661] = inform_R[662][1];				r_cell_reg[662] = inform_R[661][1];				r_cell_reg[663] = inform_R[663][1];				r_cell_reg[664] = inform_R[664][1];				r_cell_reg[665] = inform_R[666][1];				r_cell_reg[666] = inform_R[665][1];				r_cell_reg[667] = inform_R[667][1];				r_cell_reg[668] = inform_R[668][1];				r_cell_reg[669] = inform_R[670][1];				r_cell_reg[670] = inform_R[669][1];				r_cell_reg[671] = inform_R[671][1];				r_cell_reg[672] = inform_R[672][1];				r_cell_reg[673] = inform_R[674][1];				r_cell_reg[674] = inform_R[673][1];				r_cell_reg[675] = inform_R[675][1];				r_cell_reg[676] = inform_R[676][1];				r_cell_reg[677] = inform_R[678][1];				r_cell_reg[678] = inform_R[677][1];				r_cell_reg[679] = inform_R[679][1];				r_cell_reg[680] = inform_R[680][1];				r_cell_reg[681] = inform_R[682][1];				r_cell_reg[682] = inform_R[681][1];				r_cell_reg[683] = inform_R[683][1];				r_cell_reg[684] = inform_R[684][1];				r_cell_reg[685] = inform_R[686][1];				r_cell_reg[686] = inform_R[685][1];				r_cell_reg[687] = inform_R[687][1];				r_cell_reg[688] = inform_R[688][1];				r_cell_reg[689] = inform_R[690][1];				r_cell_reg[690] = inform_R[689][1];				r_cell_reg[691] = inform_R[691][1];				r_cell_reg[692] = inform_R[692][1];				r_cell_reg[693] = inform_R[694][1];				r_cell_reg[694] = inform_R[693][1];				r_cell_reg[695] = inform_R[695][1];				r_cell_reg[696] = inform_R[696][1];				r_cell_reg[697] = inform_R[698][1];				r_cell_reg[698] = inform_R[697][1];				r_cell_reg[699] = inform_R[699][1];				r_cell_reg[700] = inform_R[700][1];				r_cell_reg[701] = inform_R[702][1];				r_cell_reg[702] = inform_R[701][1];				r_cell_reg[703] = inform_R[703][1];				r_cell_reg[704] = inform_R[704][1];				r_cell_reg[705] = inform_R[706][1];				r_cell_reg[706] = inform_R[705][1];				r_cell_reg[707] = inform_R[707][1];				r_cell_reg[708] = inform_R[708][1];				r_cell_reg[709] = inform_R[710][1];				r_cell_reg[710] = inform_R[709][1];				r_cell_reg[711] = inform_R[711][1];				r_cell_reg[712] = inform_R[712][1];				r_cell_reg[713] = inform_R[714][1];				r_cell_reg[714] = inform_R[713][1];				r_cell_reg[715] = inform_R[715][1];				r_cell_reg[716] = inform_R[716][1];				r_cell_reg[717] = inform_R[718][1];				r_cell_reg[718] = inform_R[717][1];				r_cell_reg[719] = inform_R[719][1];				r_cell_reg[720] = inform_R[720][1];				r_cell_reg[721] = inform_R[722][1];				r_cell_reg[722] = inform_R[721][1];				r_cell_reg[723] = inform_R[723][1];				r_cell_reg[724] = inform_R[724][1];				r_cell_reg[725] = inform_R[726][1];				r_cell_reg[726] = inform_R[725][1];				r_cell_reg[727] = inform_R[727][1];				r_cell_reg[728] = inform_R[728][1];				r_cell_reg[729] = inform_R[730][1];				r_cell_reg[730] = inform_R[729][1];				r_cell_reg[731] = inform_R[731][1];				r_cell_reg[732] = inform_R[732][1];				r_cell_reg[733] = inform_R[734][1];				r_cell_reg[734] = inform_R[733][1];				r_cell_reg[735] = inform_R[735][1];				r_cell_reg[736] = inform_R[736][1];				r_cell_reg[737] = inform_R[738][1];				r_cell_reg[738] = inform_R[737][1];				r_cell_reg[739] = inform_R[739][1];				r_cell_reg[740] = inform_R[740][1];				r_cell_reg[741] = inform_R[742][1];				r_cell_reg[742] = inform_R[741][1];				r_cell_reg[743] = inform_R[743][1];				r_cell_reg[744] = inform_R[744][1];				r_cell_reg[745] = inform_R[746][1];				r_cell_reg[746] = inform_R[745][1];				r_cell_reg[747] = inform_R[747][1];				r_cell_reg[748] = inform_R[748][1];				r_cell_reg[749] = inform_R[750][1];				r_cell_reg[750] = inform_R[749][1];				r_cell_reg[751] = inform_R[751][1];				r_cell_reg[752] = inform_R[752][1];				r_cell_reg[753] = inform_R[754][1];				r_cell_reg[754] = inform_R[753][1];				r_cell_reg[755] = inform_R[755][1];				r_cell_reg[756] = inform_R[756][1];				r_cell_reg[757] = inform_R[758][1];				r_cell_reg[758] = inform_R[757][1];				r_cell_reg[759] = inform_R[759][1];				r_cell_reg[760] = inform_R[760][1];				r_cell_reg[761] = inform_R[762][1];				r_cell_reg[762] = inform_R[761][1];				r_cell_reg[763] = inform_R[763][1];				r_cell_reg[764] = inform_R[764][1];				r_cell_reg[765] = inform_R[766][1];				r_cell_reg[766] = inform_R[765][1];				r_cell_reg[767] = inform_R[767][1];				r_cell_reg[768] = inform_R[768][1];				r_cell_reg[769] = inform_R[770][1];				r_cell_reg[770] = inform_R[769][1];				r_cell_reg[771] = inform_R[771][1];				r_cell_reg[772] = inform_R[772][1];				r_cell_reg[773] = inform_R[774][1];				r_cell_reg[774] = inform_R[773][1];				r_cell_reg[775] = inform_R[775][1];				r_cell_reg[776] = inform_R[776][1];				r_cell_reg[777] = inform_R[778][1];				r_cell_reg[778] = inform_R[777][1];				r_cell_reg[779] = inform_R[779][1];				r_cell_reg[780] = inform_R[780][1];				r_cell_reg[781] = inform_R[782][1];				r_cell_reg[782] = inform_R[781][1];				r_cell_reg[783] = inform_R[783][1];				r_cell_reg[784] = inform_R[784][1];				r_cell_reg[785] = inform_R[786][1];				r_cell_reg[786] = inform_R[785][1];				r_cell_reg[787] = inform_R[787][1];				r_cell_reg[788] = inform_R[788][1];				r_cell_reg[789] = inform_R[790][1];				r_cell_reg[790] = inform_R[789][1];				r_cell_reg[791] = inform_R[791][1];				r_cell_reg[792] = inform_R[792][1];				r_cell_reg[793] = inform_R[794][1];				r_cell_reg[794] = inform_R[793][1];				r_cell_reg[795] = inform_R[795][1];				r_cell_reg[796] = inform_R[796][1];				r_cell_reg[797] = inform_R[798][1];				r_cell_reg[798] = inform_R[797][1];				r_cell_reg[799] = inform_R[799][1];				r_cell_reg[800] = inform_R[800][1];				r_cell_reg[801] = inform_R[802][1];				r_cell_reg[802] = inform_R[801][1];				r_cell_reg[803] = inform_R[803][1];				r_cell_reg[804] = inform_R[804][1];				r_cell_reg[805] = inform_R[806][1];				r_cell_reg[806] = inform_R[805][1];				r_cell_reg[807] = inform_R[807][1];				r_cell_reg[808] = inform_R[808][1];				r_cell_reg[809] = inform_R[810][1];				r_cell_reg[810] = inform_R[809][1];				r_cell_reg[811] = inform_R[811][1];				r_cell_reg[812] = inform_R[812][1];				r_cell_reg[813] = inform_R[814][1];				r_cell_reg[814] = inform_R[813][1];				r_cell_reg[815] = inform_R[815][1];				r_cell_reg[816] = inform_R[816][1];				r_cell_reg[817] = inform_R[818][1];				r_cell_reg[818] = inform_R[817][1];				r_cell_reg[819] = inform_R[819][1];				r_cell_reg[820] = inform_R[820][1];				r_cell_reg[821] = inform_R[822][1];				r_cell_reg[822] = inform_R[821][1];				r_cell_reg[823] = inform_R[823][1];				r_cell_reg[824] = inform_R[824][1];				r_cell_reg[825] = inform_R[826][1];				r_cell_reg[826] = inform_R[825][1];				r_cell_reg[827] = inform_R[827][1];				r_cell_reg[828] = inform_R[828][1];				r_cell_reg[829] = inform_R[830][1];				r_cell_reg[830] = inform_R[829][1];				r_cell_reg[831] = inform_R[831][1];				r_cell_reg[832] = inform_R[832][1];				r_cell_reg[833] = inform_R[834][1];				r_cell_reg[834] = inform_R[833][1];				r_cell_reg[835] = inform_R[835][1];				r_cell_reg[836] = inform_R[836][1];				r_cell_reg[837] = inform_R[838][1];				r_cell_reg[838] = inform_R[837][1];				r_cell_reg[839] = inform_R[839][1];				r_cell_reg[840] = inform_R[840][1];				r_cell_reg[841] = inform_R[842][1];				r_cell_reg[842] = inform_R[841][1];				r_cell_reg[843] = inform_R[843][1];				r_cell_reg[844] = inform_R[844][1];				r_cell_reg[845] = inform_R[846][1];				r_cell_reg[846] = inform_R[845][1];				r_cell_reg[847] = inform_R[847][1];				r_cell_reg[848] = inform_R[848][1];				r_cell_reg[849] = inform_R[850][1];				r_cell_reg[850] = inform_R[849][1];				r_cell_reg[851] = inform_R[851][1];				r_cell_reg[852] = inform_R[852][1];				r_cell_reg[853] = inform_R[854][1];				r_cell_reg[854] = inform_R[853][1];				r_cell_reg[855] = inform_R[855][1];				r_cell_reg[856] = inform_R[856][1];				r_cell_reg[857] = inform_R[858][1];				r_cell_reg[858] = inform_R[857][1];				r_cell_reg[859] = inform_R[859][1];				r_cell_reg[860] = inform_R[860][1];				r_cell_reg[861] = inform_R[862][1];				r_cell_reg[862] = inform_R[861][1];				r_cell_reg[863] = inform_R[863][1];				r_cell_reg[864] = inform_R[864][1];				r_cell_reg[865] = inform_R[866][1];				r_cell_reg[866] = inform_R[865][1];				r_cell_reg[867] = inform_R[867][1];				r_cell_reg[868] = inform_R[868][1];				r_cell_reg[869] = inform_R[870][1];				r_cell_reg[870] = inform_R[869][1];				r_cell_reg[871] = inform_R[871][1];				r_cell_reg[872] = inform_R[872][1];				r_cell_reg[873] = inform_R[874][1];				r_cell_reg[874] = inform_R[873][1];				r_cell_reg[875] = inform_R[875][1];				r_cell_reg[876] = inform_R[876][1];				r_cell_reg[877] = inform_R[878][1];				r_cell_reg[878] = inform_R[877][1];				r_cell_reg[879] = inform_R[879][1];				r_cell_reg[880] = inform_R[880][1];				r_cell_reg[881] = inform_R[882][1];				r_cell_reg[882] = inform_R[881][1];				r_cell_reg[883] = inform_R[883][1];				r_cell_reg[884] = inform_R[884][1];				r_cell_reg[885] = inform_R[886][1];				r_cell_reg[886] = inform_R[885][1];				r_cell_reg[887] = inform_R[887][1];				r_cell_reg[888] = inform_R[888][1];				r_cell_reg[889] = inform_R[890][1];				r_cell_reg[890] = inform_R[889][1];				r_cell_reg[891] = inform_R[891][1];				r_cell_reg[892] = inform_R[892][1];				r_cell_reg[893] = inform_R[894][1];				r_cell_reg[894] = inform_R[893][1];				r_cell_reg[895] = inform_R[895][1];				r_cell_reg[896] = inform_R[896][1];				r_cell_reg[897] = inform_R[898][1];				r_cell_reg[898] = inform_R[897][1];				r_cell_reg[899] = inform_R[899][1];				r_cell_reg[900] = inform_R[900][1];				r_cell_reg[901] = inform_R[902][1];				r_cell_reg[902] = inform_R[901][1];				r_cell_reg[903] = inform_R[903][1];				r_cell_reg[904] = inform_R[904][1];				r_cell_reg[905] = inform_R[906][1];				r_cell_reg[906] = inform_R[905][1];				r_cell_reg[907] = inform_R[907][1];				r_cell_reg[908] = inform_R[908][1];				r_cell_reg[909] = inform_R[910][1];				r_cell_reg[910] = inform_R[909][1];				r_cell_reg[911] = inform_R[911][1];				r_cell_reg[912] = inform_R[912][1];				r_cell_reg[913] = inform_R[914][1];				r_cell_reg[914] = inform_R[913][1];				r_cell_reg[915] = inform_R[915][1];				r_cell_reg[916] = inform_R[916][1];				r_cell_reg[917] = inform_R[918][1];				r_cell_reg[918] = inform_R[917][1];				r_cell_reg[919] = inform_R[919][1];				r_cell_reg[920] = inform_R[920][1];				r_cell_reg[921] = inform_R[922][1];				r_cell_reg[922] = inform_R[921][1];				r_cell_reg[923] = inform_R[923][1];				r_cell_reg[924] = inform_R[924][1];				r_cell_reg[925] = inform_R[926][1];				r_cell_reg[926] = inform_R[925][1];				r_cell_reg[927] = inform_R[927][1];				r_cell_reg[928] = inform_R[928][1];				r_cell_reg[929] = inform_R[930][1];				r_cell_reg[930] = inform_R[929][1];				r_cell_reg[931] = inform_R[931][1];				r_cell_reg[932] = inform_R[932][1];				r_cell_reg[933] = inform_R[934][1];				r_cell_reg[934] = inform_R[933][1];				r_cell_reg[935] = inform_R[935][1];				r_cell_reg[936] = inform_R[936][1];				r_cell_reg[937] = inform_R[938][1];				r_cell_reg[938] = inform_R[937][1];				r_cell_reg[939] = inform_R[939][1];				r_cell_reg[940] = inform_R[940][1];				r_cell_reg[941] = inform_R[942][1];				r_cell_reg[942] = inform_R[941][1];				r_cell_reg[943] = inform_R[943][1];				r_cell_reg[944] = inform_R[944][1];				r_cell_reg[945] = inform_R[946][1];				r_cell_reg[946] = inform_R[945][1];				r_cell_reg[947] = inform_R[947][1];				r_cell_reg[948] = inform_R[948][1];				r_cell_reg[949] = inform_R[950][1];				r_cell_reg[950] = inform_R[949][1];				r_cell_reg[951] = inform_R[951][1];				r_cell_reg[952] = inform_R[952][1];				r_cell_reg[953] = inform_R[954][1];				r_cell_reg[954] = inform_R[953][1];				r_cell_reg[955] = inform_R[955][1];				r_cell_reg[956] = inform_R[956][1];				r_cell_reg[957] = inform_R[958][1];				r_cell_reg[958] = inform_R[957][1];				r_cell_reg[959] = inform_R[959][1];				r_cell_reg[960] = inform_R[960][1];				r_cell_reg[961] = inform_R[962][1];				r_cell_reg[962] = inform_R[961][1];				r_cell_reg[963] = inform_R[963][1];				r_cell_reg[964] = inform_R[964][1];				r_cell_reg[965] = inform_R[966][1];				r_cell_reg[966] = inform_R[965][1];				r_cell_reg[967] = inform_R[967][1];				r_cell_reg[968] = inform_R[968][1];				r_cell_reg[969] = inform_R[970][1];				r_cell_reg[970] = inform_R[969][1];				r_cell_reg[971] = inform_R[971][1];				r_cell_reg[972] = inform_R[972][1];				r_cell_reg[973] = inform_R[974][1];				r_cell_reg[974] = inform_R[973][1];				r_cell_reg[975] = inform_R[975][1];				r_cell_reg[976] = inform_R[976][1];				r_cell_reg[977] = inform_R[978][1];				r_cell_reg[978] = inform_R[977][1];				r_cell_reg[979] = inform_R[979][1];				r_cell_reg[980] = inform_R[980][1];				r_cell_reg[981] = inform_R[982][1];				r_cell_reg[982] = inform_R[981][1];				r_cell_reg[983] = inform_R[983][1];				r_cell_reg[984] = inform_R[984][1];				r_cell_reg[985] = inform_R[986][1];				r_cell_reg[986] = inform_R[985][1];				r_cell_reg[987] = inform_R[987][1];				r_cell_reg[988] = inform_R[988][1];				r_cell_reg[989] = inform_R[990][1];				r_cell_reg[990] = inform_R[989][1];				r_cell_reg[991] = inform_R[991][1];				r_cell_reg[992] = inform_R[992][1];				r_cell_reg[993] = inform_R[994][1];				r_cell_reg[994] = inform_R[993][1];				r_cell_reg[995] = inform_R[995][1];				r_cell_reg[996] = inform_R[996][1];				r_cell_reg[997] = inform_R[998][1];				r_cell_reg[998] = inform_R[997][1];				r_cell_reg[999] = inform_R[999][1];				r_cell_reg[1000] = inform_R[1000][1];				r_cell_reg[1001] = inform_R[1002][1];				r_cell_reg[1002] = inform_R[1001][1];				r_cell_reg[1003] = inform_R[1003][1];				r_cell_reg[1004] = inform_R[1004][1];				r_cell_reg[1005] = inform_R[1006][1];				r_cell_reg[1006] = inform_R[1005][1];				r_cell_reg[1007] = inform_R[1007][1];				r_cell_reg[1008] = inform_R[1008][1];				r_cell_reg[1009] = inform_R[1010][1];				r_cell_reg[1010] = inform_R[1009][1];				r_cell_reg[1011] = inform_R[1011][1];				r_cell_reg[1012] = inform_R[1012][1];				r_cell_reg[1013] = inform_R[1014][1];				r_cell_reg[1014] = inform_R[1013][1];				r_cell_reg[1015] = inform_R[1015][1];				r_cell_reg[1016] = inform_R[1016][1];				r_cell_reg[1017] = inform_R[1018][1];				r_cell_reg[1018] = inform_R[1017][1];				r_cell_reg[1019] = inform_R[1019][1];				r_cell_reg[1020] = inform_R[1020][1];				r_cell_reg[1021] = inform_R[1022][1];				r_cell_reg[1022] = inform_R[1021][1];				r_cell_reg[1023] = inform_R[1023][1];				l_cell_reg[0] = inform_L[0][2];				l_cell_reg[1] = inform_L[2][2];				l_cell_reg[2] = inform_L[1][2];				l_cell_reg[3] = inform_L[3][2];				l_cell_reg[4] = inform_L[4][2];				l_cell_reg[5] = inform_L[6][2];				l_cell_reg[6] = inform_L[5][2];				l_cell_reg[7] = inform_L[7][2];				l_cell_reg[8] = inform_L[8][2];				l_cell_reg[9] = inform_L[10][2];				l_cell_reg[10] = inform_L[9][2];				l_cell_reg[11] = inform_L[11][2];				l_cell_reg[12] = inform_L[12][2];				l_cell_reg[13] = inform_L[14][2];				l_cell_reg[14] = inform_L[13][2];				l_cell_reg[15] = inform_L[15][2];				l_cell_reg[16] = inform_L[16][2];				l_cell_reg[17] = inform_L[18][2];				l_cell_reg[18] = inform_L[17][2];				l_cell_reg[19] = inform_L[19][2];				l_cell_reg[20] = inform_L[20][2];				l_cell_reg[21] = inform_L[22][2];				l_cell_reg[22] = inform_L[21][2];				l_cell_reg[23] = inform_L[23][2];				l_cell_reg[24] = inform_L[24][2];				l_cell_reg[25] = inform_L[26][2];				l_cell_reg[26] = inform_L[25][2];				l_cell_reg[27] = inform_L[27][2];				l_cell_reg[28] = inform_L[28][2];				l_cell_reg[29] = inform_L[30][2];				l_cell_reg[30] = inform_L[29][2];				l_cell_reg[31] = inform_L[31][2];				l_cell_reg[32] = inform_L[32][2];				l_cell_reg[33] = inform_L[34][2];				l_cell_reg[34] = inform_L[33][2];				l_cell_reg[35] = inform_L[35][2];				l_cell_reg[36] = inform_L[36][2];				l_cell_reg[37] = inform_L[38][2];				l_cell_reg[38] = inform_L[37][2];				l_cell_reg[39] = inform_L[39][2];				l_cell_reg[40] = inform_L[40][2];				l_cell_reg[41] = inform_L[42][2];				l_cell_reg[42] = inform_L[41][2];				l_cell_reg[43] = inform_L[43][2];				l_cell_reg[44] = inform_L[44][2];				l_cell_reg[45] = inform_L[46][2];				l_cell_reg[46] = inform_L[45][2];				l_cell_reg[47] = inform_L[47][2];				l_cell_reg[48] = inform_L[48][2];				l_cell_reg[49] = inform_L[50][2];				l_cell_reg[50] = inform_L[49][2];				l_cell_reg[51] = inform_L[51][2];				l_cell_reg[52] = inform_L[52][2];				l_cell_reg[53] = inform_L[54][2];				l_cell_reg[54] = inform_L[53][2];				l_cell_reg[55] = inform_L[55][2];				l_cell_reg[56] = inform_L[56][2];				l_cell_reg[57] = inform_L[58][2];				l_cell_reg[58] = inform_L[57][2];				l_cell_reg[59] = inform_L[59][2];				l_cell_reg[60] = inform_L[60][2];				l_cell_reg[61] = inform_L[62][2];				l_cell_reg[62] = inform_L[61][2];				l_cell_reg[63] = inform_L[63][2];				l_cell_reg[64] = inform_L[64][2];				l_cell_reg[65] = inform_L[66][2];				l_cell_reg[66] = inform_L[65][2];				l_cell_reg[67] = inform_L[67][2];				l_cell_reg[68] = inform_L[68][2];				l_cell_reg[69] = inform_L[70][2];				l_cell_reg[70] = inform_L[69][2];				l_cell_reg[71] = inform_L[71][2];				l_cell_reg[72] = inform_L[72][2];				l_cell_reg[73] = inform_L[74][2];				l_cell_reg[74] = inform_L[73][2];				l_cell_reg[75] = inform_L[75][2];				l_cell_reg[76] = inform_L[76][2];				l_cell_reg[77] = inform_L[78][2];				l_cell_reg[78] = inform_L[77][2];				l_cell_reg[79] = inform_L[79][2];				l_cell_reg[80] = inform_L[80][2];				l_cell_reg[81] = inform_L[82][2];				l_cell_reg[82] = inform_L[81][2];				l_cell_reg[83] = inform_L[83][2];				l_cell_reg[84] = inform_L[84][2];				l_cell_reg[85] = inform_L[86][2];				l_cell_reg[86] = inform_L[85][2];				l_cell_reg[87] = inform_L[87][2];				l_cell_reg[88] = inform_L[88][2];				l_cell_reg[89] = inform_L[90][2];				l_cell_reg[90] = inform_L[89][2];				l_cell_reg[91] = inform_L[91][2];				l_cell_reg[92] = inform_L[92][2];				l_cell_reg[93] = inform_L[94][2];				l_cell_reg[94] = inform_L[93][2];				l_cell_reg[95] = inform_L[95][2];				l_cell_reg[96] = inform_L[96][2];				l_cell_reg[97] = inform_L[98][2];				l_cell_reg[98] = inform_L[97][2];				l_cell_reg[99] = inform_L[99][2];				l_cell_reg[100] = inform_L[100][2];				l_cell_reg[101] = inform_L[102][2];				l_cell_reg[102] = inform_L[101][2];				l_cell_reg[103] = inform_L[103][2];				l_cell_reg[104] = inform_L[104][2];				l_cell_reg[105] = inform_L[106][2];				l_cell_reg[106] = inform_L[105][2];				l_cell_reg[107] = inform_L[107][2];				l_cell_reg[108] = inform_L[108][2];				l_cell_reg[109] = inform_L[110][2];				l_cell_reg[110] = inform_L[109][2];				l_cell_reg[111] = inform_L[111][2];				l_cell_reg[112] = inform_L[112][2];				l_cell_reg[113] = inform_L[114][2];				l_cell_reg[114] = inform_L[113][2];				l_cell_reg[115] = inform_L[115][2];				l_cell_reg[116] = inform_L[116][2];				l_cell_reg[117] = inform_L[118][2];				l_cell_reg[118] = inform_L[117][2];				l_cell_reg[119] = inform_L[119][2];				l_cell_reg[120] = inform_L[120][2];				l_cell_reg[121] = inform_L[122][2];				l_cell_reg[122] = inform_L[121][2];				l_cell_reg[123] = inform_L[123][2];				l_cell_reg[124] = inform_L[124][2];				l_cell_reg[125] = inform_L[126][2];				l_cell_reg[126] = inform_L[125][2];				l_cell_reg[127] = inform_L[127][2];				l_cell_reg[128] = inform_L[128][2];				l_cell_reg[129] = inform_L[130][2];				l_cell_reg[130] = inform_L[129][2];				l_cell_reg[131] = inform_L[131][2];				l_cell_reg[132] = inform_L[132][2];				l_cell_reg[133] = inform_L[134][2];				l_cell_reg[134] = inform_L[133][2];				l_cell_reg[135] = inform_L[135][2];				l_cell_reg[136] = inform_L[136][2];				l_cell_reg[137] = inform_L[138][2];				l_cell_reg[138] = inform_L[137][2];				l_cell_reg[139] = inform_L[139][2];				l_cell_reg[140] = inform_L[140][2];				l_cell_reg[141] = inform_L[142][2];				l_cell_reg[142] = inform_L[141][2];				l_cell_reg[143] = inform_L[143][2];				l_cell_reg[144] = inform_L[144][2];				l_cell_reg[145] = inform_L[146][2];				l_cell_reg[146] = inform_L[145][2];				l_cell_reg[147] = inform_L[147][2];				l_cell_reg[148] = inform_L[148][2];				l_cell_reg[149] = inform_L[150][2];				l_cell_reg[150] = inform_L[149][2];				l_cell_reg[151] = inform_L[151][2];				l_cell_reg[152] = inform_L[152][2];				l_cell_reg[153] = inform_L[154][2];				l_cell_reg[154] = inform_L[153][2];				l_cell_reg[155] = inform_L[155][2];				l_cell_reg[156] = inform_L[156][2];				l_cell_reg[157] = inform_L[158][2];				l_cell_reg[158] = inform_L[157][2];				l_cell_reg[159] = inform_L[159][2];				l_cell_reg[160] = inform_L[160][2];				l_cell_reg[161] = inform_L[162][2];				l_cell_reg[162] = inform_L[161][2];				l_cell_reg[163] = inform_L[163][2];				l_cell_reg[164] = inform_L[164][2];				l_cell_reg[165] = inform_L[166][2];				l_cell_reg[166] = inform_L[165][2];				l_cell_reg[167] = inform_L[167][2];				l_cell_reg[168] = inform_L[168][2];				l_cell_reg[169] = inform_L[170][2];				l_cell_reg[170] = inform_L[169][2];				l_cell_reg[171] = inform_L[171][2];				l_cell_reg[172] = inform_L[172][2];				l_cell_reg[173] = inform_L[174][2];				l_cell_reg[174] = inform_L[173][2];				l_cell_reg[175] = inform_L[175][2];				l_cell_reg[176] = inform_L[176][2];				l_cell_reg[177] = inform_L[178][2];				l_cell_reg[178] = inform_L[177][2];				l_cell_reg[179] = inform_L[179][2];				l_cell_reg[180] = inform_L[180][2];				l_cell_reg[181] = inform_L[182][2];				l_cell_reg[182] = inform_L[181][2];				l_cell_reg[183] = inform_L[183][2];				l_cell_reg[184] = inform_L[184][2];				l_cell_reg[185] = inform_L[186][2];				l_cell_reg[186] = inform_L[185][2];				l_cell_reg[187] = inform_L[187][2];				l_cell_reg[188] = inform_L[188][2];				l_cell_reg[189] = inform_L[190][2];				l_cell_reg[190] = inform_L[189][2];				l_cell_reg[191] = inform_L[191][2];				l_cell_reg[192] = inform_L[192][2];				l_cell_reg[193] = inform_L[194][2];				l_cell_reg[194] = inform_L[193][2];				l_cell_reg[195] = inform_L[195][2];				l_cell_reg[196] = inform_L[196][2];				l_cell_reg[197] = inform_L[198][2];				l_cell_reg[198] = inform_L[197][2];				l_cell_reg[199] = inform_L[199][2];				l_cell_reg[200] = inform_L[200][2];				l_cell_reg[201] = inform_L[202][2];				l_cell_reg[202] = inform_L[201][2];				l_cell_reg[203] = inform_L[203][2];				l_cell_reg[204] = inform_L[204][2];				l_cell_reg[205] = inform_L[206][2];				l_cell_reg[206] = inform_L[205][2];				l_cell_reg[207] = inform_L[207][2];				l_cell_reg[208] = inform_L[208][2];				l_cell_reg[209] = inform_L[210][2];				l_cell_reg[210] = inform_L[209][2];				l_cell_reg[211] = inform_L[211][2];				l_cell_reg[212] = inform_L[212][2];				l_cell_reg[213] = inform_L[214][2];				l_cell_reg[214] = inform_L[213][2];				l_cell_reg[215] = inform_L[215][2];				l_cell_reg[216] = inform_L[216][2];				l_cell_reg[217] = inform_L[218][2];				l_cell_reg[218] = inform_L[217][2];				l_cell_reg[219] = inform_L[219][2];				l_cell_reg[220] = inform_L[220][2];				l_cell_reg[221] = inform_L[222][2];				l_cell_reg[222] = inform_L[221][2];				l_cell_reg[223] = inform_L[223][2];				l_cell_reg[224] = inform_L[224][2];				l_cell_reg[225] = inform_L[226][2];				l_cell_reg[226] = inform_L[225][2];				l_cell_reg[227] = inform_L[227][2];				l_cell_reg[228] = inform_L[228][2];				l_cell_reg[229] = inform_L[230][2];				l_cell_reg[230] = inform_L[229][2];				l_cell_reg[231] = inform_L[231][2];				l_cell_reg[232] = inform_L[232][2];				l_cell_reg[233] = inform_L[234][2];				l_cell_reg[234] = inform_L[233][2];				l_cell_reg[235] = inform_L[235][2];				l_cell_reg[236] = inform_L[236][2];				l_cell_reg[237] = inform_L[238][2];				l_cell_reg[238] = inform_L[237][2];				l_cell_reg[239] = inform_L[239][2];				l_cell_reg[240] = inform_L[240][2];				l_cell_reg[241] = inform_L[242][2];				l_cell_reg[242] = inform_L[241][2];				l_cell_reg[243] = inform_L[243][2];				l_cell_reg[244] = inform_L[244][2];				l_cell_reg[245] = inform_L[246][2];				l_cell_reg[246] = inform_L[245][2];				l_cell_reg[247] = inform_L[247][2];				l_cell_reg[248] = inform_L[248][2];				l_cell_reg[249] = inform_L[250][2];				l_cell_reg[250] = inform_L[249][2];				l_cell_reg[251] = inform_L[251][2];				l_cell_reg[252] = inform_L[252][2];				l_cell_reg[253] = inform_L[254][2];				l_cell_reg[254] = inform_L[253][2];				l_cell_reg[255] = inform_L[255][2];				l_cell_reg[256] = inform_L[256][2];				l_cell_reg[257] = inform_L[258][2];				l_cell_reg[258] = inform_L[257][2];				l_cell_reg[259] = inform_L[259][2];				l_cell_reg[260] = inform_L[260][2];				l_cell_reg[261] = inform_L[262][2];				l_cell_reg[262] = inform_L[261][2];				l_cell_reg[263] = inform_L[263][2];				l_cell_reg[264] = inform_L[264][2];				l_cell_reg[265] = inform_L[266][2];				l_cell_reg[266] = inform_L[265][2];				l_cell_reg[267] = inform_L[267][2];				l_cell_reg[268] = inform_L[268][2];				l_cell_reg[269] = inform_L[270][2];				l_cell_reg[270] = inform_L[269][2];				l_cell_reg[271] = inform_L[271][2];				l_cell_reg[272] = inform_L[272][2];				l_cell_reg[273] = inform_L[274][2];				l_cell_reg[274] = inform_L[273][2];				l_cell_reg[275] = inform_L[275][2];				l_cell_reg[276] = inform_L[276][2];				l_cell_reg[277] = inform_L[278][2];				l_cell_reg[278] = inform_L[277][2];				l_cell_reg[279] = inform_L[279][2];				l_cell_reg[280] = inform_L[280][2];				l_cell_reg[281] = inform_L[282][2];				l_cell_reg[282] = inform_L[281][2];				l_cell_reg[283] = inform_L[283][2];				l_cell_reg[284] = inform_L[284][2];				l_cell_reg[285] = inform_L[286][2];				l_cell_reg[286] = inform_L[285][2];				l_cell_reg[287] = inform_L[287][2];				l_cell_reg[288] = inform_L[288][2];				l_cell_reg[289] = inform_L[290][2];				l_cell_reg[290] = inform_L[289][2];				l_cell_reg[291] = inform_L[291][2];				l_cell_reg[292] = inform_L[292][2];				l_cell_reg[293] = inform_L[294][2];				l_cell_reg[294] = inform_L[293][2];				l_cell_reg[295] = inform_L[295][2];				l_cell_reg[296] = inform_L[296][2];				l_cell_reg[297] = inform_L[298][2];				l_cell_reg[298] = inform_L[297][2];				l_cell_reg[299] = inform_L[299][2];				l_cell_reg[300] = inform_L[300][2];				l_cell_reg[301] = inform_L[302][2];				l_cell_reg[302] = inform_L[301][2];				l_cell_reg[303] = inform_L[303][2];				l_cell_reg[304] = inform_L[304][2];				l_cell_reg[305] = inform_L[306][2];				l_cell_reg[306] = inform_L[305][2];				l_cell_reg[307] = inform_L[307][2];				l_cell_reg[308] = inform_L[308][2];				l_cell_reg[309] = inform_L[310][2];				l_cell_reg[310] = inform_L[309][2];				l_cell_reg[311] = inform_L[311][2];				l_cell_reg[312] = inform_L[312][2];				l_cell_reg[313] = inform_L[314][2];				l_cell_reg[314] = inform_L[313][2];				l_cell_reg[315] = inform_L[315][2];				l_cell_reg[316] = inform_L[316][2];				l_cell_reg[317] = inform_L[318][2];				l_cell_reg[318] = inform_L[317][2];				l_cell_reg[319] = inform_L[319][2];				l_cell_reg[320] = inform_L[320][2];				l_cell_reg[321] = inform_L[322][2];				l_cell_reg[322] = inform_L[321][2];				l_cell_reg[323] = inform_L[323][2];				l_cell_reg[324] = inform_L[324][2];				l_cell_reg[325] = inform_L[326][2];				l_cell_reg[326] = inform_L[325][2];				l_cell_reg[327] = inform_L[327][2];				l_cell_reg[328] = inform_L[328][2];				l_cell_reg[329] = inform_L[330][2];				l_cell_reg[330] = inform_L[329][2];				l_cell_reg[331] = inform_L[331][2];				l_cell_reg[332] = inform_L[332][2];				l_cell_reg[333] = inform_L[334][2];				l_cell_reg[334] = inform_L[333][2];				l_cell_reg[335] = inform_L[335][2];				l_cell_reg[336] = inform_L[336][2];				l_cell_reg[337] = inform_L[338][2];				l_cell_reg[338] = inform_L[337][2];				l_cell_reg[339] = inform_L[339][2];				l_cell_reg[340] = inform_L[340][2];				l_cell_reg[341] = inform_L[342][2];				l_cell_reg[342] = inform_L[341][2];				l_cell_reg[343] = inform_L[343][2];				l_cell_reg[344] = inform_L[344][2];				l_cell_reg[345] = inform_L[346][2];				l_cell_reg[346] = inform_L[345][2];				l_cell_reg[347] = inform_L[347][2];				l_cell_reg[348] = inform_L[348][2];				l_cell_reg[349] = inform_L[350][2];				l_cell_reg[350] = inform_L[349][2];				l_cell_reg[351] = inform_L[351][2];				l_cell_reg[352] = inform_L[352][2];				l_cell_reg[353] = inform_L[354][2];				l_cell_reg[354] = inform_L[353][2];				l_cell_reg[355] = inform_L[355][2];				l_cell_reg[356] = inform_L[356][2];				l_cell_reg[357] = inform_L[358][2];				l_cell_reg[358] = inform_L[357][2];				l_cell_reg[359] = inform_L[359][2];				l_cell_reg[360] = inform_L[360][2];				l_cell_reg[361] = inform_L[362][2];				l_cell_reg[362] = inform_L[361][2];				l_cell_reg[363] = inform_L[363][2];				l_cell_reg[364] = inform_L[364][2];				l_cell_reg[365] = inform_L[366][2];				l_cell_reg[366] = inform_L[365][2];				l_cell_reg[367] = inform_L[367][2];				l_cell_reg[368] = inform_L[368][2];				l_cell_reg[369] = inform_L[370][2];				l_cell_reg[370] = inform_L[369][2];				l_cell_reg[371] = inform_L[371][2];				l_cell_reg[372] = inform_L[372][2];				l_cell_reg[373] = inform_L[374][2];				l_cell_reg[374] = inform_L[373][2];				l_cell_reg[375] = inform_L[375][2];				l_cell_reg[376] = inform_L[376][2];				l_cell_reg[377] = inform_L[378][2];				l_cell_reg[378] = inform_L[377][2];				l_cell_reg[379] = inform_L[379][2];				l_cell_reg[380] = inform_L[380][2];				l_cell_reg[381] = inform_L[382][2];				l_cell_reg[382] = inform_L[381][2];				l_cell_reg[383] = inform_L[383][2];				l_cell_reg[384] = inform_L[384][2];				l_cell_reg[385] = inform_L[386][2];				l_cell_reg[386] = inform_L[385][2];				l_cell_reg[387] = inform_L[387][2];				l_cell_reg[388] = inform_L[388][2];				l_cell_reg[389] = inform_L[390][2];				l_cell_reg[390] = inform_L[389][2];				l_cell_reg[391] = inform_L[391][2];				l_cell_reg[392] = inform_L[392][2];				l_cell_reg[393] = inform_L[394][2];				l_cell_reg[394] = inform_L[393][2];				l_cell_reg[395] = inform_L[395][2];				l_cell_reg[396] = inform_L[396][2];				l_cell_reg[397] = inform_L[398][2];				l_cell_reg[398] = inform_L[397][2];				l_cell_reg[399] = inform_L[399][2];				l_cell_reg[400] = inform_L[400][2];				l_cell_reg[401] = inform_L[402][2];				l_cell_reg[402] = inform_L[401][2];				l_cell_reg[403] = inform_L[403][2];				l_cell_reg[404] = inform_L[404][2];				l_cell_reg[405] = inform_L[406][2];				l_cell_reg[406] = inform_L[405][2];				l_cell_reg[407] = inform_L[407][2];				l_cell_reg[408] = inform_L[408][2];				l_cell_reg[409] = inform_L[410][2];				l_cell_reg[410] = inform_L[409][2];				l_cell_reg[411] = inform_L[411][2];				l_cell_reg[412] = inform_L[412][2];				l_cell_reg[413] = inform_L[414][2];				l_cell_reg[414] = inform_L[413][2];				l_cell_reg[415] = inform_L[415][2];				l_cell_reg[416] = inform_L[416][2];				l_cell_reg[417] = inform_L[418][2];				l_cell_reg[418] = inform_L[417][2];				l_cell_reg[419] = inform_L[419][2];				l_cell_reg[420] = inform_L[420][2];				l_cell_reg[421] = inform_L[422][2];				l_cell_reg[422] = inform_L[421][2];				l_cell_reg[423] = inform_L[423][2];				l_cell_reg[424] = inform_L[424][2];				l_cell_reg[425] = inform_L[426][2];				l_cell_reg[426] = inform_L[425][2];				l_cell_reg[427] = inform_L[427][2];				l_cell_reg[428] = inform_L[428][2];				l_cell_reg[429] = inform_L[430][2];				l_cell_reg[430] = inform_L[429][2];				l_cell_reg[431] = inform_L[431][2];				l_cell_reg[432] = inform_L[432][2];				l_cell_reg[433] = inform_L[434][2];				l_cell_reg[434] = inform_L[433][2];				l_cell_reg[435] = inform_L[435][2];				l_cell_reg[436] = inform_L[436][2];				l_cell_reg[437] = inform_L[438][2];				l_cell_reg[438] = inform_L[437][2];				l_cell_reg[439] = inform_L[439][2];				l_cell_reg[440] = inform_L[440][2];				l_cell_reg[441] = inform_L[442][2];				l_cell_reg[442] = inform_L[441][2];				l_cell_reg[443] = inform_L[443][2];				l_cell_reg[444] = inform_L[444][2];				l_cell_reg[445] = inform_L[446][2];				l_cell_reg[446] = inform_L[445][2];				l_cell_reg[447] = inform_L[447][2];				l_cell_reg[448] = inform_L[448][2];				l_cell_reg[449] = inform_L[450][2];				l_cell_reg[450] = inform_L[449][2];				l_cell_reg[451] = inform_L[451][2];				l_cell_reg[452] = inform_L[452][2];				l_cell_reg[453] = inform_L[454][2];				l_cell_reg[454] = inform_L[453][2];				l_cell_reg[455] = inform_L[455][2];				l_cell_reg[456] = inform_L[456][2];				l_cell_reg[457] = inform_L[458][2];				l_cell_reg[458] = inform_L[457][2];				l_cell_reg[459] = inform_L[459][2];				l_cell_reg[460] = inform_L[460][2];				l_cell_reg[461] = inform_L[462][2];				l_cell_reg[462] = inform_L[461][2];				l_cell_reg[463] = inform_L[463][2];				l_cell_reg[464] = inform_L[464][2];				l_cell_reg[465] = inform_L[466][2];				l_cell_reg[466] = inform_L[465][2];				l_cell_reg[467] = inform_L[467][2];				l_cell_reg[468] = inform_L[468][2];				l_cell_reg[469] = inform_L[470][2];				l_cell_reg[470] = inform_L[469][2];				l_cell_reg[471] = inform_L[471][2];				l_cell_reg[472] = inform_L[472][2];				l_cell_reg[473] = inform_L[474][2];				l_cell_reg[474] = inform_L[473][2];				l_cell_reg[475] = inform_L[475][2];				l_cell_reg[476] = inform_L[476][2];				l_cell_reg[477] = inform_L[478][2];				l_cell_reg[478] = inform_L[477][2];				l_cell_reg[479] = inform_L[479][2];				l_cell_reg[480] = inform_L[480][2];				l_cell_reg[481] = inform_L[482][2];				l_cell_reg[482] = inform_L[481][2];				l_cell_reg[483] = inform_L[483][2];				l_cell_reg[484] = inform_L[484][2];				l_cell_reg[485] = inform_L[486][2];				l_cell_reg[486] = inform_L[485][2];				l_cell_reg[487] = inform_L[487][2];				l_cell_reg[488] = inform_L[488][2];				l_cell_reg[489] = inform_L[490][2];				l_cell_reg[490] = inform_L[489][2];				l_cell_reg[491] = inform_L[491][2];				l_cell_reg[492] = inform_L[492][2];				l_cell_reg[493] = inform_L[494][2];				l_cell_reg[494] = inform_L[493][2];				l_cell_reg[495] = inform_L[495][2];				l_cell_reg[496] = inform_L[496][2];				l_cell_reg[497] = inform_L[498][2];				l_cell_reg[498] = inform_L[497][2];				l_cell_reg[499] = inform_L[499][2];				l_cell_reg[500] = inform_L[500][2];				l_cell_reg[501] = inform_L[502][2];				l_cell_reg[502] = inform_L[501][2];				l_cell_reg[503] = inform_L[503][2];				l_cell_reg[504] = inform_L[504][2];				l_cell_reg[505] = inform_L[506][2];				l_cell_reg[506] = inform_L[505][2];				l_cell_reg[507] = inform_L[507][2];				l_cell_reg[508] = inform_L[508][2];				l_cell_reg[509] = inform_L[510][2];				l_cell_reg[510] = inform_L[509][2];				l_cell_reg[511] = inform_L[511][2];				l_cell_reg[512] = inform_L[512][2];				l_cell_reg[513] = inform_L[514][2];				l_cell_reg[514] = inform_L[513][2];				l_cell_reg[515] = inform_L[515][2];				l_cell_reg[516] = inform_L[516][2];				l_cell_reg[517] = inform_L[518][2];				l_cell_reg[518] = inform_L[517][2];				l_cell_reg[519] = inform_L[519][2];				l_cell_reg[520] = inform_L[520][2];				l_cell_reg[521] = inform_L[522][2];				l_cell_reg[522] = inform_L[521][2];				l_cell_reg[523] = inform_L[523][2];				l_cell_reg[524] = inform_L[524][2];				l_cell_reg[525] = inform_L[526][2];				l_cell_reg[526] = inform_L[525][2];				l_cell_reg[527] = inform_L[527][2];				l_cell_reg[528] = inform_L[528][2];				l_cell_reg[529] = inform_L[530][2];				l_cell_reg[530] = inform_L[529][2];				l_cell_reg[531] = inform_L[531][2];				l_cell_reg[532] = inform_L[532][2];				l_cell_reg[533] = inform_L[534][2];				l_cell_reg[534] = inform_L[533][2];				l_cell_reg[535] = inform_L[535][2];				l_cell_reg[536] = inform_L[536][2];				l_cell_reg[537] = inform_L[538][2];				l_cell_reg[538] = inform_L[537][2];				l_cell_reg[539] = inform_L[539][2];				l_cell_reg[540] = inform_L[540][2];				l_cell_reg[541] = inform_L[542][2];				l_cell_reg[542] = inform_L[541][2];				l_cell_reg[543] = inform_L[543][2];				l_cell_reg[544] = inform_L[544][2];				l_cell_reg[545] = inform_L[546][2];				l_cell_reg[546] = inform_L[545][2];				l_cell_reg[547] = inform_L[547][2];				l_cell_reg[548] = inform_L[548][2];				l_cell_reg[549] = inform_L[550][2];				l_cell_reg[550] = inform_L[549][2];				l_cell_reg[551] = inform_L[551][2];				l_cell_reg[552] = inform_L[552][2];				l_cell_reg[553] = inform_L[554][2];				l_cell_reg[554] = inform_L[553][2];				l_cell_reg[555] = inform_L[555][2];				l_cell_reg[556] = inform_L[556][2];				l_cell_reg[557] = inform_L[558][2];				l_cell_reg[558] = inform_L[557][2];				l_cell_reg[559] = inform_L[559][2];				l_cell_reg[560] = inform_L[560][2];				l_cell_reg[561] = inform_L[562][2];				l_cell_reg[562] = inform_L[561][2];				l_cell_reg[563] = inform_L[563][2];				l_cell_reg[564] = inform_L[564][2];				l_cell_reg[565] = inform_L[566][2];				l_cell_reg[566] = inform_L[565][2];				l_cell_reg[567] = inform_L[567][2];				l_cell_reg[568] = inform_L[568][2];				l_cell_reg[569] = inform_L[570][2];				l_cell_reg[570] = inform_L[569][2];				l_cell_reg[571] = inform_L[571][2];				l_cell_reg[572] = inform_L[572][2];				l_cell_reg[573] = inform_L[574][2];				l_cell_reg[574] = inform_L[573][2];				l_cell_reg[575] = inform_L[575][2];				l_cell_reg[576] = inform_L[576][2];				l_cell_reg[577] = inform_L[578][2];				l_cell_reg[578] = inform_L[577][2];				l_cell_reg[579] = inform_L[579][2];				l_cell_reg[580] = inform_L[580][2];				l_cell_reg[581] = inform_L[582][2];				l_cell_reg[582] = inform_L[581][2];				l_cell_reg[583] = inform_L[583][2];				l_cell_reg[584] = inform_L[584][2];				l_cell_reg[585] = inform_L[586][2];				l_cell_reg[586] = inform_L[585][2];				l_cell_reg[587] = inform_L[587][2];				l_cell_reg[588] = inform_L[588][2];				l_cell_reg[589] = inform_L[590][2];				l_cell_reg[590] = inform_L[589][2];				l_cell_reg[591] = inform_L[591][2];				l_cell_reg[592] = inform_L[592][2];				l_cell_reg[593] = inform_L[594][2];				l_cell_reg[594] = inform_L[593][2];				l_cell_reg[595] = inform_L[595][2];				l_cell_reg[596] = inform_L[596][2];				l_cell_reg[597] = inform_L[598][2];				l_cell_reg[598] = inform_L[597][2];				l_cell_reg[599] = inform_L[599][2];				l_cell_reg[600] = inform_L[600][2];				l_cell_reg[601] = inform_L[602][2];				l_cell_reg[602] = inform_L[601][2];				l_cell_reg[603] = inform_L[603][2];				l_cell_reg[604] = inform_L[604][2];				l_cell_reg[605] = inform_L[606][2];				l_cell_reg[606] = inform_L[605][2];				l_cell_reg[607] = inform_L[607][2];				l_cell_reg[608] = inform_L[608][2];				l_cell_reg[609] = inform_L[610][2];				l_cell_reg[610] = inform_L[609][2];				l_cell_reg[611] = inform_L[611][2];				l_cell_reg[612] = inform_L[612][2];				l_cell_reg[613] = inform_L[614][2];				l_cell_reg[614] = inform_L[613][2];				l_cell_reg[615] = inform_L[615][2];				l_cell_reg[616] = inform_L[616][2];				l_cell_reg[617] = inform_L[618][2];				l_cell_reg[618] = inform_L[617][2];				l_cell_reg[619] = inform_L[619][2];				l_cell_reg[620] = inform_L[620][2];				l_cell_reg[621] = inform_L[622][2];				l_cell_reg[622] = inform_L[621][2];				l_cell_reg[623] = inform_L[623][2];				l_cell_reg[624] = inform_L[624][2];				l_cell_reg[625] = inform_L[626][2];				l_cell_reg[626] = inform_L[625][2];				l_cell_reg[627] = inform_L[627][2];				l_cell_reg[628] = inform_L[628][2];				l_cell_reg[629] = inform_L[630][2];				l_cell_reg[630] = inform_L[629][2];				l_cell_reg[631] = inform_L[631][2];				l_cell_reg[632] = inform_L[632][2];				l_cell_reg[633] = inform_L[634][2];				l_cell_reg[634] = inform_L[633][2];				l_cell_reg[635] = inform_L[635][2];				l_cell_reg[636] = inform_L[636][2];				l_cell_reg[637] = inform_L[638][2];				l_cell_reg[638] = inform_L[637][2];				l_cell_reg[639] = inform_L[639][2];				l_cell_reg[640] = inform_L[640][2];				l_cell_reg[641] = inform_L[642][2];				l_cell_reg[642] = inform_L[641][2];				l_cell_reg[643] = inform_L[643][2];				l_cell_reg[644] = inform_L[644][2];				l_cell_reg[645] = inform_L[646][2];				l_cell_reg[646] = inform_L[645][2];				l_cell_reg[647] = inform_L[647][2];				l_cell_reg[648] = inform_L[648][2];				l_cell_reg[649] = inform_L[650][2];				l_cell_reg[650] = inform_L[649][2];				l_cell_reg[651] = inform_L[651][2];				l_cell_reg[652] = inform_L[652][2];				l_cell_reg[653] = inform_L[654][2];				l_cell_reg[654] = inform_L[653][2];				l_cell_reg[655] = inform_L[655][2];				l_cell_reg[656] = inform_L[656][2];				l_cell_reg[657] = inform_L[658][2];				l_cell_reg[658] = inform_L[657][2];				l_cell_reg[659] = inform_L[659][2];				l_cell_reg[660] = inform_L[660][2];				l_cell_reg[661] = inform_L[662][2];				l_cell_reg[662] = inform_L[661][2];				l_cell_reg[663] = inform_L[663][2];				l_cell_reg[664] = inform_L[664][2];				l_cell_reg[665] = inform_L[666][2];				l_cell_reg[666] = inform_L[665][2];				l_cell_reg[667] = inform_L[667][2];				l_cell_reg[668] = inform_L[668][2];				l_cell_reg[669] = inform_L[670][2];				l_cell_reg[670] = inform_L[669][2];				l_cell_reg[671] = inform_L[671][2];				l_cell_reg[672] = inform_L[672][2];				l_cell_reg[673] = inform_L[674][2];				l_cell_reg[674] = inform_L[673][2];				l_cell_reg[675] = inform_L[675][2];				l_cell_reg[676] = inform_L[676][2];				l_cell_reg[677] = inform_L[678][2];				l_cell_reg[678] = inform_L[677][2];				l_cell_reg[679] = inform_L[679][2];				l_cell_reg[680] = inform_L[680][2];				l_cell_reg[681] = inform_L[682][2];				l_cell_reg[682] = inform_L[681][2];				l_cell_reg[683] = inform_L[683][2];				l_cell_reg[684] = inform_L[684][2];				l_cell_reg[685] = inform_L[686][2];				l_cell_reg[686] = inform_L[685][2];				l_cell_reg[687] = inform_L[687][2];				l_cell_reg[688] = inform_L[688][2];				l_cell_reg[689] = inform_L[690][2];				l_cell_reg[690] = inform_L[689][2];				l_cell_reg[691] = inform_L[691][2];				l_cell_reg[692] = inform_L[692][2];				l_cell_reg[693] = inform_L[694][2];				l_cell_reg[694] = inform_L[693][2];				l_cell_reg[695] = inform_L[695][2];				l_cell_reg[696] = inform_L[696][2];				l_cell_reg[697] = inform_L[698][2];				l_cell_reg[698] = inform_L[697][2];				l_cell_reg[699] = inform_L[699][2];				l_cell_reg[700] = inform_L[700][2];				l_cell_reg[701] = inform_L[702][2];				l_cell_reg[702] = inform_L[701][2];				l_cell_reg[703] = inform_L[703][2];				l_cell_reg[704] = inform_L[704][2];				l_cell_reg[705] = inform_L[706][2];				l_cell_reg[706] = inform_L[705][2];				l_cell_reg[707] = inform_L[707][2];				l_cell_reg[708] = inform_L[708][2];				l_cell_reg[709] = inform_L[710][2];				l_cell_reg[710] = inform_L[709][2];				l_cell_reg[711] = inform_L[711][2];				l_cell_reg[712] = inform_L[712][2];				l_cell_reg[713] = inform_L[714][2];				l_cell_reg[714] = inform_L[713][2];				l_cell_reg[715] = inform_L[715][2];				l_cell_reg[716] = inform_L[716][2];				l_cell_reg[717] = inform_L[718][2];				l_cell_reg[718] = inform_L[717][2];				l_cell_reg[719] = inform_L[719][2];				l_cell_reg[720] = inform_L[720][2];				l_cell_reg[721] = inform_L[722][2];				l_cell_reg[722] = inform_L[721][2];				l_cell_reg[723] = inform_L[723][2];				l_cell_reg[724] = inform_L[724][2];				l_cell_reg[725] = inform_L[726][2];				l_cell_reg[726] = inform_L[725][2];				l_cell_reg[727] = inform_L[727][2];				l_cell_reg[728] = inform_L[728][2];				l_cell_reg[729] = inform_L[730][2];				l_cell_reg[730] = inform_L[729][2];				l_cell_reg[731] = inform_L[731][2];				l_cell_reg[732] = inform_L[732][2];				l_cell_reg[733] = inform_L[734][2];				l_cell_reg[734] = inform_L[733][2];				l_cell_reg[735] = inform_L[735][2];				l_cell_reg[736] = inform_L[736][2];				l_cell_reg[737] = inform_L[738][2];				l_cell_reg[738] = inform_L[737][2];				l_cell_reg[739] = inform_L[739][2];				l_cell_reg[740] = inform_L[740][2];				l_cell_reg[741] = inform_L[742][2];				l_cell_reg[742] = inform_L[741][2];				l_cell_reg[743] = inform_L[743][2];				l_cell_reg[744] = inform_L[744][2];				l_cell_reg[745] = inform_L[746][2];				l_cell_reg[746] = inform_L[745][2];				l_cell_reg[747] = inform_L[747][2];				l_cell_reg[748] = inform_L[748][2];				l_cell_reg[749] = inform_L[750][2];				l_cell_reg[750] = inform_L[749][2];				l_cell_reg[751] = inform_L[751][2];				l_cell_reg[752] = inform_L[752][2];				l_cell_reg[753] = inform_L[754][2];				l_cell_reg[754] = inform_L[753][2];				l_cell_reg[755] = inform_L[755][2];				l_cell_reg[756] = inform_L[756][2];				l_cell_reg[757] = inform_L[758][2];				l_cell_reg[758] = inform_L[757][2];				l_cell_reg[759] = inform_L[759][2];				l_cell_reg[760] = inform_L[760][2];				l_cell_reg[761] = inform_L[762][2];				l_cell_reg[762] = inform_L[761][2];				l_cell_reg[763] = inform_L[763][2];				l_cell_reg[764] = inform_L[764][2];				l_cell_reg[765] = inform_L[766][2];				l_cell_reg[766] = inform_L[765][2];				l_cell_reg[767] = inform_L[767][2];				l_cell_reg[768] = inform_L[768][2];				l_cell_reg[769] = inform_L[770][2];				l_cell_reg[770] = inform_L[769][2];				l_cell_reg[771] = inform_L[771][2];				l_cell_reg[772] = inform_L[772][2];				l_cell_reg[773] = inform_L[774][2];				l_cell_reg[774] = inform_L[773][2];				l_cell_reg[775] = inform_L[775][2];				l_cell_reg[776] = inform_L[776][2];				l_cell_reg[777] = inform_L[778][2];				l_cell_reg[778] = inform_L[777][2];				l_cell_reg[779] = inform_L[779][2];				l_cell_reg[780] = inform_L[780][2];				l_cell_reg[781] = inform_L[782][2];				l_cell_reg[782] = inform_L[781][2];				l_cell_reg[783] = inform_L[783][2];				l_cell_reg[784] = inform_L[784][2];				l_cell_reg[785] = inform_L[786][2];				l_cell_reg[786] = inform_L[785][2];				l_cell_reg[787] = inform_L[787][2];				l_cell_reg[788] = inform_L[788][2];				l_cell_reg[789] = inform_L[790][2];				l_cell_reg[790] = inform_L[789][2];				l_cell_reg[791] = inform_L[791][2];				l_cell_reg[792] = inform_L[792][2];				l_cell_reg[793] = inform_L[794][2];				l_cell_reg[794] = inform_L[793][2];				l_cell_reg[795] = inform_L[795][2];				l_cell_reg[796] = inform_L[796][2];				l_cell_reg[797] = inform_L[798][2];				l_cell_reg[798] = inform_L[797][2];				l_cell_reg[799] = inform_L[799][2];				l_cell_reg[800] = inform_L[800][2];				l_cell_reg[801] = inform_L[802][2];				l_cell_reg[802] = inform_L[801][2];				l_cell_reg[803] = inform_L[803][2];				l_cell_reg[804] = inform_L[804][2];				l_cell_reg[805] = inform_L[806][2];				l_cell_reg[806] = inform_L[805][2];				l_cell_reg[807] = inform_L[807][2];				l_cell_reg[808] = inform_L[808][2];				l_cell_reg[809] = inform_L[810][2];				l_cell_reg[810] = inform_L[809][2];				l_cell_reg[811] = inform_L[811][2];				l_cell_reg[812] = inform_L[812][2];				l_cell_reg[813] = inform_L[814][2];				l_cell_reg[814] = inform_L[813][2];				l_cell_reg[815] = inform_L[815][2];				l_cell_reg[816] = inform_L[816][2];				l_cell_reg[817] = inform_L[818][2];				l_cell_reg[818] = inform_L[817][2];				l_cell_reg[819] = inform_L[819][2];				l_cell_reg[820] = inform_L[820][2];				l_cell_reg[821] = inform_L[822][2];				l_cell_reg[822] = inform_L[821][2];				l_cell_reg[823] = inform_L[823][2];				l_cell_reg[824] = inform_L[824][2];				l_cell_reg[825] = inform_L[826][2];				l_cell_reg[826] = inform_L[825][2];				l_cell_reg[827] = inform_L[827][2];				l_cell_reg[828] = inform_L[828][2];				l_cell_reg[829] = inform_L[830][2];				l_cell_reg[830] = inform_L[829][2];				l_cell_reg[831] = inform_L[831][2];				l_cell_reg[832] = inform_L[832][2];				l_cell_reg[833] = inform_L[834][2];				l_cell_reg[834] = inform_L[833][2];				l_cell_reg[835] = inform_L[835][2];				l_cell_reg[836] = inform_L[836][2];				l_cell_reg[837] = inform_L[838][2];				l_cell_reg[838] = inform_L[837][2];				l_cell_reg[839] = inform_L[839][2];				l_cell_reg[840] = inform_L[840][2];				l_cell_reg[841] = inform_L[842][2];				l_cell_reg[842] = inform_L[841][2];				l_cell_reg[843] = inform_L[843][2];				l_cell_reg[844] = inform_L[844][2];				l_cell_reg[845] = inform_L[846][2];				l_cell_reg[846] = inform_L[845][2];				l_cell_reg[847] = inform_L[847][2];				l_cell_reg[848] = inform_L[848][2];				l_cell_reg[849] = inform_L[850][2];				l_cell_reg[850] = inform_L[849][2];				l_cell_reg[851] = inform_L[851][2];				l_cell_reg[852] = inform_L[852][2];				l_cell_reg[853] = inform_L[854][2];				l_cell_reg[854] = inform_L[853][2];				l_cell_reg[855] = inform_L[855][2];				l_cell_reg[856] = inform_L[856][2];				l_cell_reg[857] = inform_L[858][2];				l_cell_reg[858] = inform_L[857][2];				l_cell_reg[859] = inform_L[859][2];				l_cell_reg[860] = inform_L[860][2];				l_cell_reg[861] = inform_L[862][2];				l_cell_reg[862] = inform_L[861][2];				l_cell_reg[863] = inform_L[863][2];				l_cell_reg[864] = inform_L[864][2];				l_cell_reg[865] = inform_L[866][2];				l_cell_reg[866] = inform_L[865][2];				l_cell_reg[867] = inform_L[867][2];				l_cell_reg[868] = inform_L[868][2];				l_cell_reg[869] = inform_L[870][2];				l_cell_reg[870] = inform_L[869][2];				l_cell_reg[871] = inform_L[871][2];				l_cell_reg[872] = inform_L[872][2];				l_cell_reg[873] = inform_L[874][2];				l_cell_reg[874] = inform_L[873][2];				l_cell_reg[875] = inform_L[875][2];				l_cell_reg[876] = inform_L[876][2];				l_cell_reg[877] = inform_L[878][2];				l_cell_reg[878] = inform_L[877][2];				l_cell_reg[879] = inform_L[879][2];				l_cell_reg[880] = inform_L[880][2];				l_cell_reg[881] = inform_L[882][2];				l_cell_reg[882] = inform_L[881][2];				l_cell_reg[883] = inform_L[883][2];				l_cell_reg[884] = inform_L[884][2];				l_cell_reg[885] = inform_L[886][2];				l_cell_reg[886] = inform_L[885][2];				l_cell_reg[887] = inform_L[887][2];				l_cell_reg[888] = inform_L[888][2];				l_cell_reg[889] = inform_L[890][2];				l_cell_reg[890] = inform_L[889][2];				l_cell_reg[891] = inform_L[891][2];				l_cell_reg[892] = inform_L[892][2];				l_cell_reg[893] = inform_L[894][2];				l_cell_reg[894] = inform_L[893][2];				l_cell_reg[895] = inform_L[895][2];				l_cell_reg[896] = inform_L[896][2];				l_cell_reg[897] = inform_L[898][2];				l_cell_reg[898] = inform_L[897][2];				l_cell_reg[899] = inform_L[899][2];				l_cell_reg[900] = inform_L[900][2];				l_cell_reg[901] = inform_L[902][2];				l_cell_reg[902] = inform_L[901][2];				l_cell_reg[903] = inform_L[903][2];				l_cell_reg[904] = inform_L[904][2];				l_cell_reg[905] = inform_L[906][2];				l_cell_reg[906] = inform_L[905][2];				l_cell_reg[907] = inform_L[907][2];				l_cell_reg[908] = inform_L[908][2];				l_cell_reg[909] = inform_L[910][2];				l_cell_reg[910] = inform_L[909][2];				l_cell_reg[911] = inform_L[911][2];				l_cell_reg[912] = inform_L[912][2];				l_cell_reg[913] = inform_L[914][2];				l_cell_reg[914] = inform_L[913][2];				l_cell_reg[915] = inform_L[915][2];				l_cell_reg[916] = inform_L[916][2];				l_cell_reg[917] = inform_L[918][2];				l_cell_reg[918] = inform_L[917][2];				l_cell_reg[919] = inform_L[919][2];				l_cell_reg[920] = inform_L[920][2];				l_cell_reg[921] = inform_L[922][2];				l_cell_reg[922] = inform_L[921][2];				l_cell_reg[923] = inform_L[923][2];				l_cell_reg[924] = inform_L[924][2];				l_cell_reg[925] = inform_L[926][2];				l_cell_reg[926] = inform_L[925][2];				l_cell_reg[927] = inform_L[927][2];				l_cell_reg[928] = inform_L[928][2];				l_cell_reg[929] = inform_L[930][2];				l_cell_reg[930] = inform_L[929][2];				l_cell_reg[931] = inform_L[931][2];				l_cell_reg[932] = inform_L[932][2];				l_cell_reg[933] = inform_L[934][2];				l_cell_reg[934] = inform_L[933][2];				l_cell_reg[935] = inform_L[935][2];				l_cell_reg[936] = inform_L[936][2];				l_cell_reg[937] = inform_L[938][2];				l_cell_reg[938] = inform_L[937][2];				l_cell_reg[939] = inform_L[939][2];				l_cell_reg[940] = inform_L[940][2];				l_cell_reg[941] = inform_L[942][2];				l_cell_reg[942] = inform_L[941][2];				l_cell_reg[943] = inform_L[943][2];				l_cell_reg[944] = inform_L[944][2];				l_cell_reg[945] = inform_L[946][2];				l_cell_reg[946] = inform_L[945][2];				l_cell_reg[947] = inform_L[947][2];				l_cell_reg[948] = inform_L[948][2];				l_cell_reg[949] = inform_L[950][2];				l_cell_reg[950] = inform_L[949][2];				l_cell_reg[951] = inform_L[951][2];				l_cell_reg[952] = inform_L[952][2];				l_cell_reg[953] = inform_L[954][2];				l_cell_reg[954] = inform_L[953][2];				l_cell_reg[955] = inform_L[955][2];				l_cell_reg[956] = inform_L[956][2];				l_cell_reg[957] = inform_L[958][2];				l_cell_reg[958] = inform_L[957][2];				l_cell_reg[959] = inform_L[959][2];				l_cell_reg[960] = inform_L[960][2];				l_cell_reg[961] = inform_L[962][2];				l_cell_reg[962] = inform_L[961][2];				l_cell_reg[963] = inform_L[963][2];				l_cell_reg[964] = inform_L[964][2];				l_cell_reg[965] = inform_L[966][2];				l_cell_reg[966] = inform_L[965][2];				l_cell_reg[967] = inform_L[967][2];				l_cell_reg[968] = inform_L[968][2];				l_cell_reg[969] = inform_L[970][2];				l_cell_reg[970] = inform_L[969][2];				l_cell_reg[971] = inform_L[971][2];				l_cell_reg[972] = inform_L[972][2];				l_cell_reg[973] = inform_L[974][2];				l_cell_reg[974] = inform_L[973][2];				l_cell_reg[975] = inform_L[975][2];				l_cell_reg[976] = inform_L[976][2];				l_cell_reg[977] = inform_L[978][2];				l_cell_reg[978] = inform_L[977][2];				l_cell_reg[979] = inform_L[979][2];				l_cell_reg[980] = inform_L[980][2];				l_cell_reg[981] = inform_L[982][2];				l_cell_reg[982] = inform_L[981][2];				l_cell_reg[983] = inform_L[983][2];				l_cell_reg[984] = inform_L[984][2];				l_cell_reg[985] = inform_L[986][2];				l_cell_reg[986] = inform_L[985][2];				l_cell_reg[987] = inform_L[987][2];				l_cell_reg[988] = inform_L[988][2];				l_cell_reg[989] = inform_L[990][2];				l_cell_reg[990] = inform_L[989][2];				l_cell_reg[991] = inform_L[991][2];				l_cell_reg[992] = inform_L[992][2];				l_cell_reg[993] = inform_L[994][2];				l_cell_reg[994] = inform_L[993][2];				l_cell_reg[995] = inform_L[995][2];				l_cell_reg[996] = inform_L[996][2];				l_cell_reg[997] = inform_L[998][2];				l_cell_reg[998] = inform_L[997][2];				l_cell_reg[999] = inform_L[999][2];				l_cell_reg[1000] = inform_L[1000][2];				l_cell_reg[1001] = inform_L[1002][2];				l_cell_reg[1002] = inform_L[1001][2];				l_cell_reg[1003] = inform_L[1003][2];				l_cell_reg[1004] = inform_L[1004][2];				l_cell_reg[1005] = inform_L[1006][2];				l_cell_reg[1006] = inform_L[1005][2];				l_cell_reg[1007] = inform_L[1007][2];				l_cell_reg[1008] = inform_L[1008][2];				l_cell_reg[1009] = inform_L[1010][2];				l_cell_reg[1010] = inform_L[1009][2];				l_cell_reg[1011] = inform_L[1011][2];				l_cell_reg[1012] = inform_L[1012][2];				l_cell_reg[1013] = inform_L[1014][2];				l_cell_reg[1014] = inform_L[1013][2];				l_cell_reg[1015] = inform_L[1015][2];				l_cell_reg[1016] = inform_L[1016][2];				l_cell_reg[1017] = inform_L[1018][2];				l_cell_reg[1018] = inform_L[1017][2];				l_cell_reg[1019] = inform_L[1019][2];				l_cell_reg[1020] = inform_L[1020][2];				l_cell_reg[1021] = inform_L[1022][2];				l_cell_reg[1022] = inform_L[1021][2];				l_cell_reg[1023] = inform_L[1023][2];			end
			3:			begin				r_cell_reg[0] = inform_R[0][2];				r_cell_reg[1] = inform_R[4][2];				r_cell_reg[2] = inform_R[1][2];				r_cell_reg[3] = inform_R[5][2];				r_cell_reg[4] = inform_R[2][2];				r_cell_reg[5] = inform_R[6][2];				r_cell_reg[6] = inform_R[3][2];				r_cell_reg[7] = inform_R[7][2];				r_cell_reg[8] = inform_R[8][2];				r_cell_reg[9] = inform_R[12][2];				r_cell_reg[10] = inform_R[9][2];				r_cell_reg[11] = inform_R[13][2];				r_cell_reg[12] = inform_R[10][2];				r_cell_reg[13] = inform_R[14][2];				r_cell_reg[14] = inform_R[11][2];				r_cell_reg[15] = inform_R[15][2];				r_cell_reg[16] = inform_R[16][2];				r_cell_reg[17] = inform_R[20][2];				r_cell_reg[18] = inform_R[17][2];				r_cell_reg[19] = inform_R[21][2];				r_cell_reg[20] = inform_R[18][2];				r_cell_reg[21] = inform_R[22][2];				r_cell_reg[22] = inform_R[19][2];				r_cell_reg[23] = inform_R[23][2];				r_cell_reg[24] = inform_R[24][2];				r_cell_reg[25] = inform_R[28][2];				r_cell_reg[26] = inform_R[25][2];				r_cell_reg[27] = inform_R[29][2];				r_cell_reg[28] = inform_R[26][2];				r_cell_reg[29] = inform_R[30][2];				r_cell_reg[30] = inform_R[27][2];				r_cell_reg[31] = inform_R[31][2];				r_cell_reg[32] = inform_R[32][2];				r_cell_reg[33] = inform_R[36][2];				r_cell_reg[34] = inform_R[33][2];				r_cell_reg[35] = inform_R[37][2];				r_cell_reg[36] = inform_R[34][2];				r_cell_reg[37] = inform_R[38][2];				r_cell_reg[38] = inform_R[35][2];				r_cell_reg[39] = inform_R[39][2];				r_cell_reg[40] = inform_R[40][2];				r_cell_reg[41] = inform_R[44][2];				r_cell_reg[42] = inform_R[41][2];				r_cell_reg[43] = inform_R[45][2];				r_cell_reg[44] = inform_R[42][2];				r_cell_reg[45] = inform_R[46][2];				r_cell_reg[46] = inform_R[43][2];				r_cell_reg[47] = inform_R[47][2];				r_cell_reg[48] = inform_R[48][2];				r_cell_reg[49] = inform_R[52][2];				r_cell_reg[50] = inform_R[49][2];				r_cell_reg[51] = inform_R[53][2];				r_cell_reg[52] = inform_R[50][2];				r_cell_reg[53] = inform_R[54][2];				r_cell_reg[54] = inform_R[51][2];				r_cell_reg[55] = inform_R[55][2];				r_cell_reg[56] = inform_R[56][2];				r_cell_reg[57] = inform_R[60][2];				r_cell_reg[58] = inform_R[57][2];				r_cell_reg[59] = inform_R[61][2];				r_cell_reg[60] = inform_R[58][2];				r_cell_reg[61] = inform_R[62][2];				r_cell_reg[62] = inform_R[59][2];				r_cell_reg[63] = inform_R[63][2];				r_cell_reg[64] = inform_R[64][2];				r_cell_reg[65] = inform_R[68][2];				r_cell_reg[66] = inform_R[65][2];				r_cell_reg[67] = inform_R[69][2];				r_cell_reg[68] = inform_R[66][2];				r_cell_reg[69] = inform_R[70][2];				r_cell_reg[70] = inform_R[67][2];				r_cell_reg[71] = inform_R[71][2];				r_cell_reg[72] = inform_R[72][2];				r_cell_reg[73] = inform_R[76][2];				r_cell_reg[74] = inform_R[73][2];				r_cell_reg[75] = inform_R[77][2];				r_cell_reg[76] = inform_R[74][2];				r_cell_reg[77] = inform_R[78][2];				r_cell_reg[78] = inform_R[75][2];				r_cell_reg[79] = inform_R[79][2];				r_cell_reg[80] = inform_R[80][2];				r_cell_reg[81] = inform_R[84][2];				r_cell_reg[82] = inform_R[81][2];				r_cell_reg[83] = inform_R[85][2];				r_cell_reg[84] = inform_R[82][2];				r_cell_reg[85] = inform_R[86][2];				r_cell_reg[86] = inform_R[83][2];				r_cell_reg[87] = inform_R[87][2];				r_cell_reg[88] = inform_R[88][2];				r_cell_reg[89] = inform_R[92][2];				r_cell_reg[90] = inform_R[89][2];				r_cell_reg[91] = inform_R[93][2];				r_cell_reg[92] = inform_R[90][2];				r_cell_reg[93] = inform_R[94][2];				r_cell_reg[94] = inform_R[91][2];				r_cell_reg[95] = inform_R[95][2];				r_cell_reg[96] = inform_R[96][2];				r_cell_reg[97] = inform_R[100][2];				r_cell_reg[98] = inform_R[97][2];				r_cell_reg[99] = inform_R[101][2];				r_cell_reg[100] = inform_R[98][2];				r_cell_reg[101] = inform_R[102][2];				r_cell_reg[102] = inform_R[99][2];				r_cell_reg[103] = inform_R[103][2];				r_cell_reg[104] = inform_R[104][2];				r_cell_reg[105] = inform_R[108][2];				r_cell_reg[106] = inform_R[105][2];				r_cell_reg[107] = inform_R[109][2];				r_cell_reg[108] = inform_R[106][2];				r_cell_reg[109] = inform_R[110][2];				r_cell_reg[110] = inform_R[107][2];				r_cell_reg[111] = inform_R[111][2];				r_cell_reg[112] = inform_R[112][2];				r_cell_reg[113] = inform_R[116][2];				r_cell_reg[114] = inform_R[113][2];				r_cell_reg[115] = inform_R[117][2];				r_cell_reg[116] = inform_R[114][2];				r_cell_reg[117] = inform_R[118][2];				r_cell_reg[118] = inform_R[115][2];				r_cell_reg[119] = inform_R[119][2];				r_cell_reg[120] = inform_R[120][2];				r_cell_reg[121] = inform_R[124][2];				r_cell_reg[122] = inform_R[121][2];				r_cell_reg[123] = inform_R[125][2];				r_cell_reg[124] = inform_R[122][2];				r_cell_reg[125] = inform_R[126][2];				r_cell_reg[126] = inform_R[123][2];				r_cell_reg[127] = inform_R[127][2];				r_cell_reg[128] = inform_R[128][2];				r_cell_reg[129] = inform_R[132][2];				r_cell_reg[130] = inform_R[129][2];				r_cell_reg[131] = inform_R[133][2];				r_cell_reg[132] = inform_R[130][2];				r_cell_reg[133] = inform_R[134][2];				r_cell_reg[134] = inform_R[131][2];				r_cell_reg[135] = inform_R[135][2];				r_cell_reg[136] = inform_R[136][2];				r_cell_reg[137] = inform_R[140][2];				r_cell_reg[138] = inform_R[137][2];				r_cell_reg[139] = inform_R[141][2];				r_cell_reg[140] = inform_R[138][2];				r_cell_reg[141] = inform_R[142][2];				r_cell_reg[142] = inform_R[139][2];				r_cell_reg[143] = inform_R[143][2];				r_cell_reg[144] = inform_R[144][2];				r_cell_reg[145] = inform_R[148][2];				r_cell_reg[146] = inform_R[145][2];				r_cell_reg[147] = inform_R[149][2];				r_cell_reg[148] = inform_R[146][2];				r_cell_reg[149] = inform_R[150][2];				r_cell_reg[150] = inform_R[147][2];				r_cell_reg[151] = inform_R[151][2];				r_cell_reg[152] = inform_R[152][2];				r_cell_reg[153] = inform_R[156][2];				r_cell_reg[154] = inform_R[153][2];				r_cell_reg[155] = inform_R[157][2];				r_cell_reg[156] = inform_R[154][2];				r_cell_reg[157] = inform_R[158][2];				r_cell_reg[158] = inform_R[155][2];				r_cell_reg[159] = inform_R[159][2];				r_cell_reg[160] = inform_R[160][2];				r_cell_reg[161] = inform_R[164][2];				r_cell_reg[162] = inform_R[161][2];				r_cell_reg[163] = inform_R[165][2];				r_cell_reg[164] = inform_R[162][2];				r_cell_reg[165] = inform_R[166][2];				r_cell_reg[166] = inform_R[163][2];				r_cell_reg[167] = inform_R[167][2];				r_cell_reg[168] = inform_R[168][2];				r_cell_reg[169] = inform_R[172][2];				r_cell_reg[170] = inform_R[169][2];				r_cell_reg[171] = inform_R[173][2];				r_cell_reg[172] = inform_R[170][2];				r_cell_reg[173] = inform_R[174][2];				r_cell_reg[174] = inform_R[171][2];				r_cell_reg[175] = inform_R[175][2];				r_cell_reg[176] = inform_R[176][2];				r_cell_reg[177] = inform_R[180][2];				r_cell_reg[178] = inform_R[177][2];				r_cell_reg[179] = inform_R[181][2];				r_cell_reg[180] = inform_R[178][2];				r_cell_reg[181] = inform_R[182][2];				r_cell_reg[182] = inform_R[179][2];				r_cell_reg[183] = inform_R[183][2];				r_cell_reg[184] = inform_R[184][2];				r_cell_reg[185] = inform_R[188][2];				r_cell_reg[186] = inform_R[185][2];				r_cell_reg[187] = inform_R[189][2];				r_cell_reg[188] = inform_R[186][2];				r_cell_reg[189] = inform_R[190][2];				r_cell_reg[190] = inform_R[187][2];				r_cell_reg[191] = inform_R[191][2];				r_cell_reg[192] = inform_R[192][2];				r_cell_reg[193] = inform_R[196][2];				r_cell_reg[194] = inform_R[193][2];				r_cell_reg[195] = inform_R[197][2];				r_cell_reg[196] = inform_R[194][2];				r_cell_reg[197] = inform_R[198][2];				r_cell_reg[198] = inform_R[195][2];				r_cell_reg[199] = inform_R[199][2];				r_cell_reg[200] = inform_R[200][2];				r_cell_reg[201] = inform_R[204][2];				r_cell_reg[202] = inform_R[201][2];				r_cell_reg[203] = inform_R[205][2];				r_cell_reg[204] = inform_R[202][2];				r_cell_reg[205] = inform_R[206][2];				r_cell_reg[206] = inform_R[203][2];				r_cell_reg[207] = inform_R[207][2];				r_cell_reg[208] = inform_R[208][2];				r_cell_reg[209] = inform_R[212][2];				r_cell_reg[210] = inform_R[209][2];				r_cell_reg[211] = inform_R[213][2];				r_cell_reg[212] = inform_R[210][2];				r_cell_reg[213] = inform_R[214][2];				r_cell_reg[214] = inform_R[211][2];				r_cell_reg[215] = inform_R[215][2];				r_cell_reg[216] = inform_R[216][2];				r_cell_reg[217] = inform_R[220][2];				r_cell_reg[218] = inform_R[217][2];				r_cell_reg[219] = inform_R[221][2];				r_cell_reg[220] = inform_R[218][2];				r_cell_reg[221] = inform_R[222][2];				r_cell_reg[222] = inform_R[219][2];				r_cell_reg[223] = inform_R[223][2];				r_cell_reg[224] = inform_R[224][2];				r_cell_reg[225] = inform_R[228][2];				r_cell_reg[226] = inform_R[225][2];				r_cell_reg[227] = inform_R[229][2];				r_cell_reg[228] = inform_R[226][2];				r_cell_reg[229] = inform_R[230][2];				r_cell_reg[230] = inform_R[227][2];				r_cell_reg[231] = inform_R[231][2];				r_cell_reg[232] = inform_R[232][2];				r_cell_reg[233] = inform_R[236][2];				r_cell_reg[234] = inform_R[233][2];				r_cell_reg[235] = inform_R[237][2];				r_cell_reg[236] = inform_R[234][2];				r_cell_reg[237] = inform_R[238][2];				r_cell_reg[238] = inform_R[235][2];				r_cell_reg[239] = inform_R[239][2];				r_cell_reg[240] = inform_R[240][2];				r_cell_reg[241] = inform_R[244][2];				r_cell_reg[242] = inform_R[241][2];				r_cell_reg[243] = inform_R[245][2];				r_cell_reg[244] = inform_R[242][2];				r_cell_reg[245] = inform_R[246][2];				r_cell_reg[246] = inform_R[243][2];				r_cell_reg[247] = inform_R[247][2];				r_cell_reg[248] = inform_R[248][2];				r_cell_reg[249] = inform_R[252][2];				r_cell_reg[250] = inform_R[249][2];				r_cell_reg[251] = inform_R[253][2];				r_cell_reg[252] = inform_R[250][2];				r_cell_reg[253] = inform_R[254][2];				r_cell_reg[254] = inform_R[251][2];				r_cell_reg[255] = inform_R[255][2];				r_cell_reg[256] = inform_R[256][2];				r_cell_reg[257] = inform_R[260][2];				r_cell_reg[258] = inform_R[257][2];				r_cell_reg[259] = inform_R[261][2];				r_cell_reg[260] = inform_R[258][2];				r_cell_reg[261] = inform_R[262][2];				r_cell_reg[262] = inform_R[259][2];				r_cell_reg[263] = inform_R[263][2];				r_cell_reg[264] = inform_R[264][2];				r_cell_reg[265] = inform_R[268][2];				r_cell_reg[266] = inform_R[265][2];				r_cell_reg[267] = inform_R[269][2];				r_cell_reg[268] = inform_R[266][2];				r_cell_reg[269] = inform_R[270][2];				r_cell_reg[270] = inform_R[267][2];				r_cell_reg[271] = inform_R[271][2];				r_cell_reg[272] = inform_R[272][2];				r_cell_reg[273] = inform_R[276][2];				r_cell_reg[274] = inform_R[273][2];				r_cell_reg[275] = inform_R[277][2];				r_cell_reg[276] = inform_R[274][2];				r_cell_reg[277] = inform_R[278][2];				r_cell_reg[278] = inform_R[275][2];				r_cell_reg[279] = inform_R[279][2];				r_cell_reg[280] = inform_R[280][2];				r_cell_reg[281] = inform_R[284][2];				r_cell_reg[282] = inform_R[281][2];				r_cell_reg[283] = inform_R[285][2];				r_cell_reg[284] = inform_R[282][2];				r_cell_reg[285] = inform_R[286][2];				r_cell_reg[286] = inform_R[283][2];				r_cell_reg[287] = inform_R[287][2];				r_cell_reg[288] = inform_R[288][2];				r_cell_reg[289] = inform_R[292][2];				r_cell_reg[290] = inform_R[289][2];				r_cell_reg[291] = inform_R[293][2];				r_cell_reg[292] = inform_R[290][2];				r_cell_reg[293] = inform_R[294][2];				r_cell_reg[294] = inform_R[291][2];				r_cell_reg[295] = inform_R[295][2];				r_cell_reg[296] = inform_R[296][2];				r_cell_reg[297] = inform_R[300][2];				r_cell_reg[298] = inform_R[297][2];				r_cell_reg[299] = inform_R[301][2];				r_cell_reg[300] = inform_R[298][2];				r_cell_reg[301] = inform_R[302][2];				r_cell_reg[302] = inform_R[299][2];				r_cell_reg[303] = inform_R[303][2];				r_cell_reg[304] = inform_R[304][2];				r_cell_reg[305] = inform_R[308][2];				r_cell_reg[306] = inform_R[305][2];				r_cell_reg[307] = inform_R[309][2];				r_cell_reg[308] = inform_R[306][2];				r_cell_reg[309] = inform_R[310][2];				r_cell_reg[310] = inform_R[307][2];				r_cell_reg[311] = inform_R[311][2];				r_cell_reg[312] = inform_R[312][2];				r_cell_reg[313] = inform_R[316][2];				r_cell_reg[314] = inform_R[313][2];				r_cell_reg[315] = inform_R[317][2];				r_cell_reg[316] = inform_R[314][2];				r_cell_reg[317] = inform_R[318][2];				r_cell_reg[318] = inform_R[315][2];				r_cell_reg[319] = inform_R[319][2];				r_cell_reg[320] = inform_R[320][2];				r_cell_reg[321] = inform_R[324][2];				r_cell_reg[322] = inform_R[321][2];				r_cell_reg[323] = inform_R[325][2];				r_cell_reg[324] = inform_R[322][2];				r_cell_reg[325] = inform_R[326][2];				r_cell_reg[326] = inform_R[323][2];				r_cell_reg[327] = inform_R[327][2];				r_cell_reg[328] = inform_R[328][2];				r_cell_reg[329] = inform_R[332][2];				r_cell_reg[330] = inform_R[329][2];				r_cell_reg[331] = inform_R[333][2];				r_cell_reg[332] = inform_R[330][2];				r_cell_reg[333] = inform_R[334][2];				r_cell_reg[334] = inform_R[331][2];				r_cell_reg[335] = inform_R[335][2];				r_cell_reg[336] = inform_R[336][2];				r_cell_reg[337] = inform_R[340][2];				r_cell_reg[338] = inform_R[337][2];				r_cell_reg[339] = inform_R[341][2];				r_cell_reg[340] = inform_R[338][2];				r_cell_reg[341] = inform_R[342][2];				r_cell_reg[342] = inform_R[339][2];				r_cell_reg[343] = inform_R[343][2];				r_cell_reg[344] = inform_R[344][2];				r_cell_reg[345] = inform_R[348][2];				r_cell_reg[346] = inform_R[345][2];				r_cell_reg[347] = inform_R[349][2];				r_cell_reg[348] = inform_R[346][2];				r_cell_reg[349] = inform_R[350][2];				r_cell_reg[350] = inform_R[347][2];				r_cell_reg[351] = inform_R[351][2];				r_cell_reg[352] = inform_R[352][2];				r_cell_reg[353] = inform_R[356][2];				r_cell_reg[354] = inform_R[353][2];				r_cell_reg[355] = inform_R[357][2];				r_cell_reg[356] = inform_R[354][2];				r_cell_reg[357] = inform_R[358][2];				r_cell_reg[358] = inform_R[355][2];				r_cell_reg[359] = inform_R[359][2];				r_cell_reg[360] = inform_R[360][2];				r_cell_reg[361] = inform_R[364][2];				r_cell_reg[362] = inform_R[361][2];				r_cell_reg[363] = inform_R[365][2];				r_cell_reg[364] = inform_R[362][2];				r_cell_reg[365] = inform_R[366][2];				r_cell_reg[366] = inform_R[363][2];				r_cell_reg[367] = inform_R[367][2];				r_cell_reg[368] = inform_R[368][2];				r_cell_reg[369] = inform_R[372][2];				r_cell_reg[370] = inform_R[369][2];				r_cell_reg[371] = inform_R[373][2];				r_cell_reg[372] = inform_R[370][2];				r_cell_reg[373] = inform_R[374][2];				r_cell_reg[374] = inform_R[371][2];				r_cell_reg[375] = inform_R[375][2];				r_cell_reg[376] = inform_R[376][2];				r_cell_reg[377] = inform_R[380][2];				r_cell_reg[378] = inform_R[377][2];				r_cell_reg[379] = inform_R[381][2];				r_cell_reg[380] = inform_R[378][2];				r_cell_reg[381] = inform_R[382][2];				r_cell_reg[382] = inform_R[379][2];				r_cell_reg[383] = inform_R[383][2];				r_cell_reg[384] = inform_R[384][2];				r_cell_reg[385] = inform_R[388][2];				r_cell_reg[386] = inform_R[385][2];				r_cell_reg[387] = inform_R[389][2];				r_cell_reg[388] = inform_R[386][2];				r_cell_reg[389] = inform_R[390][2];				r_cell_reg[390] = inform_R[387][2];				r_cell_reg[391] = inform_R[391][2];				r_cell_reg[392] = inform_R[392][2];				r_cell_reg[393] = inform_R[396][2];				r_cell_reg[394] = inform_R[393][2];				r_cell_reg[395] = inform_R[397][2];				r_cell_reg[396] = inform_R[394][2];				r_cell_reg[397] = inform_R[398][2];				r_cell_reg[398] = inform_R[395][2];				r_cell_reg[399] = inform_R[399][2];				r_cell_reg[400] = inform_R[400][2];				r_cell_reg[401] = inform_R[404][2];				r_cell_reg[402] = inform_R[401][2];				r_cell_reg[403] = inform_R[405][2];				r_cell_reg[404] = inform_R[402][2];				r_cell_reg[405] = inform_R[406][2];				r_cell_reg[406] = inform_R[403][2];				r_cell_reg[407] = inform_R[407][2];				r_cell_reg[408] = inform_R[408][2];				r_cell_reg[409] = inform_R[412][2];				r_cell_reg[410] = inform_R[409][2];				r_cell_reg[411] = inform_R[413][2];				r_cell_reg[412] = inform_R[410][2];				r_cell_reg[413] = inform_R[414][2];				r_cell_reg[414] = inform_R[411][2];				r_cell_reg[415] = inform_R[415][2];				r_cell_reg[416] = inform_R[416][2];				r_cell_reg[417] = inform_R[420][2];				r_cell_reg[418] = inform_R[417][2];				r_cell_reg[419] = inform_R[421][2];				r_cell_reg[420] = inform_R[418][2];				r_cell_reg[421] = inform_R[422][2];				r_cell_reg[422] = inform_R[419][2];				r_cell_reg[423] = inform_R[423][2];				r_cell_reg[424] = inform_R[424][2];				r_cell_reg[425] = inform_R[428][2];				r_cell_reg[426] = inform_R[425][2];				r_cell_reg[427] = inform_R[429][2];				r_cell_reg[428] = inform_R[426][2];				r_cell_reg[429] = inform_R[430][2];				r_cell_reg[430] = inform_R[427][2];				r_cell_reg[431] = inform_R[431][2];				r_cell_reg[432] = inform_R[432][2];				r_cell_reg[433] = inform_R[436][2];				r_cell_reg[434] = inform_R[433][2];				r_cell_reg[435] = inform_R[437][2];				r_cell_reg[436] = inform_R[434][2];				r_cell_reg[437] = inform_R[438][2];				r_cell_reg[438] = inform_R[435][2];				r_cell_reg[439] = inform_R[439][2];				r_cell_reg[440] = inform_R[440][2];				r_cell_reg[441] = inform_R[444][2];				r_cell_reg[442] = inform_R[441][2];				r_cell_reg[443] = inform_R[445][2];				r_cell_reg[444] = inform_R[442][2];				r_cell_reg[445] = inform_R[446][2];				r_cell_reg[446] = inform_R[443][2];				r_cell_reg[447] = inform_R[447][2];				r_cell_reg[448] = inform_R[448][2];				r_cell_reg[449] = inform_R[452][2];				r_cell_reg[450] = inform_R[449][2];				r_cell_reg[451] = inform_R[453][2];				r_cell_reg[452] = inform_R[450][2];				r_cell_reg[453] = inform_R[454][2];				r_cell_reg[454] = inform_R[451][2];				r_cell_reg[455] = inform_R[455][2];				r_cell_reg[456] = inform_R[456][2];				r_cell_reg[457] = inform_R[460][2];				r_cell_reg[458] = inform_R[457][2];				r_cell_reg[459] = inform_R[461][2];				r_cell_reg[460] = inform_R[458][2];				r_cell_reg[461] = inform_R[462][2];				r_cell_reg[462] = inform_R[459][2];				r_cell_reg[463] = inform_R[463][2];				r_cell_reg[464] = inform_R[464][2];				r_cell_reg[465] = inform_R[468][2];				r_cell_reg[466] = inform_R[465][2];				r_cell_reg[467] = inform_R[469][2];				r_cell_reg[468] = inform_R[466][2];				r_cell_reg[469] = inform_R[470][2];				r_cell_reg[470] = inform_R[467][2];				r_cell_reg[471] = inform_R[471][2];				r_cell_reg[472] = inform_R[472][2];				r_cell_reg[473] = inform_R[476][2];				r_cell_reg[474] = inform_R[473][2];				r_cell_reg[475] = inform_R[477][2];				r_cell_reg[476] = inform_R[474][2];				r_cell_reg[477] = inform_R[478][2];				r_cell_reg[478] = inform_R[475][2];				r_cell_reg[479] = inform_R[479][2];				r_cell_reg[480] = inform_R[480][2];				r_cell_reg[481] = inform_R[484][2];				r_cell_reg[482] = inform_R[481][2];				r_cell_reg[483] = inform_R[485][2];				r_cell_reg[484] = inform_R[482][2];				r_cell_reg[485] = inform_R[486][2];				r_cell_reg[486] = inform_R[483][2];				r_cell_reg[487] = inform_R[487][2];				r_cell_reg[488] = inform_R[488][2];				r_cell_reg[489] = inform_R[492][2];				r_cell_reg[490] = inform_R[489][2];				r_cell_reg[491] = inform_R[493][2];				r_cell_reg[492] = inform_R[490][2];				r_cell_reg[493] = inform_R[494][2];				r_cell_reg[494] = inform_R[491][2];				r_cell_reg[495] = inform_R[495][2];				r_cell_reg[496] = inform_R[496][2];				r_cell_reg[497] = inform_R[500][2];				r_cell_reg[498] = inform_R[497][2];				r_cell_reg[499] = inform_R[501][2];				r_cell_reg[500] = inform_R[498][2];				r_cell_reg[501] = inform_R[502][2];				r_cell_reg[502] = inform_R[499][2];				r_cell_reg[503] = inform_R[503][2];				r_cell_reg[504] = inform_R[504][2];				r_cell_reg[505] = inform_R[508][2];				r_cell_reg[506] = inform_R[505][2];				r_cell_reg[507] = inform_R[509][2];				r_cell_reg[508] = inform_R[506][2];				r_cell_reg[509] = inform_R[510][2];				r_cell_reg[510] = inform_R[507][2];				r_cell_reg[511] = inform_R[511][2];				r_cell_reg[512] = inform_R[512][2];				r_cell_reg[513] = inform_R[516][2];				r_cell_reg[514] = inform_R[513][2];				r_cell_reg[515] = inform_R[517][2];				r_cell_reg[516] = inform_R[514][2];				r_cell_reg[517] = inform_R[518][2];				r_cell_reg[518] = inform_R[515][2];				r_cell_reg[519] = inform_R[519][2];				r_cell_reg[520] = inform_R[520][2];				r_cell_reg[521] = inform_R[524][2];				r_cell_reg[522] = inform_R[521][2];				r_cell_reg[523] = inform_R[525][2];				r_cell_reg[524] = inform_R[522][2];				r_cell_reg[525] = inform_R[526][2];				r_cell_reg[526] = inform_R[523][2];				r_cell_reg[527] = inform_R[527][2];				r_cell_reg[528] = inform_R[528][2];				r_cell_reg[529] = inform_R[532][2];				r_cell_reg[530] = inform_R[529][2];				r_cell_reg[531] = inform_R[533][2];				r_cell_reg[532] = inform_R[530][2];				r_cell_reg[533] = inform_R[534][2];				r_cell_reg[534] = inform_R[531][2];				r_cell_reg[535] = inform_R[535][2];				r_cell_reg[536] = inform_R[536][2];				r_cell_reg[537] = inform_R[540][2];				r_cell_reg[538] = inform_R[537][2];				r_cell_reg[539] = inform_R[541][2];				r_cell_reg[540] = inform_R[538][2];				r_cell_reg[541] = inform_R[542][2];				r_cell_reg[542] = inform_R[539][2];				r_cell_reg[543] = inform_R[543][2];				r_cell_reg[544] = inform_R[544][2];				r_cell_reg[545] = inform_R[548][2];				r_cell_reg[546] = inform_R[545][2];				r_cell_reg[547] = inform_R[549][2];				r_cell_reg[548] = inform_R[546][2];				r_cell_reg[549] = inform_R[550][2];				r_cell_reg[550] = inform_R[547][2];				r_cell_reg[551] = inform_R[551][2];				r_cell_reg[552] = inform_R[552][2];				r_cell_reg[553] = inform_R[556][2];				r_cell_reg[554] = inform_R[553][2];				r_cell_reg[555] = inform_R[557][2];				r_cell_reg[556] = inform_R[554][2];				r_cell_reg[557] = inform_R[558][2];				r_cell_reg[558] = inform_R[555][2];				r_cell_reg[559] = inform_R[559][2];				r_cell_reg[560] = inform_R[560][2];				r_cell_reg[561] = inform_R[564][2];				r_cell_reg[562] = inform_R[561][2];				r_cell_reg[563] = inform_R[565][2];				r_cell_reg[564] = inform_R[562][2];				r_cell_reg[565] = inform_R[566][2];				r_cell_reg[566] = inform_R[563][2];				r_cell_reg[567] = inform_R[567][2];				r_cell_reg[568] = inform_R[568][2];				r_cell_reg[569] = inform_R[572][2];				r_cell_reg[570] = inform_R[569][2];				r_cell_reg[571] = inform_R[573][2];				r_cell_reg[572] = inform_R[570][2];				r_cell_reg[573] = inform_R[574][2];				r_cell_reg[574] = inform_R[571][2];				r_cell_reg[575] = inform_R[575][2];				r_cell_reg[576] = inform_R[576][2];				r_cell_reg[577] = inform_R[580][2];				r_cell_reg[578] = inform_R[577][2];				r_cell_reg[579] = inform_R[581][2];				r_cell_reg[580] = inform_R[578][2];				r_cell_reg[581] = inform_R[582][2];				r_cell_reg[582] = inform_R[579][2];				r_cell_reg[583] = inform_R[583][2];				r_cell_reg[584] = inform_R[584][2];				r_cell_reg[585] = inform_R[588][2];				r_cell_reg[586] = inform_R[585][2];				r_cell_reg[587] = inform_R[589][2];				r_cell_reg[588] = inform_R[586][2];				r_cell_reg[589] = inform_R[590][2];				r_cell_reg[590] = inform_R[587][2];				r_cell_reg[591] = inform_R[591][2];				r_cell_reg[592] = inform_R[592][2];				r_cell_reg[593] = inform_R[596][2];				r_cell_reg[594] = inform_R[593][2];				r_cell_reg[595] = inform_R[597][2];				r_cell_reg[596] = inform_R[594][2];				r_cell_reg[597] = inform_R[598][2];				r_cell_reg[598] = inform_R[595][2];				r_cell_reg[599] = inform_R[599][2];				r_cell_reg[600] = inform_R[600][2];				r_cell_reg[601] = inform_R[604][2];				r_cell_reg[602] = inform_R[601][2];				r_cell_reg[603] = inform_R[605][2];				r_cell_reg[604] = inform_R[602][2];				r_cell_reg[605] = inform_R[606][2];				r_cell_reg[606] = inform_R[603][2];				r_cell_reg[607] = inform_R[607][2];				r_cell_reg[608] = inform_R[608][2];				r_cell_reg[609] = inform_R[612][2];				r_cell_reg[610] = inform_R[609][2];				r_cell_reg[611] = inform_R[613][2];				r_cell_reg[612] = inform_R[610][2];				r_cell_reg[613] = inform_R[614][2];				r_cell_reg[614] = inform_R[611][2];				r_cell_reg[615] = inform_R[615][2];				r_cell_reg[616] = inform_R[616][2];				r_cell_reg[617] = inform_R[620][2];				r_cell_reg[618] = inform_R[617][2];				r_cell_reg[619] = inform_R[621][2];				r_cell_reg[620] = inform_R[618][2];				r_cell_reg[621] = inform_R[622][2];				r_cell_reg[622] = inform_R[619][2];				r_cell_reg[623] = inform_R[623][2];				r_cell_reg[624] = inform_R[624][2];				r_cell_reg[625] = inform_R[628][2];				r_cell_reg[626] = inform_R[625][2];				r_cell_reg[627] = inform_R[629][2];				r_cell_reg[628] = inform_R[626][2];				r_cell_reg[629] = inform_R[630][2];				r_cell_reg[630] = inform_R[627][2];				r_cell_reg[631] = inform_R[631][2];				r_cell_reg[632] = inform_R[632][2];				r_cell_reg[633] = inform_R[636][2];				r_cell_reg[634] = inform_R[633][2];				r_cell_reg[635] = inform_R[637][2];				r_cell_reg[636] = inform_R[634][2];				r_cell_reg[637] = inform_R[638][2];				r_cell_reg[638] = inform_R[635][2];				r_cell_reg[639] = inform_R[639][2];				r_cell_reg[640] = inform_R[640][2];				r_cell_reg[641] = inform_R[644][2];				r_cell_reg[642] = inform_R[641][2];				r_cell_reg[643] = inform_R[645][2];				r_cell_reg[644] = inform_R[642][2];				r_cell_reg[645] = inform_R[646][2];				r_cell_reg[646] = inform_R[643][2];				r_cell_reg[647] = inform_R[647][2];				r_cell_reg[648] = inform_R[648][2];				r_cell_reg[649] = inform_R[652][2];				r_cell_reg[650] = inform_R[649][2];				r_cell_reg[651] = inform_R[653][2];				r_cell_reg[652] = inform_R[650][2];				r_cell_reg[653] = inform_R[654][2];				r_cell_reg[654] = inform_R[651][2];				r_cell_reg[655] = inform_R[655][2];				r_cell_reg[656] = inform_R[656][2];				r_cell_reg[657] = inform_R[660][2];				r_cell_reg[658] = inform_R[657][2];				r_cell_reg[659] = inform_R[661][2];				r_cell_reg[660] = inform_R[658][2];				r_cell_reg[661] = inform_R[662][2];				r_cell_reg[662] = inform_R[659][2];				r_cell_reg[663] = inform_R[663][2];				r_cell_reg[664] = inform_R[664][2];				r_cell_reg[665] = inform_R[668][2];				r_cell_reg[666] = inform_R[665][2];				r_cell_reg[667] = inform_R[669][2];				r_cell_reg[668] = inform_R[666][2];				r_cell_reg[669] = inform_R[670][2];				r_cell_reg[670] = inform_R[667][2];				r_cell_reg[671] = inform_R[671][2];				r_cell_reg[672] = inform_R[672][2];				r_cell_reg[673] = inform_R[676][2];				r_cell_reg[674] = inform_R[673][2];				r_cell_reg[675] = inform_R[677][2];				r_cell_reg[676] = inform_R[674][2];				r_cell_reg[677] = inform_R[678][2];				r_cell_reg[678] = inform_R[675][2];				r_cell_reg[679] = inform_R[679][2];				r_cell_reg[680] = inform_R[680][2];				r_cell_reg[681] = inform_R[684][2];				r_cell_reg[682] = inform_R[681][2];				r_cell_reg[683] = inform_R[685][2];				r_cell_reg[684] = inform_R[682][2];				r_cell_reg[685] = inform_R[686][2];				r_cell_reg[686] = inform_R[683][2];				r_cell_reg[687] = inform_R[687][2];				r_cell_reg[688] = inform_R[688][2];				r_cell_reg[689] = inform_R[692][2];				r_cell_reg[690] = inform_R[689][2];				r_cell_reg[691] = inform_R[693][2];				r_cell_reg[692] = inform_R[690][2];				r_cell_reg[693] = inform_R[694][2];				r_cell_reg[694] = inform_R[691][2];				r_cell_reg[695] = inform_R[695][2];				r_cell_reg[696] = inform_R[696][2];				r_cell_reg[697] = inform_R[700][2];				r_cell_reg[698] = inform_R[697][2];				r_cell_reg[699] = inform_R[701][2];				r_cell_reg[700] = inform_R[698][2];				r_cell_reg[701] = inform_R[702][2];				r_cell_reg[702] = inform_R[699][2];				r_cell_reg[703] = inform_R[703][2];				r_cell_reg[704] = inform_R[704][2];				r_cell_reg[705] = inform_R[708][2];				r_cell_reg[706] = inform_R[705][2];				r_cell_reg[707] = inform_R[709][2];				r_cell_reg[708] = inform_R[706][2];				r_cell_reg[709] = inform_R[710][2];				r_cell_reg[710] = inform_R[707][2];				r_cell_reg[711] = inform_R[711][2];				r_cell_reg[712] = inform_R[712][2];				r_cell_reg[713] = inform_R[716][2];				r_cell_reg[714] = inform_R[713][2];				r_cell_reg[715] = inform_R[717][2];				r_cell_reg[716] = inform_R[714][2];				r_cell_reg[717] = inform_R[718][2];				r_cell_reg[718] = inform_R[715][2];				r_cell_reg[719] = inform_R[719][2];				r_cell_reg[720] = inform_R[720][2];				r_cell_reg[721] = inform_R[724][2];				r_cell_reg[722] = inform_R[721][2];				r_cell_reg[723] = inform_R[725][2];				r_cell_reg[724] = inform_R[722][2];				r_cell_reg[725] = inform_R[726][2];				r_cell_reg[726] = inform_R[723][2];				r_cell_reg[727] = inform_R[727][2];				r_cell_reg[728] = inform_R[728][2];				r_cell_reg[729] = inform_R[732][2];				r_cell_reg[730] = inform_R[729][2];				r_cell_reg[731] = inform_R[733][2];				r_cell_reg[732] = inform_R[730][2];				r_cell_reg[733] = inform_R[734][2];				r_cell_reg[734] = inform_R[731][2];				r_cell_reg[735] = inform_R[735][2];				r_cell_reg[736] = inform_R[736][2];				r_cell_reg[737] = inform_R[740][2];				r_cell_reg[738] = inform_R[737][2];				r_cell_reg[739] = inform_R[741][2];				r_cell_reg[740] = inform_R[738][2];				r_cell_reg[741] = inform_R[742][2];				r_cell_reg[742] = inform_R[739][2];				r_cell_reg[743] = inform_R[743][2];				r_cell_reg[744] = inform_R[744][2];				r_cell_reg[745] = inform_R[748][2];				r_cell_reg[746] = inform_R[745][2];				r_cell_reg[747] = inform_R[749][2];				r_cell_reg[748] = inform_R[746][2];				r_cell_reg[749] = inform_R[750][2];				r_cell_reg[750] = inform_R[747][2];				r_cell_reg[751] = inform_R[751][2];				r_cell_reg[752] = inform_R[752][2];				r_cell_reg[753] = inform_R[756][2];				r_cell_reg[754] = inform_R[753][2];				r_cell_reg[755] = inform_R[757][2];				r_cell_reg[756] = inform_R[754][2];				r_cell_reg[757] = inform_R[758][2];				r_cell_reg[758] = inform_R[755][2];				r_cell_reg[759] = inform_R[759][2];				r_cell_reg[760] = inform_R[760][2];				r_cell_reg[761] = inform_R[764][2];				r_cell_reg[762] = inform_R[761][2];				r_cell_reg[763] = inform_R[765][2];				r_cell_reg[764] = inform_R[762][2];				r_cell_reg[765] = inform_R[766][2];				r_cell_reg[766] = inform_R[763][2];				r_cell_reg[767] = inform_R[767][2];				r_cell_reg[768] = inform_R[768][2];				r_cell_reg[769] = inform_R[772][2];				r_cell_reg[770] = inform_R[769][2];				r_cell_reg[771] = inform_R[773][2];				r_cell_reg[772] = inform_R[770][2];				r_cell_reg[773] = inform_R[774][2];				r_cell_reg[774] = inform_R[771][2];				r_cell_reg[775] = inform_R[775][2];				r_cell_reg[776] = inform_R[776][2];				r_cell_reg[777] = inform_R[780][2];				r_cell_reg[778] = inform_R[777][2];				r_cell_reg[779] = inform_R[781][2];				r_cell_reg[780] = inform_R[778][2];				r_cell_reg[781] = inform_R[782][2];				r_cell_reg[782] = inform_R[779][2];				r_cell_reg[783] = inform_R[783][2];				r_cell_reg[784] = inform_R[784][2];				r_cell_reg[785] = inform_R[788][2];				r_cell_reg[786] = inform_R[785][2];				r_cell_reg[787] = inform_R[789][2];				r_cell_reg[788] = inform_R[786][2];				r_cell_reg[789] = inform_R[790][2];				r_cell_reg[790] = inform_R[787][2];				r_cell_reg[791] = inform_R[791][2];				r_cell_reg[792] = inform_R[792][2];				r_cell_reg[793] = inform_R[796][2];				r_cell_reg[794] = inform_R[793][2];				r_cell_reg[795] = inform_R[797][2];				r_cell_reg[796] = inform_R[794][2];				r_cell_reg[797] = inform_R[798][2];				r_cell_reg[798] = inform_R[795][2];				r_cell_reg[799] = inform_R[799][2];				r_cell_reg[800] = inform_R[800][2];				r_cell_reg[801] = inform_R[804][2];				r_cell_reg[802] = inform_R[801][2];				r_cell_reg[803] = inform_R[805][2];				r_cell_reg[804] = inform_R[802][2];				r_cell_reg[805] = inform_R[806][2];				r_cell_reg[806] = inform_R[803][2];				r_cell_reg[807] = inform_R[807][2];				r_cell_reg[808] = inform_R[808][2];				r_cell_reg[809] = inform_R[812][2];				r_cell_reg[810] = inform_R[809][2];				r_cell_reg[811] = inform_R[813][2];				r_cell_reg[812] = inform_R[810][2];				r_cell_reg[813] = inform_R[814][2];				r_cell_reg[814] = inform_R[811][2];				r_cell_reg[815] = inform_R[815][2];				r_cell_reg[816] = inform_R[816][2];				r_cell_reg[817] = inform_R[820][2];				r_cell_reg[818] = inform_R[817][2];				r_cell_reg[819] = inform_R[821][2];				r_cell_reg[820] = inform_R[818][2];				r_cell_reg[821] = inform_R[822][2];				r_cell_reg[822] = inform_R[819][2];				r_cell_reg[823] = inform_R[823][2];				r_cell_reg[824] = inform_R[824][2];				r_cell_reg[825] = inform_R[828][2];				r_cell_reg[826] = inform_R[825][2];				r_cell_reg[827] = inform_R[829][2];				r_cell_reg[828] = inform_R[826][2];				r_cell_reg[829] = inform_R[830][2];				r_cell_reg[830] = inform_R[827][2];				r_cell_reg[831] = inform_R[831][2];				r_cell_reg[832] = inform_R[832][2];				r_cell_reg[833] = inform_R[836][2];				r_cell_reg[834] = inform_R[833][2];				r_cell_reg[835] = inform_R[837][2];				r_cell_reg[836] = inform_R[834][2];				r_cell_reg[837] = inform_R[838][2];				r_cell_reg[838] = inform_R[835][2];				r_cell_reg[839] = inform_R[839][2];				r_cell_reg[840] = inform_R[840][2];				r_cell_reg[841] = inform_R[844][2];				r_cell_reg[842] = inform_R[841][2];				r_cell_reg[843] = inform_R[845][2];				r_cell_reg[844] = inform_R[842][2];				r_cell_reg[845] = inform_R[846][2];				r_cell_reg[846] = inform_R[843][2];				r_cell_reg[847] = inform_R[847][2];				r_cell_reg[848] = inform_R[848][2];				r_cell_reg[849] = inform_R[852][2];				r_cell_reg[850] = inform_R[849][2];				r_cell_reg[851] = inform_R[853][2];				r_cell_reg[852] = inform_R[850][2];				r_cell_reg[853] = inform_R[854][2];				r_cell_reg[854] = inform_R[851][2];				r_cell_reg[855] = inform_R[855][2];				r_cell_reg[856] = inform_R[856][2];				r_cell_reg[857] = inform_R[860][2];				r_cell_reg[858] = inform_R[857][2];				r_cell_reg[859] = inform_R[861][2];				r_cell_reg[860] = inform_R[858][2];				r_cell_reg[861] = inform_R[862][2];				r_cell_reg[862] = inform_R[859][2];				r_cell_reg[863] = inform_R[863][2];				r_cell_reg[864] = inform_R[864][2];				r_cell_reg[865] = inform_R[868][2];				r_cell_reg[866] = inform_R[865][2];				r_cell_reg[867] = inform_R[869][2];				r_cell_reg[868] = inform_R[866][2];				r_cell_reg[869] = inform_R[870][2];				r_cell_reg[870] = inform_R[867][2];				r_cell_reg[871] = inform_R[871][2];				r_cell_reg[872] = inform_R[872][2];				r_cell_reg[873] = inform_R[876][2];				r_cell_reg[874] = inform_R[873][2];				r_cell_reg[875] = inform_R[877][2];				r_cell_reg[876] = inform_R[874][2];				r_cell_reg[877] = inform_R[878][2];				r_cell_reg[878] = inform_R[875][2];				r_cell_reg[879] = inform_R[879][2];				r_cell_reg[880] = inform_R[880][2];				r_cell_reg[881] = inform_R[884][2];				r_cell_reg[882] = inform_R[881][2];				r_cell_reg[883] = inform_R[885][2];				r_cell_reg[884] = inform_R[882][2];				r_cell_reg[885] = inform_R[886][2];				r_cell_reg[886] = inform_R[883][2];				r_cell_reg[887] = inform_R[887][2];				r_cell_reg[888] = inform_R[888][2];				r_cell_reg[889] = inform_R[892][2];				r_cell_reg[890] = inform_R[889][2];				r_cell_reg[891] = inform_R[893][2];				r_cell_reg[892] = inform_R[890][2];				r_cell_reg[893] = inform_R[894][2];				r_cell_reg[894] = inform_R[891][2];				r_cell_reg[895] = inform_R[895][2];				r_cell_reg[896] = inform_R[896][2];				r_cell_reg[897] = inform_R[900][2];				r_cell_reg[898] = inform_R[897][2];				r_cell_reg[899] = inform_R[901][2];				r_cell_reg[900] = inform_R[898][2];				r_cell_reg[901] = inform_R[902][2];				r_cell_reg[902] = inform_R[899][2];				r_cell_reg[903] = inform_R[903][2];				r_cell_reg[904] = inform_R[904][2];				r_cell_reg[905] = inform_R[908][2];				r_cell_reg[906] = inform_R[905][2];				r_cell_reg[907] = inform_R[909][2];				r_cell_reg[908] = inform_R[906][2];				r_cell_reg[909] = inform_R[910][2];				r_cell_reg[910] = inform_R[907][2];				r_cell_reg[911] = inform_R[911][2];				r_cell_reg[912] = inform_R[912][2];				r_cell_reg[913] = inform_R[916][2];				r_cell_reg[914] = inform_R[913][2];				r_cell_reg[915] = inform_R[917][2];				r_cell_reg[916] = inform_R[914][2];				r_cell_reg[917] = inform_R[918][2];				r_cell_reg[918] = inform_R[915][2];				r_cell_reg[919] = inform_R[919][2];				r_cell_reg[920] = inform_R[920][2];				r_cell_reg[921] = inform_R[924][2];				r_cell_reg[922] = inform_R[921][2];				r_cell_reg[923] = inform_R[925][2];				r_cell_reg[924] = inform_R[922][2];				r_cell_reg[925] = inform_R[926][2];				r_cell_reg[926] = inform_R[923][2];				r_cell_reg[927] = inform_R[927][2];				r_cell_reg[928] = inform_R[928][2];				r_cell_reg[929] = inform_R[932][2];				r_cell_reg[930] = inform_R[929][2];				r_cell_reg[931] = inform_R[933][2];				r_cell_reg[932] = inform_R[930][2];				r_cell_reg[933] = inform_R[934][2];				r_cell_reg[934] = inform_R[931][2];				r_cell_reg[935] = inform_R[935][2];				r_cell_reg[936] = inform_R[936][2];				r_cell_reg[937] = inform_R[940][2];				r_cell_reg[938] = inform_R[937][2];				r_cell_reg[939] = inform_R[941][2];				r_cell_reg[940] = inform_R[938][2];				r_cell_reg[941] = inform_R[942][2];				r_cell_reg[942] = inform_R[939][2];				r_cell_reg[943] = inform_R[943][2];				r_cell_reg[944] = inform_R[944][2];				r_cell_reg[945] = inform_R[948][2];				r_cell_reg[946] = inform_R[945][2];				r_cell_reg[947] = inform_R[949][2];				r_cell_reg[948] = inform_R[946][2];				r_cell_reg[949] = inform_R[950][2];				r_cell_reg[950] = inform_R[947][2];				r_cell_reg[951] = inform_R[951][2];				r_cell_reg[952] = inform_R[952][2];				r_cell_reg[953] = inform_R[956][2];				r_cell_reg[954] = inform_R[953][2];				r_cell_reg[955] = inform_R[957][2];				r_cell_reg[956] = inform_R[954][2];				r_cell_reg[957] = inform_R[958][2];				r_cell_reg[958] = inform_R[955][2];				r_cell_reg[959] = inform_R[959][2];				r_cell_reg[960] = inform_R[960][2];				r_cell_reg[961] = inform_R[964][2];				r_cell_reg[962] = inform_R[961][2];				r_cell_reg[963] = inform_R[965][2];				r_cell_reg[964] = inform_R[962][2];				r_cell_reg[965] = inform_R[966][2];				r_cell_reg[966] = inform_R[963][2];				r_cell_reg[967] = inform_R[967][2];				r_cell_reg[968] = inform_R[968][2];				r_cell_reg[969] = inform_R[972][2];				r_cell_reg[970] = inform_R[969][2];				r_cell_reg[971] = inform_R[973][2];				r_cell_reg[972] = inform_R[970][2];				r_cell_reg[973] = inform_R[974][2];				r_cell_reg[974] = inform_R[971][2];				r_cell_reg[975] = inform_R[975][2];				r_cell_reg[976] = inform_R[976][2];				r_cell_reg[977] = inform_R[980][2];				r_cell_reg[978] = inform_R[977][2];				r_cell_reg[979] = inform_R[981][2];				r_cell_reg[980] = inform_R[978][2];				r_cell_reg[981] = inform_R[982][2];				r_cell_reg[982] = inform_R[979][2];				r_cell_reg[983] = inform_R[983][2];				r_cell_reg[984] = inform_R[984][2];				r_cell_reg[985] = inform_R[988][2];				r_cell_reg[986] = inform_R[985][2];				r_cell_reg[987] = inform_R[989][2];				r_cell_reg[988] = inform_R[986][2];				r_cell_reg[989] = inform_R[990][2];				r_cell_reg[990] = inform_R[987][2];				r_cell_reg[991] = inform_R[991][2];				r_cell_reg[992] = inform_R[992][2];				r_cell_reg[993] = inform_R[996][2];				r_cell_reg[994] = inform_R[993][2];				r_cell_reg[995] = inform_R[997][2];				r_cell_reg[996] = inform_R[994][2];				r_cell_reg[997] = inform_R[998][2];				r_cell_reg[998] = inform_R[995][2];				r_cell_reg[999] = inform_R[999][2];				r_cell_reg[1000] = inform_R[1000][2];				r_cell_reg[1001] = inform_R[1004][2];				r_cell_reg[1002] = inform_R[1001][2];				r_cell_reg[1003] = inform_R[1005][2];				r_cell_reg[1004] = inform_R[1002][2];				r_cell_reg[1005] = inform_R[1006][2];				r_cell_reg[1006] = inform_R[1003][2];				r_cell_reg[1007] = inform_R[1007][2];				r_cell_reg[1008] = inform_R[1008][2];				r_cell_reg[1009] = inform_R[1012][2];				r_cell_reg[1010] = inform_R[1009][2];				r_cell_reg[1011] = inform_R[1013][2];				r_cell_reg[1012] = inform_R[1010][2];				r_cell_reg[1013] = inform_R[1014][2];				r_cell_reg[1014] = inform_R[1011][2];				r_cell_reg[1015] = inform_R[1015][2];				r_cell_reg[1016] = inform_R[1016][2];				r_cell_reg[1017] = inform_R[1020][2];				r_cell_reg[1018] = inform_R[1017][2];				r_cell_reg[1019] = inform_R[1021][2];				r_cell_reg[1020] = inform_R[1018][2];				r_cell_reg[1021] = inform_R[1022][2];				r_cell_reg[1022] = inform_R[1019][2];				r_cell_reg[1023] = inform_R[1023][2];				l_cell_reg[0] = inform_L[0][3];				l_cell_reg[1] = inform_L[4][3];				l_cell_reg[2] = inform_L[1][3];				l_cell_reg[3] = inform_L[5][3];				l_cell_reg[4] = inform_L[2][3];				l_cell_reg[5] = inform_L[6][3];				l_cell_reg[6] = inform_L[3][3];				l_cell_reg[7] = inform_L[7][3];				l_cell_reg[8] = inform_L[8][3];				l_cell_reg[9] = inform_L[12][3];				l_cell_reg[10] = inform_L[9][3];				l_cell_reg[11] = inform_L[13][3];				l_cell_reg[12] = inform_L[10][3];				l_cell_reg[13] = inform_L[14][3];				l_cell_reg[14] = inform_L[11][3];				l_cell_reg[15] = inform_L[15][3];				l_cell_reg[16] = inform_L[16][3];				l_cell_reg[17] = inform_L[20][3];				l_cell_reg[18] = inform_L[17][3];				l_cell_reg[19] = inform_L[21][3];				l_cell_reg[20] = inform_L[18][3];				l_cell_reg[21] = inform_L[22][3];				l_cell_reg[22] = inform_L[19][3];				l_cell_reg[23] = inform_L[23][3];				l_cell_reg[24] = inform_L[24][3];				l_cell_reg[25] = inform_L[28][3];				l_cell_reg[26] = inform_L[25][3];				l_cell_reg[27] = inform_L[29][3];				l_cell_reg[28] = inform_L[26][3];				l_cell_reg[29] = inform_L[30][3];				l_cell_reg[30] = inform_L[27][3];				l_cell_reg[31] = inform_L[31][3];				l_cell_reg[32] = inform_L[32][3];				l_cell_reg[33] = inform_L[36][3];				l_cell_reg[34] = inform_L[33][3];				l_cell_reg[35] = inform_L[37][3];				l_cell_reg[36] = inform_L[34][3];				l_cell_reg[37] = inform_L[38][3];				l_cell_reg[38] = inform_L[35][3];				l_cell_reg[39] = inform_L[39][3];				l_cell_reg[40] = inform_L[40][3];				l_cell_reg[41] = inform_L[44][3];				l_cell_reg[42] = inform_L[41][3];				l_cell_reg[43] = inform_L[45][3];				l_cell_reg[44] = inform_L[42][3];				l_cell_reg[45] = inform_L[46][3];				l_cell_reg[46] = inform_L[43][3];				l_cell_reg[47] = inform_L[47][3];				l_cell_reg[48] = inform_L[48][3];				l_cell_reg[49] = inform_L[52][3];				l_cell_reg[50] = inform_L[49][3];				l_cell_reg[51] = inform_L[53][3];				l_cell_reg[52] = inform_L[50][3];				l_cell_reg[53] = inform_L[54][3];				l_cell_reg[54] = inform_L[51][3];				l_cell_reg[55] = inform_L[55][3];				l_cell_reg[56] = inform_L[56][3];				l_cell_reg[57] = inform_L[60][3];				l_cell_reg[58] = inform_L[57][3];				l_cell_reg[59] = inform_L[61][3];				l_cell_reg[60] = inform_L[58][3];				l_cell_reg[61] = inform_L[62][3];				l_cell_reg[62] = inform_L[59][3];				l_cell_reg[63] = inform_L[63][3];				l_cell_reg[64] = inform_L[64][3];				l_cell_reg[65] = inform_L[68][3];				l_cell_reg[66] = inform_L[65][3];				l_cell_reg[67] = inform_L[69][3];				l_cell_reg[68] = inform_L[66][3];				l_cell_reg[69] = inform_L[70][3];				l_cell_reg[70] = inform_L[67][3];				l_cell_reg[71] = inform_L[71][3];				l_cell_reg[72] = inform_L[72][3];				l_cell_reg[73] = inform_L[76][3];				l_cell_reg[74] = inform_L[73][3];				l_cell_reg[75] = inform_L[77][3];				l_cell_reg[76] = inform_L[74][3];				l_cell_reg[77] = inform_L[78][3];				l_cell_reg[78] = inform_L[75][3];				l_cell_reg[79] = inform_L[79][3];				l_cell_reg[80] = inform_L[80][3];				l_cell_reg[81] = inform_L[84][3];				l_cell_reg[82] = inform_L[81][3];				l_cell_reg[83] = inform_L[85][3];				l_cell_reg[84] = inform_L[82][3];				l_cell_reg[85] = inform_L[86][3];				l_cell_reg[86] = inform_L[83][3];				l_cell_reg[87] = inform_L[87][3];				l_cell_reg[88] = inform_L[88][3];				l_cell_reg[89] = inform_L[92][3];				l_cell_reg[90] = inform_L[89][3];				l_cell_reg[91] = inform_L[93][3];				l_cell_reg[92] = inform_L[90][3];				l_cell_reg[93] = inform_L[94][3];				l_cell_reg[94] = inform_L[91][3];				l_cell_reg[95] = inform_L[95][3];				l_cell_reg[96] = inform_L[96][3];				l_cell_reg[97] = inform_L[100][3];				l_cell_reg[98] = inform_L[97][3];				l_cell_reg[99] = inform_L[101][3];				l_cell_reg[100] = inform_L[98][3];				l_cell_reg[101] = inform_L[102][3];				l_cell_reg[102] = inform_L[99][3];				l_cell_reg[103] = inform_L[103][3];				l_cell_reg[104] = inform_L[104][3];				l_cell_reg[105] = inform_L[108][3];				l_cell_reg[106] = inform_L[105][3];				l_cell_reg[107] = inform_L[109][3];				l_cell_reg[108] = inform_L[106][3];				l_cell_reg[109] = inform_L[110][3];				l_cell_reg[110] = inform_L[107][3];				l_cell_reg[111] = inform_L[111][3];				l_cell_reg[112] = inform_L[112][3];				l_cell_reg[113] = inform_L[116][3];				l_cell_reg[114] = inform_L[113][3];				l_cell_reg[115] = inform_L[117][3];				l_cell_reg[116] = inform_L[114][3];				l_cell_reg[117] = inform_L[118][3];				l_cell_reg[118] = inform_L[115][3];				l_cell_reg[119] = inform_L[119][3];				l_cell_reg[120] = inform_L[120][3];				l_cell_reg[121] = inform_L[124][3];				l_cell_reg[122] = inform_L[121][3];				l_cell_reg[123] = inform_L[125][3];				l_cell_reg[124] = inform_L[122][3];				l_cell_reg[125] = inform_L[126][3];				l_cell_reg[126] = inform_L[123][3];				l_cell_reg[127] = inform_L[127][3];				l_cell_reg[128] = inform_L[128][3];				l_cell_reg[129] = inform_L[132][3];				l_cell_reg[130] = inform_L[129][3];				l_cell_reg[131] = inform_L[133][3];				l_cell_reg[132] = inform_L[130][3];				l_cell_reg[133] = inform_L[134][3];				l_cell_reg[134] = inform_L[131][3];				l_cell_reg[135] = inform_L[135][3];				l_cell_reg[136] = inform_L[136][3];				l_cell_reg[137] = inform_L[140][3];				l_cell_reg[138] = inform_L[137][3];				l_cell_reg[139] = inform_L[141][3];				l_cell_reg[140] = inform_L[138][3];				l_cell_reg[141] = inform_L[142][3];				l_cell_reg[142] = inform_L[139][3];				l_cell_reg[143] = inform_L[143][3];				l_cell_reg[144] = inform_L[144][3];				l_cell_reg[145] = inform_L[148][3];				l_cell_reg[146] = inform_L[145][3];				l_cell_reg[147] = inform_L[149][3];				l_cell_reg[148] = inform_L[146][3];				l_cell_reg[149] = inform_L[150][3];				l_cell_reg[150] = inform_L[147][3];				l_cell_reg[151] = inform_L[151][3];				l_cell_reg[152] = inform_L[152][3];				l_cell_reg[153] = inform_L[156][3];				l_cell_reg[154] = inform_L[153][3];				l_cell_reg[155] = inform_L[157][3];				l_cell_reg[156] = inform_L[154][3];				l_cell_reg[157] = inform_L[158][3];				l_cell_reg[158] = inform_L[155][3];				l_cell_reg[159] = inform_L[159][3];				l_cell_reg[160] = inform_L[160][3];				l_cell_reg[161] = inform_L[164][3];				l_cell_reg[162] = inform_L[161][3];				l_cell_reg[163] = inform_L[165][3];				l_cell_reg[164] = inform_L[162][3];				l_cell_reg[165] = inform_L[166][3];				l_cell_reg[166] = inform_L[163][3];				l_cell_reg[167] = inform_L[167][3];				l_cell_reg[168] = inform_L[168][3];				l_cell_reg[169] = inform_L[172][3];				l_cell_reg[170] = inform_L[169][3];				l_cell_reg[171] = inform_L[173][3];				l_cell_reg[172] = inform_L[170][3];				l_cell_reg[173] = inform_L[174][3];				l_cell_reg[174] = inform_L[171][3];				l_cell_reg[175] = inform_L[175][3];				l_cell_reg[176] = inform_L[176][3];				l_cell_reg[177] = inform_L[180][3];				l_cell_reg[178] = inform_L[177][3];				l_cell_reg[179] = inform_L[181][3];				l_cell_reg[180] = inform_L[178][3];				l_cell_reg[181] = inform_L[182][3];				l_cell_reg[182] = inform_L[179][3];				l_cell_reg[183] = inform_L[183][3];				l_cell_reg[184] = inform_L[184][3];				l_cell_reg[185] = inform_L[188][3];				l_cell_reg[186] = inform_L[185][3];				l_cell_reg[187] = inform_L[189][3];				l_cell_reg[188] = inform_L[186][3];				l_cell_reg[189] = inform_L[190][3];				l_cell_reg[190] = inform_L[187][3];				l_cell_reg[191] = inform_L[191][3];				l_cell_reg[192] = inform_L[192][3];				l_cell_reg[193] = inform_L[196][3];				l_cell_reg[194] = inform_L[193][3];				l_cell_reg[195] = inform_L[197][3];				l_cell_reg[196] = inform_L[194][3];				l_cell_reg[197] = inform_L[198][3];				l_cell_reg[198] = inform_L[195][3];				l_cell_reg[199] = inform_L[199][3];				l_cell_reg[200] = inform_L[200][3];				l_cell_reg[201] = inform_L[204][3];				l_cell_reg[202] = inform_L[201][3];				l_cell_reg[203] = inform_L[205][3];				l_cell_reg[204] = inform_L[202][3];				l_cell_reg[205] = inform_L[206][3];				l_cell_reg[206] = inform_L[203][3];				l_cell_reg[207] = inform_L[207][3];				l_cell_reg[208] = inform_L[208][3];				l_cell_reg[209] = inform_L[212][3];				l_cell_reg[210] = inform_L[209][3];				l_cell_reg[211] = inform_L[213][3];				l_cell_reg[212] = inform_L[210][3];				l_cell_reg[213] = inform_L[214][3];				l_cell_reg[214] = inform_L[211][3];				l_cell_reg[215] = inform_L[215][3];				l_cell_reg[216] = inform_L[216][3];				l_cell_reg[217] = inform_L[220][3];				l_cell_reg[218] = inform_L[217][3];				l_cell_reg[219] = inform_L[221][3];				l_cell_reg[220] = inform_L[218][3];				l_cell_reg[221] = inform_L[222][3];				l_cell_reg[222] = inform_L[219][3];				l_cell_reg[223] = inform_L[223][3];				l_cell_reg[224] = inform_L[224][3];				l_cell_reg[225] = inform_L[228][3];				l_cell_reg[226] = inform_L[225][3];				l_cell_reg[227] = inform_L[229][3];				l_cell_reg[228] = inform_L[226][3];				l_cell_reg[229] = inform_L[230][3];				l_cell_reg[230] = inform_L[227][3];				l_cell_reg[231] = inform_L[231][3];				l_cell_reg[232] = inform_L[232][3];				l_cell_reg[233] = inform_L[236][3];				l_cell_reg[234] = inform_L[233][3];				l_cell_reg[235] = inform_L[237][3];				l_cell_reg[236] = inform_L[234][3];				l_cell_reg[237] = inform_L[238][3];				l_cell_reg[238] = inform_L[235][3];				l_cell_reg[239] = inform_L[239][3];				l_cell_reg[240] = inform_L[240][3];				l_cell_reg[241] = inform_L[244][3];				l_cell_reg[242] = inform_L[241][3];				l_cell_reg[243] = inform_L[245][3];				l_cell_reg[244] = inform_L[242][3];				l_cell_reg[245] = inform_L[246][3];				l_cell_reg[246] = inform_L[243][3];				l_cell_reg[247] = inform_L[247][3];				l_cell_reg[248] = inform_L[248][3];				l_cell_reg[249] = inform_L[252][3];				l_cell_reg[250] = inform_L[249][3];				l_cell_reg[251] = inform_L[253][3];				l_cell_reg[252] = inform_L[250][3];				l_cell_reg[253] = inform_L[254][3];				l_cell_reg[254] = inform_L[251][3];				l_cell_reg[255] = inform_L[255][3];				l_cell_reg[256] = inform_L[256][3];				l_cell_reg[257] = inform_L[260][3];				l_cell_reg[258] = inform_L[257][3];				l_cell_reg[259] = inform_L[261][3];				l_cell_reg[260] = inform_L[258][3];				l_cell_reg[261] = inform_L[262][3];				l_cell_reg[262] = inform_L[259][3];				l_cell_reg[263] = inform_L[263][3];				l_cell_reg[264] = inform_L[264][3];				l_cell_reg[265] = inform_L[268][3];				l_cell_reg[266] = inform_L[265][3];				l_cell_reg[267] = inform_L[269][3];				l_cell_reg[268] = inform_L[266][3];				l_cell_reg[269] = inform_L[270][3];				l_cell_reg[270] = inform_L[267][3];				l_cell_reg[271] = inform_L[271][3];				l_cell_reg[272] = inform_L[272][3];				l_cell_reg[273] = inform_L[276][3];				l_cell_reg[274] = inform_L[273][3];				l_cell_reg[275] = inform_L[277][3];				l_cell_reg[276] = inform_L[274][3];				l_cell_reg[277] = inform_L[278][3];				l_cell_reg[278] = inform_L[275][3];				l_cell_reg[279] = inform_L[279][3];				l_cell_reg[280] = inform_L[280][3];				l_cell_reg[281] = inform_L[284][3];				l_cell_reg[282] = inform_L[281][3];				l_cell_reg[283] = inform_L[285][3];				l_cell_reg[284] = inform_L[282][3];				l_cell_reg[285] = inform_L[286][3];				l_cell_reg[286] = inform_L[283][3];				l_cell_reg[287] = inform_L[287][3];				l_cell_reg[288] = inform_L[288][3];				l_cell_reg[289] = inform_L[292][3];				l_cell_reg[290] = inform_L[289][3];				l_cell_reg[291] = inform_L[293][3];				l_cell_reg[292] = inform_L[290][3];				l_cell_reg[293] = inform_L[294][3];				l_cell_reg[294] = inform_L[291][3];				l_cell_reg[295] = inform_L[295][3];				l_cell_reg[296] = inform_L[296][3];				l_cell_reg[297] = inform_L[300][3];				l_cell_reg[298] = inform_L[297][3];				l_cell_reg[299] = inform_L[301][3];				l_cell_reg[300] = inform_L[298][3];				l_cell_reg[301] = inform_L[302][3];				l_cell_reg[302] = inform_L[299][3];				l_cell_reg[303] = inform_L[303][3];				l_cell_reg[304] = inform_L[304][3];				l_cell_reg[305] = inform_L[308][3];				l_cell_reg[306] = inform_L[305][3];				l_cell_reg[307] = inform_L[309][3];				l_cell_reg[308] = inform_L[306][3];				l_cell_reg[309] = inform_L[310][3];				l_cell_reg[310] = inform_L[307][3];				l_cell_reg[311] = inform_L[311][3];				l_cell_reg[312] = inform_L[312][3];				l_cell_reg[313] = inform_L[316][3];				l_cell_reg[314] = inform_L[313][3];				l_cell_reg[315] = inform_L[317][3];				l_cell_reg[316] = inform_L[314][3];				l_cell_reg[317] = inform_L[318][3];				l_cell_reg[318] = inform_L[315][3];				l_cell_reg[319] = inform_L[319][3];				l_cell_reg[320] = inform_L[320][3];				l_cell_reg[321] = inform_L[324][3];				l_cell_reg[322] = inform_L[321][3];				l_cell_reg[323] = inform_L[325][3];				l_cell_reg[324] = inform_L[322][3];				l_cell_reg[325] = inform_L[326][3];				l_cell_reg[326] = inform_L[323][3];				l_cell_reg[327] = inform_L[327][3];				l_cell_reg[328] = inform_L[328][3];				l_cell_reg[329] = inform_L[332][3];				l_cell_reg[330] = inform_L[329][3];				l_cell_reg[331] = inform_L[333][3];				l_cell_reg[332] = inform_L[330][3];				l_cell_reg[333] = inform_L[334][3];				l_cell_reg[334] = inform_L[331][3];				l_cell_reg[335] = inform_L[335][3];				l_cell_reg[336] = inform_L[336][3];				l_cell_reg[337] = inform_L[340][3];				l_cell_reg[338] = inform_L[337][3];				l_cell_reg[339] = inform_L[341][3];				l_cell_reg[340] = inform_L[338][3];				l_cell_reg[341] = inform_L[342][3];				l_cell_reg[342] = inform_L[339][3];				l_cell_reg[343] = inform_L[343][3];				l_cell_reg[344] = inform_L[344][3];				l_cell_reg[345] = inform_L[348][3];				l_cell_reg[346] = inform_L[345][3];				l_cell_reg[347] = inform_L[349][3];				l_cell_reg[348] = inform_L[346][3];				l_cell_reg[349] = inform_L[350][3];				l_cell_reg[350] = inform_L[347][3];				l_cell_reg[351] = inform_L[351][3];				l_cell_reg[352] = inform_L[352][3];				l_cell_reg[353] = inform_L[356][3];				l_cell_reg[354] = inform_L[353][3];				l_cell_reg[355] = inform_L[357][3];				l_cell_reg[356] = inform_L[354][3];				l_cell_reg[357] = inform_L[358][3];				l_cell_reg[358] = inform_L[355][3];				l_cell_reg[359] = inform_L[359][3];				l_cell_reg[360] = inform_L[360][3];				l_cell_reg[361] = inform_L[364][3];				l_cell_reg[362] = inform_L[361][3];				l_cell_reg[363] = inform_L[365][3];				l_cell_reg[364] = inform_L[362][3];				l_cell_reg[365] = inform_L[366][3];				l_cell_reg[366] = inform_L[363][3];				l_cell_reg[367] = inform_L[367][3];				l_cell_reg[368] = inform_L[368][3];				l_cell_reg[369] = inform_L[372][3];				l_cell_reg[370] = inform_L[369][3];				l_cell_reg[371] = inform_L[373][3];				l_cell_reg[372] = inform_L[370][3];				l_cell_reg[373] = inform_L[374][3];				l_cell_reg[374] = inform_L[371][3];				l_cell_reg[375] = inform_L[375][3];				l_cell_reg[376] = inform_L[376][3];				l_cell_reg[377] = inform_L[380][3];				l_cell_reg[378] = inform_L[377][3];				l_cell_reg[379] = inform_L[381][3];				l_cell_reg[380] = inform_L[378][3];				l_cell_reg[381] = inform_L[382][3];				l_cell_reg[382] = inform_L[379][3];				l_cell_reg[383] = inform_L[383][3];				l_cell_reg[384] = inform_L[384][3];				l_cell_reg[385] = inform_L[388][3];				l_cell_reg[386] = inform_L[385][3];				l_cell_reg[387] = inform_L[389][3];				l_cell_reg[388] = inform_L[386][3];				l_cell_reg[389] = inform_L[390][3];				l_cell_reg[390] = inform_L[387][3];				l_cell_reg[391] = inform_L[391][3];				l_cell_reg[392] = inform_L[392][3];				l_cell_reg[393] = inform_L[396][3];				l_cell_reg[394] = inform_L[393][3];				l_cell_reg[395] = inform_L[397][3];				l_cell_reg[396] = inform_L[394][3];				l_cell_reg[397] = inform_L[398][3];				l_cell_reg[398] = inform_L[395][3];				l_cell_reg[399] = inform_L[399][3];				l_cell_reg[400] = inform_L[400][3];				l_cell_reg[401] = inform_L[404][3];				l_cell_reg[402] = inform_L[401][3];				l_cell_reg[403] = inform_L[405][3];				l_cell_reg[404] = inform_L[402][3];				l_cell_reg[405] = inform_L[406][3];				l_cell_reg[406] = inform_L[403][3];				l_cell_reg[407] = inform_L[407][3];				l_cell_reg[408] = inform_L[408][3];				l_cell_reg[409] = inform_L[412][3];				l_cell_reg[410] = inform_L[409][3];				l_cell_reg[411] = inform_L[413][3];				l_cell_reg[412] = inform_L[410][3];				l_cell_reg[413] = inform_L[414][3];				l_cell_reg[414] = inform_L[411][3];				l_cell_reg[415] = inform_L[415][3];				l_cell_reg[416] = inform_L[416][3];				l_cell_reg[417] = inform_L[420][3];				l_cell_reg[418] = inform_L[417][3];				l_cell_reg[419] = inform_L[421][3];				l_cell_reg[420] = inform_L[418][3];				l_cell_reg[421] = inform_L[422][3];				l_cell_reg[422] = inform_L[419][3];				l_cell_reg[423] = inform_L[423][3];				l_cell_reg[424] = inform_L[424][3];				l_cell_reg[425] = inform_L[428][3];				l_cell_reg[426] = inform_L[425][3];				l_cell_reg[427] = inform_L[429][3];				l_cell_reg[428] = inform_L[426][3];				l_cell_reg[429] = inform_L[430][3];				l_cell_reg[430] = inform_L[427][3];				l_cell_reg[431] = inform_L[431][3];				l_cell_reg[432] = inform_L[432][3];				l_cell_reg[433] = inform_L[436][3];				l_cell_reg[434] = inform_L[433][3];				l_cell_reg[435] = inform_L[437][3];				l_cell_reg[436] = inform_L[434][3];				l_cell_reg[437] = inform_L[438][3];				l_cell_reg[438] = inform_L[435][3];				l_cell_reg[439] = inform_L[439][3];				l_cell_reg[440] = inform_L[440][3];				l_cell_reg[441] = inform_L[444][3];				l_cell_reg[442] = inform_L[441][3];				l_cell_reg[443] = inform_L[445][3];				l_cell_reg[444] = inform_L[442][3];				l_cell_reg[445] = inform_L[446][3];				l_cell_reg[446] = inform_L[443][3];				l_cell_reg[447] = inform_L[447][3];				l_cell_reg[448] = inform_L[448][3];				l_cell_reg[449] = inform_L[452][3];				l_cell_reg[450] = inform_L[449][3];				l_cell_reg[451] = inform_L[453][3];				l_cell_reg[452] = inform_L[450][3];				l_cell_reg[453] = inform_L[454][3];				l_cell_reg[454] = inform_L[451][3];				l_cell_reg[455] = inform_L[455][3];				l_cell_reg[456] = inform_L[456][3];				l_cell_reg[457] = inform_L[460][3];				l_cell_reg[458] = inform_L[457][3];				l_cell_reg[459] = inform_L[461][3];				l_cell_reg[460] = inform_L[458][3];				l_cell_reg[461] = inform_L[462][3];				l_cell_reg[462] = inform_L[459][3];				l_cell_reg[463] = inform_L[463][3];				l_cell_reg[464] = inform_L[464][3];				l_cell_reg[465] = inform_L[468][3];				l_cell_reg[466] = inform_L[465][3];				l_cell_reg[467] = inform_L[469][3];				l_cell_reg[468] = inform_L[466][3];				l_cell_reg[469] = inform_L[470][3];				l_cell_reg[470] = inform_L[467][3];				l_cell_reg[471] = inform_L[471][3];				l_cell_reg[472] = inform_L[472][3];				l_cell_reg[473] = inform_L[476][3];				l_cell_reg[474] = inform_L[473][3];				l_cell_reg[475] = inform_L[477][3];				l_cell_reg[476] = inform_L[474][3];				l_cell_reg[477] = inform_L[478][3];				l_cell_reg[478] = inform_L[475][3];				l_cell_reg[479] = inform_L[479][3];				l_cell_reg[480] = inform_L[480][3];				l_cell_reg[481] = inform_L[484][3];				l_cell_reg[482] = inform_L[481][3];				l_cell_reg[483] = inform_L[485][3];				l_cell_reg[484] = inform_L[482][3];				l_cell_reg[485] = inform_L[486][3];				l_cell_reg[486] = inform_L[483][3];				l_cell_reg[487] = inform_L[487][3];				l_cell_reg[488] = inform_L[488][3];				l_cell_reg[489] = inform_L[492][3];				l_cell_reg[490] = inform_L[489][3];				l_cell_reg[491] = inform_L[493][3];				l_cell_reg[492] = inform_L[490][3];				l_cell_reg[493] = inform_L[494][3];				l_cell_reg[494] = inform_L[491][3];				l_cell_reg[495] = inform_L[495][3];				l_cell_reg[496] = inform_L[496][3];				l_cell_reg[497] = inform_L[500][3];				l_cell_reg[498] = inform_L[497][3];				l_cell_reg[499] = inform_L[501][3];				l_cell_reg[500] = inform_L[498][3];				l_cell_reg[501] = inform_L[502][3];				l_cell_reg[502] = inform_L[499][3];				l_cell_reg[503] = inform_L[503][3];				l_cell_reg[504] = inform_L[504][3];				l_cell_reg[505] = inform_L[508][3];				l_cell_reg[506] = inform_L[505][3];				l_cell_reg[507] = inform_L[509][3];				l_cell_reg[508] = inform_L[506][3];				l_cell_reg[509] = inform_L[510][3];				l_cell_reg[510] = inform_L[507][3];				l_cell_reg[511] = inform_L[511][3];				l_cell_reg[512] = inform_L[512][3];				l_cell_reg[513] = inform_L[516][3];				l_cell_reg[514] = inform_L[513][3];				l_cell_reg[515] = inform_L[517][3];				l_cell_reg[516] = inform_L[514][3];				l_cell_reg[517] = inform_L[518][3];				l_cell_reg[518] = inform_L[515][3];				l_cell_reg[519] = inform_L[519][3];				l_cell_reg[520] = inform_L[520][3];				l_cell_reg[521] = inform_L[524][3];				l_cell_reg[522] = inform_L[521][3];				l_cell_reg[523] = inform_L[525][3];				l_cell_reg[524] = inform_L[522][3];				l_cell_reg[525] = inform_L[526][3];				l_cell_reg[526] = inform_L[523][3];				l_cell_reg[527] = inform_L[527][3];				l_cell_reg[528] = inform_L[528][3];				l_cell_reg[529] = inform_L[532][3];				l_cell_reg[530] = inform_L[529][3];				l_cell_reg[531] = inform_L[533][3];				l_cell_reg[532] = inform_L[530][3];				l_cell_reg[533] = inform_L[534][3];				l_cell_reg[534] = inform_L[531][3];				l_cell_reg[535] = inform_L[535][3];				l_cell_reg[536] = inform_L[536][3];				l_cell_reg[537] = inform_L[540][3];				l_cell_reg[538] = inform_L[537][3];				l_cell_reg[539] = inform_L[541][3];				l_cell_reg[540] = inform_L[538][3];				l_cell_reg[541] = inform_L[542][3];				l_cell_reg[542] = inform_L[539][3];				l_cell_reg[543] = inform_L[543][3];				l_cell_reg[544] = inform_L[544][3];				l_cell_reg[545] = inform_L[548][3];				l_cell_reg[546] = inform_L[545][3];				l_cell_reg[547] = inform_L[549][3];				l_cell_reg[548] = inform_L[546][3];				l_cell_reg[549] = inform_L[550][3];				l_cell_reg[550] = inform_L[547][3];				l_cell_reg[551] = inform_L[551][3];				l_cell_reg[552] = inform_L[552][3];				l_cell_reg[553] = inform_L[556][3];				l_cell_reg[554] = inform_L[553][3];				l_cell_reg[555] = inform_L[557][3];				l_cell_reg[556] = inform_L[554][3];				l_cell_reg[557] = inform_L[558][3];				l_cell_reg[558] = inform_L[555][3];				l_cell_reg[559] = inform_L[559][3];				l_cell_reg[560] = inform_L[560][3];				l_cell_reg[561] = inform_L[564][3];				l_cell_reg[562] = inform_L[561][3];				l_cell_reg[563] = inform_L[565][3];				l_cell_reg[564] = inform_L[562][3];				l_cell_reg[565] = inform_L[566][3];				l_cell_reg[566] = inform_L[563][3];				l_cell_reg[567] = inform_L[567][3];				l_cell_reg[568] = inform_L[568][3];				l_cell_reg[569] = inform_L[572][3];				l_cell_reg[570] = inform_L[569][3];				l_cell_reg[571] = inform_L[573][3];				l_cell_reg[572] = inform_L[570][3];				l_cell_reg[573] = inform_L[574][3];				l_cell_reg[574] = inform_L[571][3];				l_cell_reg[575] = inform_L[575][3];				l_cell_reg[576] = inform_L[576][3];				l_cell_reg[577] = inform_L[580][3];				l_cell_reg[578] = inform_L[577][3];				l_cell_reg[579] = inform_L[581][3];				l_cell_reg[580] = inform_L[578][3];				l_cell_reg[581] = inform_L[582][3];				l_cell_reg[582] = inform_L[579][3];				l_cell_reg[583] = inform_L[583][3];				l_cell_reg[584] = inform_L[584][3];				l_cell_reg[585] = inform_L[588][3];				l_cell_reg[586] = inform_L[585][3];				l_cell_reg[587] = inform_L[589][3];				l_cell_reg[588] = inform_L[586][3];				l_cell_reg[589] = inform_L[590][3];				l_cell_reg[590] = inform_L[587][3];				l_cell_reg[591] = inform_L[591][3];				l_cell_reg[592] = inform_L[592][3];				l_cell_reg[593] = inform_L[596][3];				l_cell_reg[594] = inform_L[593][3];				l_cell_reg[595] = inform_L[597][3];				l_cell_reg[596] = inform_L[594][3];				l_cell_reg[597] = inform_L[598][3];				l_cell_reg[598] = inform_L[595][3];				l_cell_reg[599] = inform_L[599][3];				l_cell_reg[600] = inform_L[600][3];				l_cell_reg[601] = inform_L[604][3];				l_cell_reg[602] = inform_L[601][3];				l_cell_reg[603] = inform_L[605][3];				l_cell_reg[604] = inform_L[602][3];				l_cell_reg[605] = inform_L[606][3];				l_cell_reg[606] = inform_L[603][3];				l_cell_reg[607] = inform_L[607][3];				l_cell_reg[608] = inform_L[608][3];				l_cell_reg[609] = inform_L[612][3];				l_cell_reg[610] = inform_L[609][3];				l_cell_reg[611] = inform_L[613][3];				l_cell_reg[612] = inform_L[610][3];				l_cell_reg[613] = inform_L[614][3];				l_cell_reg[614] = inform_L[611][3];				l_cell_reg[615] = inform_L[615][3];				l_cell_reg[616] = inform_L[616][3];				l_cell_reg[617] = inform_L[620][3];				l_cell_reg[618] = inform_L[617][3];				l_cell_reg[619] = inform_L[621][3];				l_cell_reg[620] = inform_L[618][3];				l_cell_reg[621] = inform_L[622][3];				l_cell_reg[622] = inform_L[619][3];				l_cell_reg[623] = inform_L[623][3];				l_cell_reg[624] = inform_L[624][3];				l_cell_reg[625] = inform_L[628][3];				l_cell_reg[626] = inform_L[625][3];				l_cell_reg[627] = inform_L[629][3];				l_cell_reg[628] = inform_L[626][3];				l_cell_reg[629] = inform_L[630][3];				l_cell_reg[630] = inform_L[627][3];				l_cell_reg[631] = inform_L[631][3];				l_cell_reg[632] = inform_L[632][3];				l_cell_reg[633] = inform_L[636][3];				l_cell_reg[634] = inform_L[633][3];				l_cell_reg[635] = inform_L[637][3];				l_cell_reg[636] = inform_L[634][3];				l_cell_reg[637] = inform_L[638][3];				l_cell_reg[638] = inform_L[635][3];				l_cell_reg[639] = inform_L[639][3];				l_cell_reg[640] = inform_L[640][3];				l_cell_reg[641] = inform_L[644][3];				l_cell_reg[642] = inform_L[641][3];				l_cell_reg[643] = inform_L[645][3];				l_cell_reg[644] = inform_L[642][3];				l_cell_reg[645] = inform_L[646][3];				l_cell_reg[646] = inform_L[643][3];				l_cell_reg[647] = inform_L[647][3];				l_cell_reg[648] = inform_L[648][3];				l_cell_reg[649] = inform_L[652][3];				l_cell_reg[650] = inform_L[649][3];				l_cell_reg[651] = inform_L[653][3];				l_cell_reg[652] = inform_L[650][3];				l_cell_reg[653] = inform_L[654][3];				l_cell_reg[654] = inform_L[651][3];				l_cell_reg[655] = inform_L[655][3];				l_cell_reg[656] = inform_L[656][3];				l_cell_reg[657] = inform_L[660][3];				l_cell_reg[658] = inform_L[657][3];				l_cell_reg[659] = inform_L[661][3];				l_cell_reg[660] = inform_L[658][3];				l_cell_reg[661] = inform_L[662][3];				l_cell_reg[662] = inform_L[659][3];				l_cell_reg[663] = inform_L[663][3];				l_cell_reg[664] = inform_L[664][3];				l_cell_reg[665] = inform_L[668][3];				l_cell_reg[666] = inform_L[665][3];				l_cell_reg[667] = inform_L[669][3];				l_cell_reg[668] = inform_L[666][3];				l_cell_reg[669] = inform_L[670][3];				l_cell_reg[670] = inform_L[667][3];				l_cell_reg[671] = inform_L[671][3];				l_cell_reg[672] = inform_L[672][3];				l_cell_reg[673] = inform_L[676][3];				l_cell_reg[674] = inform_L[673][3];				l_cell_reg[675] = inform_L[677][3];				l_cell_reg[676] = inform_L[674][3];				l_cell_reg[677] = inform_L[678][3];				l_cell_reg[678] = inform_L[675][3];				l_cell_reg[679] = inform_L[679][3];				l_cell_reg[680] = inform_L[680][3];				l_cell_reg[681] = inform_L[684][3];				l_cell_reg[682] = inform_L[681][3];				l_cell_reg[683] = inform_L[685][3];				l_cell_reg[684] = inform_L[682][3];				l_cell_reg[685] = inform_L[686][3];				l_cell_reg[686] = inform_L[683][3];				l_cell_reg[687] = inform_L[687][3];				l_cell_reg[688] = inform_L[688][3];				l_cell_reg[689] = inform_L[692][3];				l_cell_reg[690] = inform_L[689][3];				l_cell_reg[691] = inform_L[693][3];				l_cell_reg[692] = inform_L[690][3];				l_cell_reg[693] = inform_L[694][3];				l_cell_reg[694] = inform_L[691][3];				l_cell_reg[695] = inform_L[695][3];				l_cell_reg[696] = inform_L[696][3];				l_cell_reg[697] = inform_L[700][3];				l_cell_reg[698] = inform_L[697][3];				l_cell_reg[699] = inform_L[701][3];				l_cell_reg[700] = inform_L[698][3];				l_cell_reg[701] = inform_L[702][3];				l_cell_reg[702] = inform_L[699][3];				l_cell_reg[703] = inform_L[703][3];				l_cell_reg[704] = inform_L[704][3];				l_cell_reg[705] = inform_L[708][3];				l_cell_reg[706] = inform_L[705][3];				l_cell_reg[707] = inform_L[709][3];				l_cell_reg[708] = inform_L[706][3];				l_cell_reg[709] = inform_L[710][3];				l_cell_reg[710] = inform_L[707][3];				l_cell_reg[711] = inform_L[711][3];				l_cell_reg[712] = inform_L[712][3];				l_cell_reg[713] = inform_L[716][3];				l_cell_reg[714] = inform_L[713][3];				l_cell_reg[715] = inform_L[717][3];				l_cell_reg[716] = inform_L[714][3];				l_cell_reg[717] = inform_L[718][3];				l_cell_reg[718] = inform_L[715][3];				l_cell_reg[719] = inform_L[719][3];				l_cell_reg[720] = inform_L[720][3];				l_cell_reg[721] = inform_L[724][3];				l_cell_reg[722] = inform_L[721][3];				l_cell_reg[723] = inform_L[725][3];				l_cell_reg[724] = inform_L[722][3];				l_cell_reg[725] = inform_L[726][3];				l_cell_reg[726] = inform_L[723][3];				l_cell_reg[727] = inform_L[727][3];				l_cell_reg[728] = inform_L[728][3];				l_cell_reg[729] = inform_L[732][3];				l_cell_reg[730] = inform_L[729][3];				l_cell_reg[731] = inform_L[733][3];				l_cell_reg[732] = inform_L[730][3];				l_cell_reg[733] = inform_L[734][3];				l_cell_reg[734] = inform_L[731][3];				l_cell_reg[735] = inform_L[735][3];				l_cell_reg[736] = inform_L[736][3];				l_cell_reg[737] = inform_L[740][3];				l_cell_reg[738] = inform_L[737][3];				l_cell_reg[739] = inform_L[741][3];				l_cell_reg[740] = inform_L[738][3];				l_cell_reg[741] = inform_L[742][3];				l_cell_reg[742] = inform_L[739][3];				l_cell_reg[743] = inform_L[743][3];				l_cell_reg[744] = inform_L[744][3];				l_cell_reg[745] = inform_L[748][3];				l_cell_reg[746] = inform_L[745][3];				l_cell_reg[747] = inform_L[749][3];				l_cell_reg[748] = inform_L[746][3];				l_cell_reg[749] = inform_L[750][3];				l_cell_reg[750] = inform_L[747][3];				l_cell_reg[751] = inform_L[751][3];				l_cell_reg[752] = inform_L[752][3];				l_cell_reg[753] = inform_L[756][3];				l_cell_reg[754] = inform_L[753][3];				l_cell_reg[755] = inform_L[757][3];				l_cell_reg[756] = inform_L[754][3];				l_cell_reg[757] = inform_L[758][3];				l_cell_reg[758] = inform_L[755][3];				l_cell_reg[759] = inform_L[759][3];				l_cell_reg[760] = inform_L[760][3];				l_cell_reg[761] = inform_L[764][3];				l_cell_reg[762] = inform_L[761][3];				l_cell_reg[763] = inform_L[765][3];				l_cell_reg[764] = inform_L[762][3];				l_cell_reg[765] = inform_L[766][3];				l_cell_reg[766] = inform_L[763][3];				l_cell_reg[767] = inform_L[767][3];				l_cell_reg[768] = inform_L[768][3];				l_cell_reg[769] = inform_L[772][3];				l_cell_reg[770] = inform_L[769][3];				l_cell_reg[771] = inform_L[773][3];				l_cell_reg[772] = inform_L[770][3];				l_cell_reg[773] = inform_L[774][3];				l_cell_reg[774] = inform_L[771][3];				l_cell_reg[775] = inform_L[775][3];				l_cell_reg[776] = inform_L[776][3];				l_cell_reg[777] = inform_L[780][3];				l_cell_reg[778] = inform_L[777][3];				l_cell_reg[779] = inform_L[781][3];				l_cell_reg[780] = inform_L[778][3];				l_cell_reg[781] = inform_L[782][3];				l_cell_reg[782] = inform_L[779][3];				l_cell_reg[783] = inform_L[783][3];				l_cell_reg[784] = inform_L[784][3];				l_cell_reg[785] = inform_L[788][3];				l_cell_reg[786] = inform_L[785][3];				l_cell_reg[787] = inform_L[789][3];				l_cell_reg[788] = inform_L[786][3];				l_cell_reg[789] = inform_L[790][3];				l_cell_reg[790] = inform_L[787][3];				l_cell_reg[791] = inform_L[791][3];				l_cell_reg[792] = inform_L[792][3];				l_cell_reg[793] = inform_L[796][3];				l_cell_reg[794] = inform_L[793][3];				l_cell_reg[795] = inform_L[797][3];				l_cell_reg[796] = inform_L[794][3];				l_cell_reg[797] = inform_L[798][3];				l_cell_reg[798] = inform_L[795][3];				l_cell_reg[799] = inform_L[799][3];				l_cell_reg[800] = inform_L[800][3];				l_cell_reg[801] = inform_L[804][3];				l_cell_reg[802] = inform_L[801][3];				l_cell_reg[803] = inform_L[805][3];				l_cell_reg[804] = inform_L[802][3];				l_cell_reg[805] = inform_L[806][3];				l_cell_reg[806] = inform_L[803][3];				l_cell_reg[807] = inform_L[807][3];				l_cell_reg[808] = inform_L[808][3];				l_cell_reg[809] = inform_L[812][3];				l_cell_reg[810] = inform_L[809][3];				l_cell_reg[811] = inform_L[813][3];				l_cell_reg[812] = inform_L[810][3];				l_cell_reg[813] = inform_L[814][3];				l_cell_reg[814] = inform_L[811][3];				l_cell_reg[815] = inform_L[815][3];				l_cell_reg[816] = inform_L[816][3];				l_cell_reg[817] = inform_L[820][3];				l_cell_reg[818] = inform_L[817][3];				l_cell_reg[819] = inform_L[821][3];				l_cell_reg[820] = inform_L[818][3];				l_cell_reg[821] = inform_L[822][3];				l_cell_reg[822] = inform_L[819][3];				l_cell_reg[823] = inform_L[823][3];				l_cell_reg[824] = inform_L[824][3];				l_cell_reg[825] = inform_L[828][3];				l_cell_reg[826] = inform_L[825][3];				l_cell_reg[827] = inform_L[829][3];				l_cell_reg[828] = inform_L[826][3];				l_cell_reg[829] = inform_L[830][3];				l_cell_reg[830] = inform_L[827][3];				l_cell_reg[831] = inform_L[831][3];				l_cell_reg[832] = inform_L[832][3];				l_cell_reg[833] = inform_L[836][3];				l_cell_reg[834] = inform_L[833][3];				l_cell_reg[835] = inform_L[837][3];				l_cell_reg[836] = inform_L[834][3];				l_cell_reg[837] = inform_L[838][3];				l_cell_reg[838] = inform_L[835][3];				l_cell_reg[839] = inform_L[839][3];				l_cell_reg[840] = inform_L[840][3];				l_cell_reg[841] = inform_L[844][3];				l_cell_reg[842] = inform_L[841][3];				l_cell_reg[843] = inform_L[845][3];				l_cell_reg[844] = inform_L[842][3];				l_cell_reg[845] = inform_L[846][3];				l_cell_reg[846] = inform_L[843][3];				l_cell_reg[847] = inform_L[847][3];				l_cell_reg[848] = inform_L[848][3];				l_cell_reg[849] = inform_L[852][3];				l_cell_reg[850] = inform_L[849][3];				l_cell_reg[851] = inform_L[853][3];				l_cell_reg[852] = inform_L[850][3];				l_cell_reg[853] = inform_L[854][3];				l_cell_reg[854] = inform_L[851][3];				l_cell_reg[855] = inform_L[855][3];				l_cell_reg[856] = inform_L[856][3];				l_cell_reg[857] = inform_L[860][3];				l_cell_reg[858] = inform_L[857][3];				l_cell_reg[859] = inform_L[861][3];				l_cell_reg[860] = inform_L[858][3];				l_cell_reg[861] = inform_L[862][3];				l_cell_reg[862] = inform_L[859][3];				l_cell_reg[863] = inform_L[863][3];				l_cell_reg[864] = inform_L[864][3];				l_cell_reg[865] = inform_L[868][3];				l_cell_reg[866] = inform_L[865][3];				l_cell_reg[867] = inform_L[869][3];				l_cell_reg[868] = inform_L[866][3];				l_cell_reg[869] = inform_L[870][3];				l_cell_reg[870] = inform_L[867][3];				l_cell_reg[871] = inform_L[871][3];				l_cell_reg[872] = inform_L[872][3];				l_cell_reg[873] = inform_L[876][3];				l_cell_reg[874] = inform_L[873][3];				l_cell_reg[875] = inform_L[877][3];				l_cell_reg[876] = inform_L[874][3];				l_cell_reg[877] = inform_L[878][3];				l_cell_reg[878] = inform_L[875][3];				l_cell_reg[879] = inform_L[879][3];				l_cell_reg[880] = inform_L[880][3];				l_cell_reg[881] = inform_L[884][3];				l_cell_reg[882] = inform_L[881][3];				l_cell_reg[883] = inform_L[885][3];				l_cell_reg[884] = inform_L[882][3];				l_cell_reg[885] = inform_L[886][3];				l_cell_reg[886] = inform_L[883][3];				l_cell_reg[887] = inform_L[887][3];				l_cell_reg[888] = inform_L[888][3];				l_cell_reg[889] = inform_L[892][3];				l_cell_reg[890] = inform_L[889][3];				l_cell_reg[891] = inform_L[893][3];				l_cell_reg[892] = inform_L[890][3];				l_cell_reg[893] = inform_L[894][3];				l_cell_reg[894] = inform_L[891][3];				l_cell_reg[895] = inform_L[895][3];				l_cell_reg[896] = inform_L[896][3];				l_cell_reg[897] = inform_L[900][3];				l_cell_reg[898] = inform_L[897][3];				l_cell_reg[899] = inform_L[901][3];				l_cell_reg[900] = inform_L[898][3];				l_cell_reg[901] = inform_L[902][3];				l_cell_reg[902] = inform_L[899][3];				l_cell_reg[903] = inform_L[903][3];				l_cell_reg[904] = inform_L[904][3];				l_cell_reg[905] = inform_L[908][3];				l_cell_reg[906] = inform_L[905][3];				l_cell_reg[907] = inform_L[909][3];				l_cell_reg[908] = inform_L[906][3];				l_cell_reg[909] = inform_L[910][3];				l_cell_reg[910] = inform_L[907][3];				l_cell_reg[911] = inform_L[911][3];				l_cell_reg[912] = inform_L[912][3];				l_cell_reg[913] = inform_L[916][3];				l_cell_reg[914] = inform_L[913][3];				l_cell_reg[915] = inform_L[917][3];				l_cell_reg[916] = inform_L[914][3];				l_cell_reg[917] = inform_L[918][3];				l_cell_reg[918] = inform_L[915][3];				l_cell_reg[919] = inform_L[919][3];				l_cell_reg[920] = inform_L[920][3];				l_cell_reg[921] = inform_L[924][3];				l_cell_reg[922] = inform_L[921][3];				l_cell_reg[923] = inform_L[925][3];				l_cell_reg[924] = inform_L[922][3];				l_cell_reg[925] = inform_L[926][3];				l_cell_reg[926] = inform_L[923][3];				l_cell_reg[927] = inform_L[927][3];				l_cell_reg[928] = inform_L[928][3];				l_cell_reg[929] = inform_L[932][3];				l_cell_reg[930] = inform_L[929][3];				l_cell_reg[931] = inform_L[933][3];				l_cell_reg[932] = inform_L[930][3];				l_cell_reg[933] = inform_L[934][3];				l_cell_reg[934] = inform_L[931][3];				l_cell_reg[935] = inform_L[935][3];				l_cell_reg[936] = inform_L[936][3];				l_cell_reg[937] = inform_L[940][3];				l_cell_reg[938] = inform_L[937][3];				l_cell_reg[939] = inform_L[941][3];				l_cell_reg[940] = inform_L[938][3];				l_cell_reg[941] = inform_L[942][3];				l_cell_reg[942] = inform_L[939][3];				l_cell_reg[943] = inform_L[943][3];				l_cell_reg[944] = inform_L[944][3];				l_cell_reg[945] = inform_L[948][3];				l_cell_reg[946] = inform_L[945][3];				l_cell_reg[947] = inform_L[949][3];				l_cell_reg[948] = inform_L[946][3];				l_cell_reg[949] = inform_L[950][3];				l_cell_reg[950] = inform_L[947][3];				l_cell_reg[951] = inform_L[951][3];				l_cell_reg[952] = inform_L[952][3];				l_cell_reg[953] = inform_L[956][3];				l_cell_reg[954] = inform_L[953][3];				l_cell_reg[955] = inform_L[957][3];				l_cell_reg[956] = inform_L[954][3];				l_cell_reg[957] = inform_L[958][3];				l_cell_reg[958] = inform_L[955][3];				l_cell_reg[959] = inform_L[959][3];				l_cell_reg[960] = inform_L[960][3];				l_cell_reg[961] = inform_L[964][3];				l_cell_reg[962] = inform_L[961][3];				l_cell_reg[963] = inform_L[965][3];				l_cell_reg[964] = inform_L[962][3];				l_cell_reg[965] = inform_L[966][3];				l_cell_reg[966] = inform_L[963][3];				l_cell_reg[967] = inform_L[967][3];				l_cell_reg[968] = inform_L[968][3];				l_cell_reg[969] = inform_L[972][3];				l_cell_reg[970] = inform_L[969][3];				l_cell_reg[971] = inform_L[973][3];				l_cell_reg[972] = inform_L[970][3];				l_cell_reg[973] = inform_L[974][3];				l_cell_reg[974] = inform_L[971][3];				l_cell_reg[975] = inform_L[975][3];				l_cell_reg[976] = inform_L[976][3];				l_cell_reg[977] = inform_L[980][3];				l_cell_reg[978] = inform_L[977][3];				l_cell_reg[979] = inform_L[981][3];				l_cell_reg[980] = inform_L[978][3];				l_cell_reg[981] = inform_L[982][3];				l_cell_reg[982] = inform_L[979][3];				l_cell_reg[983] = inform_L[983][3];				l_cell_reg[984] = inform_L[984][3];				l_cell_reg[985] = inform_L[988][3];				l_cell_reg[986] = inform_L[985][3];				l_cell_reg[987] = inform_L[989][3];				l_cell_reg[988] = inform_L[986][3];				l_cell_reg[989] = inform_L[990][3];				l_cell_reg[990] = inform_L[987][3];				l_cell_reg[991] = inform_L[991][3];				l_cell_reg[992] = inform_L[992][3];				l_cell_reg[993] = inform_L[996][3];				l_cell_reg[994] = inform_L[993][3];				l_cell_reg[995] = inform_L[997][3];				l_cell_reg[996] = inform_L[994][3];				l_cell_reg[997] = inform_L[998][3];				l_cell_reg[998] = inform_L[995][3];				l_cell_reg[999] = inform_L[999][3];				l_cell_reg[1000] = inform_L[1000][3];				l_cell_reg[1001] = inform_L[1004][3];				l_cell_reg[1002] = inform_L[1001][3];				l_cell_reg[1003] = inform_L[1005][3];				l_cell_reg[1004] = inform_L[1002][3];				l_cell_reg[1005] = inform_L[1006][3];				l_cell_reg[1006] = inform_L[1003][3];				l_cell_reg[1007] = inform_L[1007][3];				l_cell_reg[1008] = inform_L[1008][3];				l_cell_reg[1009] = inform_L[1012][3];				l_cell_reg[1010] = inform_L[1009][3];				l_cell_reg[1011] = inform_L[1013][3];				l_cell_reg[1012] = inform_L[1010][3];				l_cell_reg[1013] = inform_L[1014][3];				l_cell_reg[1014] = inform_L[1011][3];				l_cell_reg[1015] = inform_L[1015][3];				l_cell_reg[1016] = inform_L[1016][3];				l_cell_reg[1017] = inform_L[1020][3];				l_cell_reg[1018] = inform_L[1017][3];				l_cell_reg[1019] = inform_L[1021][3];				l_cell_reg[1020] = inform_L[1018][3];				l_cell_reg[1021] = inform_L[1022][3];				l_cell_reg[1022] = inform_L[1019][3];				l_cell_reg[1023] = inform_L[1023][3];			end
			4:			begin				r_cell_reg[0] = inform_R[0][3];				r_cell_reg[1] = inform_R[8][3];				r_cell_reg[2] = inform_R[1][3];				r_cell_reg[3] = inform_R[9][3];				r_cell_reg[4] = inform_R[2][3];				r_cell_reg[5] = inform_R[10][3];				r_cell_reg[6] = inform_R[3][3];				r_cell_reg[7] = inform_R[11][3];				r_cell_reg[8] = inform_R[4][3];				r_cell_reg[9] = inform_R[12][3];				r_cell_reg[10] = inform_R[5][3];				r_cell_reg[11] = inform_R[13][3];				r_cell_reg[12] = inform_R[6][3];				r_cell_reg[13] = inform_R[14][3];				r_cell_reg[14] = inform_R[7][3];				r_cell_reg[15] = inform_R[15][3];				r_cell_reg[16] = inform_R[16][3];				r_cell_reg[17] = inform_R[24][3];				r_cell_reg[18] = inform_R[17][3];				r_cell_reg[19] = inform_R[25][3];				r_cell_reg[20] = inform_R[18][3];				r_cell_reg[21] = inform_R[26][3];				r_cell_reg[22] = inform_R[19][3];				r_cell_reg[23] = inform_R[27][3];				r_cell_reg[24] = inform_R[20][3];				r_cell_reg[25] = inform_R[28][3];				r_cell_reg[26] = inform_R[21][3];				r_cell_reg[27] = inform_R[29][3];				r_cell_reg[28] = inform_R[22][3];				r_cell_reg[29] = inform_R[30][3];				r_cell_reg[30] = inform_R[23][3];				r_cell_reg[31] = inform_R[31][3];				r_cell_reg[32] = inform_R[32][3];				r_cell_reg[33] = inform_R[40][3];				r_cell_reg[34] = inform_R[33][3];				r_cell_reg[35] = inform_R[41][3];				r_cell_reg[36] = inform_R[34][3];				r_cell_reg[37] = inform_R[42][3];				r_cell_reg[38] = inform_R[35][3];				r_cell_reg[39] = inform_R[43][3];				r_cell_reg[40] = inform_R[36][3];				r_cell_reg[41] = inform_R[44][3];				r_cell_reg[42] = inform_R[37][3];				r_cell_reg[43] = inform_R[45][3];				r_cell_reg[44] = inform_R[38][3];				r_cell_reg[45] = inform_R[46][3];				r_cell_reg[46] = inform_R[39][3];				r_cell_reg[47] = inform_R[47][3];				r_cell_reg[48] = inform_R[48][3];				r_cell_reg[49] = inform_R[56][3];				r_cell_reg[50] = inform_R[49][3];				r_cell_reg[51] = inform_R[57][3];				r_cell_reg[52] = inform_R[50][3];				r_cell_reg[53] = inform_R[58][3];				r_cell_reg[54] = inform_R[51][3];				r_cell_reg[55] = inform_R[59][3];				r_cell_reg[56] = inform_R[52][3];				r_cell_reg[57] = inform_R[60][3];				r_cell_reg[58] = inform_R[53][3];				r_cell_reg[59] = inform_R[61][3];				r_cell_reg[60] = inform_R[54][3];				r_cell_reg[61] = inform_R[62][3];				r_cell_reg[62] = inform_R[55][3];				r_cell_reg[63] = inform_R[63][3];				r_cell_reg[64] = inform_R[64][3];				r_cell_reg[65] = inform_R[72][3];				r_cell_reg[66] = inform_R[65][3];				r_cell_reg[67] = inform_R[73][3];				r_cell_reg[68] = inform_R[66][3];				r_cell_reg[69] = inform_R[74][3];				r_cell_reg[70] = inform_R[67][3];				r_cell_reg[71] = inform_R[75][3];				r_cell_reg[72] = inform_R[68][3];				r_cell_reg[73] = inform_R[76][3];				r_cell_reg[74] = inform_R[69][3];				r_cell_reg[75] = inform_R[77][3];				r_cell_reg[76] = inform_R[70][3];				r_cell_reg[77] = inform_R[78][3];				r_cell_reg[78] = inform_R[71][3];				r_cell_reg[79] = inform_R[79][3];				r_cell_reg[80] = inform_R[80][3];				r_cell_reg[81] = inform_R[88][3];				r_cell_reg[82] = inform_R[81][3];				r_cell_reg[83] = inform_R[89][3];				r_cell_reg[84] = inform_R[82][3];				r_cell_reg[85] = inform_R[90][3];				r_cell_reg[86] = inform_R[83][3];				r_cell_reg[87] = inform_R[91][3];				r_cell_reg[88] = inform_R[84][3];				r_cell_reg[89] = inform_R[92][3];				r_cell_reg[90] = inform_R[85][3];				r_cell_reg[91] = inform_R[93][3];				r_cell_reg[92] = inform_R[86][3];				r_cell_reg[93] = inform_R[94][3];				r_cell_reg[94] = inform_R[87][3];				r_cell_reg[95] = inform_R[95][3];				r_cell_reg[96] = inform_R[96][3];				r_cell_reg[97] = inform_R[104][3];				r_cell_reg[98] = inform_R[97][3];				r_cell_reg[99] = inform_R[105][3];				r_cell_reg[100] = inform_R[98][3];				r_cell_reg[101] = inform_R[106][3];				r_cell_reg[102] = inform_R[99][3];				r_cell_reg[103] = inform_R[107][3];				r_cell_reg[104] = inform_R[100][3];				r_cell_reg[105] = inform_R[108][3];				r_cell_reg[106] = inform_R[101][3];				r_cell_reg[107] = inform_R[109][3];				r_cell_reg[108] = inform_R[102][3];				r_cell_reg[109] = inform_R[110][3];				r_cell_reg[110] = inform_R[103][3];				r_cell_reg[111] = inform_R[111][3];				r_cell_reg[112] = inform_R[112][3];				r_cell_reg[113] = inform_R[120][3];				r_cell_reg[114] = inform_R[113][3];				r_cell_reg[115] = inform_R[121][3];				r_cell_reg[116] = inform_R[114][3];				r_cell_reg[117] = inform_R[122][3];				r_cell_reg[118] = inform_R[115][3];				r_cell_reg[119] = inform_R[123][3];				r_cell_reg[120] = inform_R[116][3];				r_cell_reg[121] = inform_R[124][3];				r_cell_reg[122] = inform_R[117][3];				r_cell_reg[123] = inform_R[125][3];				r_cell_reg[124] = inform_R[118][3];				r_cell_reg[125] = inform_R[126][3];				r_cell_reg[126] = inform_R[119][3];				r_cell_reg[127] = inform_R[127][3];				r_cell_reg[128] = inform_R[128][3];				r_cell_reg[129] = inform_R[136][3];				r_cell_reg[130] = inform_R[129][3];				r_cell_reg[131] = inform_R[137][3];				r_cell_reg[132] = inform_R[130][3];				r_cell_reg[133] = inform_R[138][3];				r_cell_reg[134] = inform_R[131][3];				r_cell_reg[135] = inform_R[139][3];				r_cell_reg[136] = inform_R[132][3];				r_cell_reg[137] = inform_R[140][3];				r_cell_reg[138] = inform_R[133][3];				r_cell_reg[139] = inform_R[141][3];				r_cell_reg[140] = inform_R[134][3];				r_cell_reg[141] = inform_R[142][3];				r_cell_reg[142] = inform_R[135][3];				r_cell_reg[143] = inform_R[143][3];				r_cell_reg[144] = inform_R[144][3];				r_cell_reg[145] = inform_R[152][3];				r_cell_reg[146] = inform_R[145][3];				r_cell_reg[147] = inform_R[153][3];				r_cell_reg[148] = inform_R[146][3];				r_cell_reg[149] = inform_R[154][3];				r_cell_reg[150] = inform_R[147][3];				r_cell_reg[151] = inform_R[155][3];				r_cell_reg[152] = inform_R[148][3];				r_cell_reg[153] = inform_R[156][3];				r_cell_reg[154] = inform_R[149][3];				r_cell_reg[155] = inform_R[157][3];				r_cell_reg[156] = inform_R[150][3];				r_cell_reg[157] = inform_R[158][3];				r_cell_reg[158] = inform_R[151][3];				r_cell_reg[159] = inform_R[159][3];				r_cell_reg[160] = inform_R[160][3];				r_cell_reg[161] = inform_R[168][3];				r_cell_reg[162] = inform_R[161][3];				r_cell_reg[163] = inform_R[169][3];				r_cell_reg[164] = inform_R[162][3];				r_cell_reg[165] = inform_R[170][3];				r_cell_reg[166] = inform_R[163][3];				r_cell_reg[167] = inform_R[171][3];				r_cell_reg[168] = inform_R[164][3];				r_cell_reg[169] = inform_R[172][3];				r_cell_reg[170] = inform_R[165][3];				r_cell_reg[171] = inform_R[173][3];				r_cell_reg[172] = inform_R[166][3];				r_cell_reg[173] = inform_R[174][3];				r_cell_reg[174] = inform_R[167][3];				r_cell_reg[175] = inform_R[175][3];				r_cell_reg[176] = inform_R[176][3];				r_cell_reg[177] = inform_R[184][3];				r_cell_reg[178] = inform_R[177][3];				r_cell_reg[179] = inform_R[185][3];				r_cell_reg[180] = inform_R[178][3];				r_cell_reg[181] = inform_R[186][3];				r_cell_reg[182] = inform_R[179][3];				r_cell_reg[183] = inform_R[187][3];				r_cell_reg[184] = inform_R[180][3];				r_cell_reg[185] = inform_R[188][3];				r_cell_reg[186] = inform_R[181][3];				r_cell_reg[187] = inform_R[189][3];				r_cell_reg[188] = inform_R[182][3];				r_cell_reg[189] = inform_R[190][3];				r_cell_reg[190] = inform_R[183][3];				r_cell_reg[191] = inform_R[191][3];				r_cell_reg[192] = inform_R[192][3];				r_cell_reg[193] = inform_R[200][3];				r_cell_reg[194] = inform_R[193][3];				r_cell_reg[195] = inform_R[201][3];				r_cell_reg[196] = inform_R[194][3];				r_cell_reg[197] = inform_R[202][3];				r_cell_reg[198] = inform_R[195][3];				r_cell_reg[199] = inform_R[203][3];				r_cell_reg[200] = inform_R[196][3];				r_cell_reg[201] = inform_R[204][3];				r_cell_reg[202] = inform_R[197][3];				r_cell_reg[203] = inform_R[205][3];				r_cell_reg[204] = inform_R[198][3];				r_cell_reg[205] = inform_R[206][3];				r_cell_reg[206] = inform_R[199][3];				r_cell_reg[207] = inform_R[207][3];				r_cell_reg[208] = inform_R[208][3];				r_cell_reg[209] = inform_R[216][3];				r_cell_reg[210] = inform_R[209][3];				r_cell_reg[211] = inform_R[217][3];				r_cell_reg[212] = inform_R[210][3];				r_cell_reg[213] = inform_R[218][3];				r_cell_reg[214] = inform_R[211][3];				r_cell_reg[215] = inform_R[219][3];				r_cell_reg[216] = inform_R[212][3];				r_cell_reg[217] = inform_R[220][3];				r_cell_reg[218] = inform_R[213][3];				r_cell_reg[219] = inform_R[221][3];				r_cell_reg[220] = inform_R[214][3];				r_cell_reg[221] = inform_R[222][3];				r_cell_reg[222] = inform_R[215][3];				r_cell_reg[223] = inform_R[223][3];				r_cell_reg[224] = inform_R[224][3];				r_cell_reg[225] = inform_R[232][3];				r_cell_reg[226] = inform_R[225][3];				r_cell_reg[227] = inform_R[233][3];				r_cell_reg[228] = inform_R[226][3];				r_cell_reg[229] = inform_R[234][3];				r_cell_reg[230] = inform_R[227][3];				r_cell_reg[231] = inform_R[235][3];				r_cell_reg[232] = inform_R[228][3];				r_cell_reg[233] = inform_R[236][3];				r_cell_reg[234] = inform_R[229][3];				r_cell_reg[235] = inform_R[237][3];				r_cell_reg[236] = inform_R[230][3];				r_cell_reg[237] = inform_R[238][3];				r_cell_reg[238] = inform_R[231][3];				r_cell_reg[239] = inform_R[239][3];				r_cell_reg[240] = inform_R[240][3];				r_cell_reg[241] = inform_R[248][3];				r_cell_reg[242] = inform_R[241][3];				r_cell_reg[243] = inform_R[249][3];				r_cell_reg[244] = inform_R[242][3];				r_cell_reg[245] = inform_R[250][3];				r_cell_reg[246] = inform_R[243][3];				r_cell_reg[247] = inform_R[251][3];				r_cell_reg[248] = inform_R[244][3];				r_cell_reg[249] = inform_R[252][3];				r_cell_reg[250] = inform_R[245][3];				r_cell_reg[251] = inform_R[253][3];				r_cell_reg[252] = inform_R[246][3];				r_cell_reg[253] = inform_R[254][3];				r_cell_reg[254] = inform_R[247][3];				r_cell_reg[255] = inform_R[255][3];				r_cell_reg[256] = inform_R[256][3];				r_cell_reg[257] = inform_R[264][3];				r_cell_reg[258] = inform_R[257][3];				r_cell_reg[259] = inform_R[265][3];				r_cell_reg[260] = inform_R[258][3];				r_cell_reg[261] = inform_R[266][3];				r_cell_reg[262] = inform_R[259][3];				r_cell_reg[263] = inform_R[267][3];				r_cell_reg[264] = inform_R[260][3];				r_cell_reg[265] = inform_R[268][3];				r_cell_reg[266] = inform_R[261][3];				r_cell_reg[267] = inform_R[269][3];				r_cell_reg[268] = inform_R[262][3];				r_cell_reg[269] = inform_R[270][3];				r_cell_reg[270] = inform_R[263][3];				r_cell_reg[271] = inform_R[271][3];				r_cell_reg[272] = inform_R[272][3];				r_cell_reg[273] = inform_R[280][3];				r_cell_reg[274] = inform_R[273][3];				r_cell_reg[275] = inform_R[281][3];				r_cell_reg[276] = inform_R[274][3];				r_cell_reg[277] = inform_R[282][3];				r_cell_reg[278] = inform_R[275][3];				r_cell_reg[279] = inform_R[283][3];				r_cell_reg[280] = inform_R[276][3];				r_cell_reg[281] = inform_R[284][3];				r_cell_reg[282] = inform_R[277][3];				r_cell_reg[283] = inform_R[285][3];				r_cell_reg[284] = inform_R[278][3];				r_cell_reg[285] = inform_R[286][3];				r_cell_reg[286] = inform_R[279][3];				r_cell_reg[287] = inform_R[287][3];				r_cell_reg[288] = inform_R[288][3];				r_cell_reg[289] = inform_R[296][3];				r_cell_reg[290] = inform_R[289][3];				r_cell_reg[291] = inform_R[297][3];				r_cell_reg[292] = inform_R[290][3];				r_cell_reg[293] = inform_R[298][3];				r_cell_reg[294] = inform_R[291][3];				r_cell_reg[295] = inform_R[299][3];				r_cell_reg[296] = inform_R[292][3];				r_cell_reg[297] = inform_R[300][3];				r_cell_reg[298] = inform_R[293][3];				r_cell_reg[299] = inform_R[301][3];				r_cell_reg[300] = inform_R[294][3];				r_cell_reg[301] = inform_R[302][3];				r_cell_reg[302] = inform_R[295][3];				r_cell_reg[303] = inform_R[303][3];				r_cell_reg[304] = inform_R[304][3];				r_cell_reg[305] = inform_R[312][3];				r_cell_reg[306] = inform_R[305][3];				r_cell_reg[307] = inform_R[313][3];				r_cell_reg[308] = inform_R[306][3];				r_cell_reg[309] = inform_R[314][3];				r_cell_reg[310] = inform_R[307][3];				r_cell_reg[311] = inform_R[315][3];				r_cell_reg[312] = inform_R[308][3];				r_cell_reg[313] = inform_R[316][3];				r_cell_reg[314] = inform_R[309][3];				r_cell_reg[315] = inform_R[317][3];				r_cell_reg[316] = inform_R[310][3];				r_cell_reg[317] = inform_R[318][3];				r_cell_reg[318] = inform_R[311][3];				r_cell_reg[319] = inform_R[319][3];				r_cell_reg[320] = inform_R[320][3];				r_cell_reg[321] = inform_R[328][3];				r_cell_reg[322] = inform_R[321][3];				r_cell_reg[323] = inform_R[329][3];				r_cell_reg[324] = inform_R[322][3];				r_cell_reg[325] = inform_R[330][3];				r_cell_reg[326] = inform_R[323][3];				r_cell_reg[327] = inform_R[331][3];				r_cell_reg[328] = inform_R[324][3];				r_cell_reg[329] = inform_R[332][3];				r_cell_reg[330] = inform_R[325][3];				r_cell_reg[331] = inform_R[333][3];				r_cell_reg[332] = inform_R[326][3];				r_cell_reg[333] = inform_R[334][3];				r_cell_reg[334] = inform_R[327][3];				r_cell_reg[335] = inform_R[335][3];				r_cell_reg[336] = inform_R[336][3];				r_cell_reg[337] = inform_R[344][3];				r_cell_reg[338] = inform_R[337][3];				r_cell_reg[339] = inform_R[345][3];				r_cell_reg[340] = inform_R[338][3];				r_cell_reg[341] = inform_R[346][3];				r_cell_reg[342] = inform_R[339][3];				r_cell_reg[343] = inform_R[347][3];				r_cell_reg[344] = inform_R[340][3];				r_cell_reg[345] = inform_R[348][3];				r_cell_reg[346] = inform_R[341][3];				r_cell_reg[347] = inform_R[349][3];				r_cell_reg[348] = inform_R[342][3];				r_cell_reg[349] = inform_R[350][3];				r_cell_reg[350] = inform_R[343][3];				r_cell_reg[351] = inform_R[351][3];				r_cell_reg[352] = inform_R[352][3];				r_cell_reg[353] = inform_R[360][3];				r_cell_reg[354] = inform_R[353][3];				r_cell_reg[355] = inform_R[361][3];				r_cell_reg[356] = inform_R[354][3];				r_cell_reg[357] = inform_R[362][3];				r_cell_reg[358] = inform_R[355][3];				r_cell_reg[359] = inform_R[363][3];				r_cell_reg[360] = inform_R[356][3];				r_cell_reg[361] = inform_R[364][3];				r_cell_reg[362] = inform_R[357][3];				r_cell_reg[363] = inform_R[365][3];				r_cell_reg[364] = inform_R[358][3];				r_cell_reg[365] = inform_R[366][3];				r_cell_reg[366] = inform_R[359][3];				r_cell_reg[367] = inform_R[367][3];				r_cell_reg[368] = inform_R[368][3];				r_cell_reg[369] = inform_R[376][3];				r_cell_reg[370] = inform_R[369][3];				r_cell_reg[371] = inform_R[377][3];				r_cell_reg[372] = inform_R[370][3];				r_cell_reg[373] = inform_R[378][3];				r_cell_reg[374] = inform_R[371][3];				r_cell_reg[375] = inform_R[379][3];				r_cell_reg[376] = inform_R[372][3];				r_cell_reg[377] = inform_R[380][3];				r_cell_reg[378] = inform_R[373][3];				r_cell_reg[379] = inform_R[381][3];				r_cell_reg[380] = inform_R[374][3];				r_cell_reg[381] = inform_R[382][3];				r_cell_reg[382] = inform_R[375][3];				r_cell_reg[383] = inform_R[383][3];				r_cell_reg[384] = inform_R[384][3];				r_cell_reg[385] = inform_R[392][3];				r_cell_reg[386] = inform_R[385][3];				r_cell_reg[387] = inform_R[393][3];				r_cell_reg[388] = inform_R[386][3];				r_cell_reg[389] = inform_R[394][3];				r_cell_reg[390] = inform_R[387][3];				r_cell_reg[391] = inform_R[395][3];				r_cell_reg[392] = inform_R[388][3];				r_cell_reg[393] = inform_R[396][3];				r_cell_reg[394] = inform_R[389][3];				r_cell_reg[395] = inform_R[397][3];				r_cell_reg[396] = inform_R[390][3];				r_cell_reg[397] = inform_R[398][3];				r_cell_reg[398] = inform_R[391][3];				r_cell_reg[399] = inform_R[399][3];				r_cell_reg[400] = inform_R[400][3];				r_cell_reg[401] = inform_R[408][3];				r_cell_reg[402] = inform_R[401][3];				r_cell_reg[403] = inform_R[409][3];				r_cell_reg[404] = inform_R[402][3];				r_cell_reg[405] = inform_R[410][3];				r_cell_reg[406] = inform_R[403][3];				r_cell_reg[407] = inform_R[411][3];				r_cell_reg[408] = inform_R[404][3];				r_cell_reg[409] = inform_R[412][3];				r_cell_reg[410] = inform_R[405][3];				r_cell_reg[411] = inform_R[413][3];				r_cell_reg[412] = inform_R[406][3];				r_cell_reg[413] = inform_R[414][3];				r_cell_reg[414] = inform_R[407][3];				r_cell_reg[415] = inform_R[415][3];				r_cell_reg[416] = inform_R[416][3];				r_cell_reg[417] = inform_R[424][3];				r_cell_reg[418] = inform_R[417][3];				r_cell_reg[419] = inform_R[425][3];				r_cell_reg[420] = inform_R[418][3];				r_cell_reg[421] = inform_R[426][3];				r_cell_reg[422] = inform_R[419][3];				r_cell_reg[423] = inform_R[427][3];				r_cell_reg[424] = inform_R[420][3];				r_cell_reg[425] = inform_R[428][3];				r_cell_reg[426] = inform_R[421][3];				r_cell_reg[427] = inform_R[429][3];				r_cell_reg[428] = inform_R[422][3];				r_cell_reg[429] = inform_R[430][3];				r_cell_reg[430] = inform_R[423][3];				r_cell_reg[431] = inform_R[431][3];				r_cell_reg[432] = inform_R[432][3];				r_cell_reg[433] = inform_R[440][3];				r_cell_reg[434] = inform_R[433][3];				r_cell_reg[435] = inform_R[441][3];				r_cell_reg[436] = inform_R[434][3];				r_cell_reg[437] = inform_R[442][3];				r_cell_reg[438] = inform_R[435][3];				r_cell_reg[439] = inform_R[443][3];				r_cell_reg[440] = inform_R[436][3];				r_cell_reg[441] = inform_R[444][3];				r_cell_reg[442] = inform_R[437][3];				r_cell_reg[443] = inform_R[445][3];				r_cell_reg[444] = inform_R[438][3];				r_cell_reg[445] = inform_R[446][3];				r_cell_reg[446] = inform_R[439][3];				r_cell_reg[447] = inform_R[447][3];				r_cell_reg[448] = inform_R[448][3];				r_cell_reg[449] = inform_R[456][3];				r_cell_reg[450] = inform_R[449][3];				r_cell_reg[451] = inform_R[457][3];				r_cell_reg[452] = inform_R[450][3];				r_cell_reg[453] = inform_R[458][3];				r_cell_reg[454] = inform_R[451][3];				r_cell_reg[455] = inform_R[459][3];				r_cell_reg[456] = inform_R[452][3];				r_cell_reg[457] = inform_R[460][3];				r_cell_reg[458] = inform_R[453][3];				r_cell_reg[459] = inform_R[461][3];				r_cell_reg[460] = inform_R[454][3];				r_cell_reg[461] = inform_R[462][3];				r_cell_reg[462] = inform_R[455][3];				r_cell_reg[463] = inform_R[463][3];				r_cell_reg[464] = inform_R[464][3];				r_cell_reg[465] = inform_R[472][3];				r_cell_reg[466] = inform_R[465][3];				r_cell_reg[467] = inform_R[473][3];				r_cell_reg[468] = inform_R[466][3];				r_cell_reg[469] = inform_R[474][3];				r_cell_reg[470] = inform_R[467][3];				r_cell_reg[471] = inform_R[475][3];				r_cell_reg[472] = inform_R[468][3];				r_cell_reg[473] = inform_R[476][3];				r_cell_reg[474] = inform_R[469][3];				r_cell_reg[475] = inform_R[477][3];				r_cell_reg[476] = inform_R[470][3];				r_cell_reg[477] = inform_R[478][3];				r_cell_reg[478] = inform_R[471][3];				r_cell_reg[479] = inform_R[479][3];				r_cell_reg[480] = inform_R[480][3];				r_cell_reg[481] = inform_R[488][3];				r_cell_reg[482] = inform_R[481][3];				r_cell_reg[483] = inform_R[489][3];				r_cell_reg[484] = inform_R[482][3];				r_cell_reg[485] = inform_R[490][3];				r_cell_reg[486] = inform_R[483][3];				r_cell_reg[487] = inform_R[491][3];				r_cell_reg[488] = inform_R[484][3];				r_cell_reg[489] = inform_R[492][3];				r_cell_reg[490] = inform_R[485][3];				r_cell_reg[491] = inform_R[493][3];				r_cell_reg[492] = inform_R[486][3];				r_cell_reg[493] = inform_R[494][3];				r_cell_reg[494] = inform_R[487][3];				r_cell_reg[495] = inform_R[495][3];				r_cell_reg[496] = inform_R[496][3];				r_cell_reg[497] = inform_R[504][3];				r_cell_reg[498] = inform_R[497][3];				r_cell_reg[499] = inform_R[505][3];				r_cell_reg[500] = inform_R[498][3];				r_cell_reg[501] = inform_R[506][3];				r_cell_reg[502] = inform_R[499][3];				r_cell_reg[503] = inform_R[507][3];				r_cell_reg[504] = inform_R[500][3];				r_cell_reg[505] = inform_R[508][3];				r_cell_reg[506] = inform_R[501][3];				r_cell_reg[507] = inform_R[509][3];				r_cell_reg[508] = inform_R[502][3];				r_cell_reg[509] = inform_R[510][3];				r_cell_reg[510] = inform_R[503][3];				r_cell_reg[511] = inform_R[511][3];				r_cell_reg[512] = inform_R[512][3];				r_cell_reg[513] = inform_R[520][3];				r_cell_reg[514] = inform_R[513][3];				r_cell_reg[515] = inform_R[521][3];				r_cell_reg[516] = inform_R[514][3];				r_cell_reg[517] = inform_R[522][3];				r_cell_reg[518] = inform_R[515][3];				r_cell_reg[519] = inform_R[523][3];				r_cell_reg[520] = inform_R[516][3];				r_cell_reg[521] = inform_R[524][3];				r_cell_reg[522] = inform_R[517][3];				r_cell_reg[523] = inform_R[525][3];				r_cell_reg[524] = inform_R[518][3];				r_cell_reg[525] = inform_R[526][3];				r_cell_reg[526] = inform_R[519][3];				r_cell_reg[527] = inform_R[527][3];				r_cell_reg[528] = inform_R[528][3];				r_cell_reg[529] = inform_R[536][3];				r_cell_reg[530] = inform_R[529][3];				r_cell_reg[531] = inform_R[537][3];				r_cell_reg[532] = inform_R[530][3];				r_cell_reg[533] = inform_R[538][3];				r_cell_reg[534] = inform_R[531][3];				r_cell_reg[535] = inform_R[539][3];				r_cell_reg[536] = inform_R[532][3];				r_cell_reg[537] = inform_R[540][3];				r_cell_reg[538] = inform_R[533][3];				r_cell_reg[539] = inform_R[541][3];				r_cell_reg[540] = inform_R[534][3];				r_cell_reg[541] = inform_R[542][3];				r_cell_reg[542] = inform_R[535][3];				r_cell_reg[543] = inform_R[543][3];				r_cell_reg[544] = inform_R[544][3];				r_cell_reg[545] = inform_R[552][3];				r_cell_reg[546] = inform_R[545][3];				r_cell_reg[547] = inform_R[553][3];				r_cell_reg[548] = inform_R[546][3];				r_cell_reg[549] = inform_R[554][3];				r_cell_reg[550] = inform_R[547][3];				r_cell_reg[551] = inform_R[555][3];				r_cell_reg[552] = inform_R[548][3];				r_cell_reg[553] = inform_R[556][3];				r_cell_reg[554] = inform_R[549][3];				r_cell_reg[555] = inform_R[557][3];				r_cell_reg[556] = inform_R[550][3];				r_cell_reg[557] = inform_R[558][3];				r_cell_reg[558] = inform_R[551][3];				r_cell_reg[559] = inform_R[559][3];				r_cell_reg[560] = inform_R[560][3];				r_cell_reg[561] = inform_R[568][3];				r_cell_reg[562] = inform_R[561][3];				r_cell_reg[563] = inform_R[569][3];				r_cell_reg[564] = inform_R[562][3];				r_cell_reg[565] = inform_R[570][3];				r_cell_reg[566] = inform_R[563][3];				r_cell_reg[567] = inform_R[571][3];				r_cell_reg[568] = inform_R[564][3];				r_cell_reg[569] = inform_R[572][3];				r_cell_reg[570] = inform_R[565][3];				r_cell_reg[571] = inform_R[573][3];				r_cell_reg[572] = inform_R[566][3];				r_cell_reg[573] = inform_R[574][3];				r_cell_reg[574] = inform_R[567][3];				r_cell_reg[575] = inform_R[575][3];				r_cell_reg[576] = inform_R[576][3];				r_cell_reg[577] = inform_R[584][3];				r_cell_reg[578] = inform_R[577][3];				r_cell_reg[579] = inform_R[585][3];				r_cell_reg[580] = inform_R[578][3];				r_cell_reg[581] = inform_R[586][3];				r_cell_reg[582] = inform_R[579][3];				r_cell_reg[583] = inform_R[587][3];				r_cell_reg[584] = inform_R[580][3];				r_cell_reg[585] = inform_R[588][3];				r_cell_reg[586] = inform_R[581][3];				r_cell_reg[587] = inform_R[589][3];				r_cell_reg[588] = inform_R[582][3];				r_cell_reg[589] = inform_R[590][3];				r_cell_reg[590] = inform_R[583][3];				r_cell_reg[591] = inform_R[591][3];				r_cell_reg[592] = inform_R[592][3];				r_cell_reg[593] = inform_R[600][3];				r_cell_reg[594] = inform_R[593][3];				r_cell_reg[595] = inform_R[601][3];				r_cell_reg[596] = inform_R[594][3];				r_cell_reg[597] = inform_R[602][3];				r_cell_reg[598] = inform_R[595][3];				r_cell_reg[599] = inform_R[603][3];				r_cell_reg[600] = inform_R[596][3];				r_cell_reg[601] = inform_R[604][3];				r_cell_reg[602] = inform_R[597][3];				r_cell_reg[603] = inform_R[605][3];				r_cell_reg[604] = inform_R[598][3];				r_cell_reg[605] = inform_R[606][3];				r_cell_reg[606] = inform_R[599][3];				r_cell_reg[607] = inform_R[607][3];				r_cell_reg[608] = inform_R[608][3];				r_cell_reg[609] = inform_R[616][3];				r_cell_reg[610] = inform_R[609][3];				r_cell_reg[611] = inform_R[617][3];				r_cell_reg[612] = inform_R[610][3];				r_cell_reg[613] = inform_R[618][3];				r_cell_reg[614] = inform_R[611][3];				r_cell_reg[615] = inform_R[619][3];				r_cell_reg[616] = inform_R[612][3];				r_cell_reg[617] = inform_R[620][3];				r_cell_reg[618] = inform_R[613][3];				r_cell_reg[619] = inform_R[621][3];				r_cell_reg[620] = inform_R[614][3];				r_cell_reg[621] = inform_R[622][3];				r_cell_reg[622] = inform_R[615][3];				r_cell_reg[623] = inform_R[623][3];				r_cell_reg[624] = inform_R[624][3];				r_cell_reg[625] = inform_R[632][3];				r_cell_reg[626] = inform_R[625][3];				r_cell_reg[627] = inform_R[633][3];				r_cell_reg[628] = inform_R[626][3];				r_cell_reg[629] = inform_R[634][3];				r_cell_reg[630] = inform_R[627][3];				r_cell_reg[631] = inform_R[635][3];				r_cell_reg[632] = inform_R[628][3];				r_cell_reg[633] = inform_R[636][3];				r_cell_reg[634] = inform_R[629][3];				r_cell_reg[635] = inform_R[637][3];				r_cell_reg[636] = inform_R[630][3];				r_cell_reg[637] = inform_R[638][3];				r_cell_reg[638] = inform_R[631][3];				r_cell_reg[639] = inform_R[639][3];				r_cell_reg[640] = inform_R[640][3];				r_cell_reg[641] = inform_R[648][3];				r_cell_reg[642] = inform_R[641][3];				r_cell_reg[643] = inform_R[649][3];				r_cell_reg[644] = inform_R[642][3];				r_cell_reg[645] = inform_R[650][3];				r_cell_reg[646] = inform_R[643][3];				r_cell_reg[647] = inform_R[651][3];				r_cell_reg[648] = inform_R[644][3];				r_cell_reg[649] = inform_R[652][3];				r_cell_reg[650] = inform_R[645][3];				r_cell_reg[651] = inform_R[653][3];				r_cell_reg[652] = inform_R[646][3];				r_cell_reg[653] = inform_R[654][3];				r_cell_reg[654] = inform_R[647][3];				r_cell_reg[655] = inform_R[655][3];				r_cell_reg[656] = inform_R[656][3];				r_cell_reg[657] = inform_R[664][3];				r_cell_reg[658] = inform_R[657][3];				r_cell_reg[659] = inform_R[665][3];				r_cell_reg[660] = inform_R[658][3];				r_cell_reg[661] = inform_R[666][3];				r_cell_reg[662] = inform_R[659][3];				r_cell_reg[663] = inform_R[667][3];				r_cell_reg[664] = inform_R[660][3];				r_cell_reg[665] = inform_R[668][3];				r_cell_reg[666] = inform_R[661][3];				r_cell_reg[667] = inform_R[669][3];				r_cell_reg[668] = inform_R[662][3];				r_cell_reg[669] = inform_R[670][3];				r_cell_reg[670] = inform_R[663][3];				r_cell_reg[671] = inform_R[671][3];				r_cell_reg[672] = inform_R[672][3];				r_cell_reg[673] = inform_R[680][3];				r_cell_reg[674] = inform_R[673][3];				r_cell_reg[675] = inform_R[681][3];				r_cell_reg[676] = inform_R[674][3];				r_cell_reg[677] = inform_R[682][3];				r_cell_reg[678] = inform_R[675][3];				r_cell_reg[679] = inform_R[683][3];				r_cell_reg[680] = inform_R[676][3];				r_cell_reg[681] = inform_R[684][3];				r_cell_reg[682] = inform_R[677][3];				r_cell_reg[683] = inform_R[685][3];				r_cell_reg[684] = inform_R[678][3];				r_cell_reg[685] = inform_R[686][3];				r_cell_reg[686] = inform_R[679][3];				r_cell_reg[687] = inform_R[687][3];				r_cell_reg[688] = inform_R[688][3];				r_cell_reg[689] = inform_R[696][3];				r_cell_reg[690] = inform_R[689][3];				r_cell_reg[691] = inform_R[697][3];				r_cell_reg[692] = inform_R[690][3];				r_cell_reg[693] = inform_R[698][3];				r_cell_reg[694] = inform_R[691][3];				r_cell_reg[695] = inform_R[699][3];				r_cell_reg[696] = inform_R[692][3];				r_cell_reg[697] = inform_R[700][3];				r_cell_reg[698] = inform_R[693][3];				r_cell_reg[699] = inform_R[701][3];				r_cell_reg[700] = inform_R[694][3];				r_cell_reg[701] = inform_R[702][3];				r_cell_reg[702] = inform_R[695][3];				r_cell_reg[703] = inform_R[703][3];				r_cell_reg[704] = inform_R[704][3];				r_cell_reg[705] = inform_R[712][3];				r_cell_reg[706] = inform_R[705][3];				r_cell_reg[707] = inform_R[713][3];				r_cell_reg[708] = inform_R[706][3];				r_cell_reg[709] = inform_R[714][3];				r_cell_reg[710] = inform_R[707][3];				r_cell_reg[711] = inform_R[715][3];				r_cell_reg[712] = inform_R[708][3];				r_cell_reg[713] = inform_R[716][3];				r_cell_reg[714] = inform_R[709][3];				r_cell_reg[715] = inform_R[717][3];				r_cell_reg[716] = inform_R[710][3];				r_cell_reg[717] = inform_R[718][3];				r_cell_reg[718] = inform_R[711][3];				r_cell_reg[719] = inform_R[719][3];				r_cell_reg[720] = inform_R[720][3];				r_cell_reg[721] = inform_R[728][3];				r_cell_reg[722] = inform_R[721][3];				r_cell_reg[723] = inform_R[729][3];				r_cell_reg[724] = inform_R[722][3];				r_cell_reg[725] = inform_R[730][3];				r_cell_reg[726] = inform_R[723][3];				r_cell_reg[727] = inform_R[731][3];				r_cell_reg[728] = inform_R[724][3];				r_cell_reg[729] = inform_R[732][3];				r_cell_reg[730] = inform_R[725][3];				r_cell_reg[731] = inform_R[733][3];				r_cell_reg[732] = inform_R[726][3];				r_cell_reg[733] = inform_R[734][3];				r_cell_reg[734] = inform_R[727][3];				r_cell_reg[735] = inform_R[735][3];				r_cell_reg[736] = inform_R[736][3];				r_cell_reg[737] = inform_R[744][3];				r_cell_reg[738] = inform_R[737][3];				r_cell_reg[739] = inform_R[745][3];				r_cell_reg[740] = inform_R[738][3];				r_cell_reg[741] = inform_R[746][3];				r_cell_reg[742] = inform_R[739][3];				r_cell_reg[743] = inform_R[747][3];				r_cell_reg[744] = inform_R[740][3];				r_cell_reg[745] = inform_R[748][3];				r_cell_reg[746] = inform_R[741][3];				r_cell_reg[747] = inform_R[749][3];				r_cell_reg[748] = inform_R[742][3];				r_cell_reg[749] = inform_R[750][3];				r_cell_reg[750] = inform_R[743][3];				r_cell_reg[751] = inform_R[751][3];				r_cell_reg[752] = inform_R[752][3];				r_cell_reg[753] = inform_R[760][3];				r_cell_reg[754] = inform_R[753][3];				r_cell_reg[755] = inform_R[761][3];				r_cell_reg[756] = inform_R[754][3];				r_cell_reg[757] = inform_R[762][3];				r_cell_reg[758] = inform_R[755][3];				r_cell_reg[759] = inform_R[763][3];				r_cell_reg[760] = inform_R[756][3];				r_cell_reg[761] = inform_R[764][3];				r_cell_reg[762] = inform_R[757][3];				r_cell_reg[763] = inform_R[765][3];				r_cell_reg[764] = inform_R[758][3];				r_cell_reg[765] = inform_R[766][3];				r_cell_reg[766] = inform_R[759][3];				r_cell_reg[767] = inform_R[767][3];				r_cell_reg[768] = inform_R[768][3];				r_cell_reg[769] = inform_R[776][3];				r_cell_reg[770] = inform_R[769][3];				r_cell_reg[771] = inform_R[777][3];				r_cell_reg[772] = inform_R[770][3];				r_cell_reg[773] = inform_R[778][3];				r_cell_reg[774] = inform_R[771][3];				r_cell_reg[775] = inform_R[779][3];				r_cell_reg[776] = inform_R[772][3];				r_cell_reg[777] = inform_R[780][3];				r_cell_reg[778] = inform_R[773][3];				r_cell_reg[779] = inform_R[781][3];				r_cell_reg[780] = inform_R[774][3];				r_cell_reg[781] = inform_R[782][3];				r_cell_reg[782] = inform_R[775][3];				r_cell_reg[783] = inform_R[783][3];				r_cell_reg[784] = inform_R[784][3];				r_cell_reg[785] = inform_R[792][3];				r_cell_reg[786] = inform_R[785][3];				r_cell_reg[787] = inform_R[793][3];				r_cell_reg[788] = inform_R[786][3];				r_cell_reg[789] = inform_R[794][3];				r_cell_reg[790] = inform_R[787][3];				r_cell_reg[791] = inform_R[795][3];				r_cell_reg[792] = inform_R[788][3];				r_cell_reg[793] = inform_R[796][3];				r_cell_reg[794] = inform_R[789][3];				r_cell_reg[795] = inform_R[797][3];				r_cell_reg[796] = inform_R[790][3];				r_cell_reg[797] = inform_R[798][3];				r_cell_reg[798] = inform_R[791][3];				r_cell_reg[799] = inform_R[799][3];				r_cell_reg[800] = inform_R[800][3];				r_cell_reg[801] = inform_R[808][3];				r_cell_reg[802] = inform_R[801][3];				r_cell_reg[803] = inform_R[809][3];				r_cell_reg[804] = inform_R[802][3];				r_cell_reg[805] = inform_R[810][3];				r_cell_reg[806] = inform_R[803][3];				r_cell_reg[807] = inform_R[811][3];				r_cell_reg[808] = inform_R[804][3];				r_cell_reg[809] = inform_R[812][3];				r_cell_reg[810] = inform_R[805][3];				r_cell_reg[811] = inform_R[813][3];				r_cell_reg[812] = inform_R[806][3];				r_cell_reg[813] = inform_R[814][3];				r_cell_reg[814] = inform_R[807][3];				r_cell_reg[815] = inform_R[815][3];				r_cell_reg[816] = inform_R[816][3];				r_cell_reg[817] = inform_R[824][3];				r_cell_reg[818] = inform_R[817][3];				r_cell_reg[819] = inform_R[825][3];				r_cell_reg[820] = inform_R[818][3];				r_cell_reg[821] = inform_R[826][3];				r_cell_reg[822] = inform_R[819][3];				r_cell_reg[823] = inform_R[827][3];				r_cell_reg[824] = inform_R[820][3];				r_cell_reg[825] = inform_R[828][3];				r_cell_reg[826] = inform_R[821][3];				r_cell_reg[827] = inform_R[829][3];				r_cell_reg[828] = inform_R[822][3];				r_cell_reg[829] = inform_R[830][3];				r_cell_reg[830] = inform_R[823][3];				r_cell_reg[831] = inform_R[831][3];				r_cell_reg[832] = inform_R[832][3];				r_cell_reg[833] = inform_R[840][3];				r_cell_reg[834] = inform_R[833][3];				r_cell_reg[835] = inform_R[841][3];				r_cell_reg[836] = inform_R[834][3];				r_cell_reg[837] = inform_R[842][3];				r_cell_reg[838] = inform_R[835][3];				r_cell_reg[839] = inform_R[843][3];				r_cell_reg[840] = inform_R[836][3];				r_cell_reg[841] = inform_R[844][3];				r_cell_reg[842] = inform_R[837][3];				r_cell_reg[843] = inform_R[845][3];				r_cell_reg[844] = inform_R[838][3];				r_cell_reg[845] = inform_R[846][3];				r_cell_reg[846] = inform_R[839][3];				r_cell_reg[847] = inform_R[847][3];				r_cell_reg[848] = inform_R[848][3];				r_cell_reg[849] = inform_R[856][3];				r_cell_reg[850] = inform_R[849][3];				r_cell_reg[851] = inform_R[857][3];				r_cell_reg[852] = inform_R[850][3];				r_cell_reg[853] = inform_R[858][3];				r_cell_reg[854] = inform_R[851][3];				r_cell_reg[855] = inform_R[859][3];				r_cell_reg[856] = inform_R[852][3];				r_cell_reg[857] = inform_R[860][3];				r_cell_reg[858] = inform_R[853][3];				r_cell_reg[859] = inform_R[861][3];				r_cell_reg[860] = inform_R[854][3];				r_cell_reg[861] = inform_R[862][3];				r_cell_reg[862] = inform_R[855][3];				r_cell_reg[863] = inform_R[863][3];				r_cell_reg[864] = inform_R[864][3];				r_cell_reg[865] = inform_R[872][3];				r_cell_reg[866] = inform_R[865][3];				r_cell_reg[867] = inform_R[873][3];				r_cell_reg[868] = inform_R[866][3];				r_cell_reg[869] = inform_R[874][3];				r_cell_reg[870] = inform_R[867][3];				r_cell_reg[871] = inform_R[875][3];				r_cell_reg[872] = inform_R[868][3];				r_cell_reg[873] = inform_R[876][3];				r_cell_reg[874] = inform_R[869][3];				r_cell_reg[875] = inform_R[877][3];				r_cell_reg[876] = inform_R[870][3];				r_cell_reg[877] = inform_R[878][3];				r_cell_reg[878] = inform_R[871][3];				r_cell_reg[879] = inform_R[879][3];				r_cell_reg[880] = inform_R[880][3];				r_cell_reg[881] = inform_R[888][3];				r_cell_reg[882] = inform_R[881][3];				r_cell_reg[883] = inform_R[889][3];				r_cell_reg[884] = inform_R[882][3];				r_cell_reg[885] = inform_R[890][3];				r_cell_reg[886] = inform_R[883][3];				r_cell_reg[887] = inform_R[891][3];				r_cell_reg[888] = inform_R[884][3];				r_cell_reg[889] = inform_R[892][3];				r_cell_reg[890] = inform_R[885][3];				r_cell_reg[891] = inform_R[893][3];				r_cell_reg[892] = inform_R[886][3];				r_cell_reg[893] = inform_R[894][3];				r_cell_reg[894] = inform_R[887][3];				r_cell_reg[895] = inform_R[895][3];				r_cell_reg[896] = inform_R[896][3];				r_cell_reg[897] = inform_R[904][3];				r_cell_reg[898] = inform_R[897][3];				r_cell_reg[899] = inform_R[905][3];				r_cell_reg[900] = inform_R[898][3];				r_cell_reg[901] = inform_R[906][3];				r_cell_reg[902] = inform_R[899][3];				r_cell_reg[903] = inform_R[907][3];				r_cell_reg[904] = inform_R[900][3];				r_cell_reg[905] = inform_R[908][3];				r_cell_reg[906] = inform_R[901][3];				r_cell_reg[907] = inform_R[909][3];				r_cell_reg[908] = inform_R[902][3];				r_cell_reg[909] = inform_R[910][3];				r_cell_reg[910] = inform_R[903][3];				r_cell_reg[911] = inform_R[911][3];				r_cell_reg[912] = inform_R[912][3];				r_cell_reg[913] = inform_R[920][3];				r_cell_reg[914] = inform_R[913][3];				r_cell_reg[915] = inform_R[921][3];				r_cell_reg[916] = inform_R[914][3];				r_cell_reg[917] = inform_R[922][3];				r_cell_reg[918] = inform_R[915][3];				r_cell_reg[919] = inform_R[923][3];				r_cell_reg[920] = inform_R[916][3];				r_cell_reg[921] = inform_R[924][3];				r_cell_reg[922] = inform_R[917][3];				r_cell_reg[923] = inform_R[925][3];				r_cell_reg[924] = inform_R[918][3];				r_cell_reg[925] = inform_R[926][3];				r_cell_reg[926] = inform_R[919][3];				r_cell_reg[927] = inform_R[927][3];				r_cell_reg[928] = inform_R[928][3];				r_cell_reg[929] = inform_R[936][3];				r_cell_reg[930] = inform_R[929][3];				r_cell_reg[931] = inform_R[937][3];				r_cell_reg[932] = inform_R[930][3];				r_cell_reg[933] = inform_R[938][3];				r_cell_reg[934] = inform_R[931][3];				r_cell_reg[935] = inform_R[939][3];				r_cell_reg[936] = inform_R[932][3];				r_cell_reg[937] = inform_R[940][3];				r_cell_reg[938] = inform_R[933][3];				r_cell_reg[939] = inform_R[941][3];				r_cell_reg[940] = inform_R[934][3];				r_cell_reg[941] = inform_R[942][3];				r_cell_reg[942] = inform_R[935][3];				r_cell_reg[943] = inform_R[943][3];				r_cell_reg[944] = inform_R[944][3];				r_cell_reg[945] = inform_R[952][3];				r_cell_reg[946] = inform_R[945][3];				r_cell_reg[947] = inform_R[953][3];				r_cell_reg[948] = inform_R[946][3];				r_cell_reg[949] = inform_R[954][3];				r_cell_reg[950] = inform_R[947][3];				r_cell_reg[951] = inform_R[955][3];				r_cell_reg[952] = inform_R[948][3];				r_cell_reg[953] = inform_R[956][3];				r_cell_reg[954] = inform_R[949][3];				r_cell_reg[955] = inform_R[957][3];				r_cell_reg[956] = inform_R[950][3];				r_cell_reg[957] = inform_R[958][3];				r_cell_reg[958] = inform_R[951][3];				r_cell_reg[959] = inform_R[959][3];				r_cell_reg[960] = inform_R[960][3];				r_cell_reg[961] = inform_R[968][3];				r_cell_reg[962] = inform_R[961][3];				r_cell_reg[963] = inform_R[969][3];				r_cell_reg[964] = inform_R[962][3];				r_cell_reg[965] = inform_R[970][3];				r_cell_reg[966] = inform_R[963][3];				r_cell_reg[967] = inform_R[971][3];				r_cell_reg[968] = inform_R[964][3];				r_cell_reg[969] = inform_R[972][3];				r_cell_reg[970] = inform_R[965][3];				r_cell_reg[971] = inform_R[973][3];				r_cell_reg[972] = inform_R[966][3];				r_cell_reg[973] = inform_R[974][3];				r_cell_reg[974] = inform_R[967][3];				r_cell_reg[975] = inform_R[975][3];				r_cell_reg[976] = inform_R[976][3];				r_cell_reg[977] = inform_R[984][3];				r_cell_reg[978] = inform_R[977][3];				r_cell_reg[979] = inform_R[985][3];				r_cell_reg[980] = inform_R[978][3];				r_cell_reg[981] = inform_R[986][3];				r_cell_reg[982] = inform_R[979][3];				r_cell_reg[983] = inform_R[987][3];				r_cell_reg[984] = inform_R[980][3];				r_cell_reg[985] = inform_R[988][3];				r_cell_reg[986] = inform_R[981][3];				r_cell_reg[987] = inform_R[989][3];				r_cell_reg[988] = inform_R[982][3];				r_cell_reg[989] = inform_R[990][3];				r_cell_reg[990] = inform_R[983][3];				r_cell_reg[991] = inform_R[991][3];				r_cell_reg[992] = inform_R[992][3];				r_cell_reg[993] = inform_R[1000][3];				r_cell_reg[994] = inform_R[993][3];				r_cell_reg[995] = inform_R[1001][3];				r_cell_reg[996] = inform_R[994][3];				r_cell_reg[997] = inform_R[1002][3];				r_cell_reg[998] = inform_R[995][3];				r_cell_reg[999] = inform_R[1003][3];				r_cell_reg[1000] = inform_R[996][3];				r_cell_reg[1001] = inform_R[1004][3];				r_cell_reg[1002] = inform_R[997][3];				r_cell_reg[1003] = inform_R[1005][3];				r_cell_reg[1004] = inform_R[998][3];				r_cell_reg[1005] = inform_R[1006][3];				r_cell_reg[1006] = inform_R[999][3];				r_cell_reg[1007] = inform_R[1007][3];				r_cell_reg[1008] = inform_R[1008][3];				r_cell_reg[1009] = inform_R[1016][3];				r_cell_reg[1010] = inform_R[1009][3];				r_cell_reg[1011] = inform_R[1017][3];				r_cell_reg[1012] = inform_R[1010][3];				r_cell_reg[1013] = inform_R[1018][3];				r_cell_reg[1014] = inform_R[1011][3];				r_cell_reg[1015] = inform_R[1019][3];				r_cell_reg[1016] = inform_R[1012][3];				r_cell_reg[1017] = inform_R[1020][3];				r_cell_reg[1018] = inform_R[1013][3];				r_cell_reg[1019] = inform_R[1021][3];				r_cell_reg[1020] = inform_R[1014][3];				r_cell_reg[1021] = inform_R[1022][3];				r_cell_reg[1022] = inform_R[1015][3];				r_cell_reg[1023] = inform_R[1023][3];				l_cell_reg[0] = inform_L[0][4];				l_cell_reg[1] = inform_L[8][4];				l_cell_reg[2] = inform_L[1][4];				l_cell_reg[3] = inform_L[9][4];				l_cell_reg[4] = inform_L[2][4];				l_cell_reg[5] = inform_L[10][4];				l_cell_reg[6] = inform_L[3][4];				l_cell_reg[7] = inform_L[11][4];				l_cell_reg[8] = inform_L[4][4];				l_cell_reg[9] = inform_L[12][4];				l_cell_reg[10] = inform_L[5][4];				l_cell_reg[11] = inform_L[13][4];				l_cell_reg[12] = inform_L[6][4];				l_cell_reg[13] = inform_L[14][4];				l_cell_reg[14] = inform_L[7][4];				l_cell_reg[15] = inform_L[15][4];				l_cell_reg[16] = inform_L[16][4];				l_cell_reg[17] = inform_L[24][4];				l_cell_reg[18] = inform_L[17][4];				l_cell_reg[19] = inform_L[25][4];				l_cell_reg[20] = inform_L[18][4];				l_cell_reg[21] = inform_L[26][4];				l_cell_reg[22] = inform_L[19][4];				l_cell_reg[23] = inform_L[27][4];				l_cell_reg[24] = inform_L[20][4];				l_cell_reg[25] = inform_L[28][4];				l_cell_reg[26] = inform_L[21][4];				l_cell_reg[27] = inform_L[29][4];				l_cell_reg[28] = inform_L[22][4];				l_cell_reg[29] = inform_L[30][4];				l_cell_reg[30] = inform_L[23][4];				l_cell_reg[31] = inform_L[31][4];				l_cell_reg[32] = inform_L[32][4];				l_cell_reg[33] = inform_L[40][4];				l_cell_reg[34] = inform_L[33][4];				l_cell_reg[35] = inform_L[41][4];				l_cell_reg[36] = inform_L[34][4];				l_cell_reg[37] = inform_L[42][4];				l_cell_reg[38] = inform_L[35][4];				l_cell_reg[39] = inform_L[43][4];				l_cell_reg[40] = inform_L[36][4];				l_cell_reg[41] = inform_L[44][4];				l_cell_reg[42] = inform_L[37][4];				l_cell_reg[43] = inform_L[45][4];				l_cell_reg[44] = inform_L[38][4];				l_cell_reg[45] = inform_L[46][4];				l_cell_reg[46] = inform_L[39][4];				l_cell_reg[47] = inform_L[47][4];				l_cell_reg[48] = inform_L[48][4];				l_cell_reg[49] = inform_L[56][4];				l_cell_reg[50] = inform_L[49][4];				l_cell_reg[51] = inform_L[57][4];				l_cell_reg[52] = inform_L[50][4];				l_cell_reg[53] = inform_L[58][4];				l_cell_reg[54] = inform_L[51][4];				l_cell_reg[55] = inform_L[59][4];				l_cell_reg[56] = inform_L[52][4];				l_cell_reg[57] = inform_L[60][4];				l_cell_reg[58] = inform_L[53][4];				l_cell_reg[59] = inform_L[61][4];				l_cell_reg[60] = inform_L[54][4];				l_cell_reg[61] = inform_L[62][4];				l_cell_reg[62] = inform_L[55][4];				l_cell_reg[63] = inform_L[63][4];				l_cell_reg[64] = inform_L[64][4];				l_cell_reg[65] = inform_L[72][4];				l_cell_reg[66] = inform_L[65][4];				l_cell_reg[67] = inform_L[73][4];				l_cell_reg[68] = inform_L[66][4];				l_cell_reg[69] = inform_L[74][4];				l_cell_reg[70] = inform_L[67][4];				l_cell_reg[71] = inform_L[75][4];				l_cell_reg[72] = inform_L[68][4];				l_cell_reg[73] = inform_L[76][4];				l_cell_reg[74] = inform_L[69][4];				l_cell_reg[75] = inform_L[77][4];				l_cell_reg[76] = inform_L[70][4];				l_cell_reg[77] = inform_L[78][4];				l_cell_reg[78] = inform_L[71][4];				l_cell_reg[79] = inform_L[79][4];				l_cell_reg[80] = inform_L[80][4];				l_cell_reg[81] = inform_L[88][4];				l_cell_reg[82] = inform_L[81][4];				l_cell_reg[83] = inform_L[89][4];				l_cell_reg[84] = inform_L[82][4];				l_cell_reg[85] = inform_L[90][4];				l_cell_reg[86] = inform_L[83][4];				l_cell_reg[87] = inform_L[91][4];				l_cell_reg[88] = inform_L[84][4];				l_cell_reg[89] = inform_L[92][4];				l_cell_reg[90] = inform_L[85][4];				l_cell_reg[91] = inform_L[93][4];				l_cell_reg[92] = inform_L[86][4];				l_cell_reg[93] = inform_L[94][4];				l_cell_reg[94] = inform_L[87][4];				l_cell_reg[95] = inform_L[95][4];				l_cell_reg[96] = inform_L[96][4];				l_cell_reg[97] = inform_L[104][4];				l_cell_reg[98] = inform_L[97][4];				l_cell_reg[99] = inform_L[105][4];				l_cell_reg[100] = inform_L[98][4];				l_cell_reg[101] = inform_L[106][4];				l_cell_reg[102] = inform_L[99][4];				l_cell_reg[103] = inform_L[107][4];				l_cell_reg[104] = inform_L[100][4];				l_cell_reg[105] = inform_L[108][4];				l_cell_reg[106] = inform_L[101][4];				l_cell_reg[107] = inform_L[109][4];				l_cell_reg[108] = inform_L[102][4];				l_cell_reg[109] = inform_L[110][4];				l_cell_reg[110] = inform_L[103][4];				l_cell_reg[111] = inform_L[111][4];				l_cell_reg[112] = inform_L[112][4];				l_cell_reg[113] = inform_L[120][4];				l_cell_reg[114] = inform_L[113][4];				l_cell_reg[115] = inform_L[121][4];				l_cell_reg[116] = inform_L[114][4];				l_cell_reg[117] = inform_L[122][4];				l_cell_reg[118] = inform_L[115][4];				l_cell_reg[119] = inform_L[123][4];				l_cell_reg[120] = inform_L[116][4];				l_cell_reg[121] = inform_L[124][4];				l_cell_reg[122] = inform_L[117][4];				l_cell_reg[123] = inform_L[125][4];				l_cell_reg[124] = inform_L[118][4];				l_cell_reg[125] = inform_L[126][4];				l_cell_reg[126] = inform_L[119][4];				l_cell_reg[127] = inform_L[127][4];				l_cell_reg[128] = inform_L[128][4];				l_cell_reg[129] = inform_L[136][4];				l_cell_reg[130] = inform_L[129][4];				l_cell_reg[131] = inform_L[137][4];				l_cell_reg[132] = inform_L[130][4];				l_cell_reg[133] = inform_L[138][4];				l_cell_reg[134] = inform_L[131][4];				l_cell_reg[135] = inform_L[139][4];				l_cell_reg[136] = inform_L[132][4];				l_cell_reg[137] = inform_L[140][4];				l_cell_reg[138] = inform_L[133][4];				l_cell_reg[139] = inform_L[141][4];				l_cell_reg[140] = inform_L[134][4];				l_cell_reg[141] = inform_L[142][4];				l_cell_reg[142] = inform_L[135][4];				l_cell_reg[143] = inform_L[143][4];				l_cell_reg[144] = inform_L[144][4];				l_cell_reg[145] = inform_L[152][4];				l_cell_reg[146] = inform_L[145][4];				l_cell_reg[147] = inform_L[153][4];				l_cell_reg[148] = inform_L[146][4];				l_cell_reg[149] = inform_L[154][4];				l_cell_reg[150] = inform_L[147][4];				l_cell_reg[151] = inform_L[155][4];				l_cell_reg[152] = inform_L[148][4];				l_cell_reg[153] = inform_L[156][4];				l_cell_reg[154] = inform_L[149][4];				l_cell_reg[155] = inform_L[157][4];				l_cell_reg[156] = inform_L[150][4];				l_cell_reg[157] = inform_L[158][4];				l_cell_reg[158] = inform_L[151][4];				l_cell_reg[159] = inform_L[159][4];				l_cell_reg[160] = inform_L[160][4];				l_cell_reg[161] = inform_L[168][4];				l_cell_reg[162] = inform_L[161][4];				l_cell_reg[163] = inform_L[169][4];				l_cell_reg[164] = inform_L[162][4];				l_cell_reg[165] = inform_L[170][4];				l_cell_reg[166] = inform_L[163][4];				l_cell_reg[167] = inform_L[171][4];				l_cell_reg[168] = inform_L[164][4];				l_cell_reg[169] = inform_L[172][4];				l_cell_reg[170] = inform_L[165][4];				l_cell_reg[171] = inform_L[173][4];				l_cell_reg[172] = inform_L[166][4];				l_cell_reg[173] = inform_L[174][4];				l_cell_reg[174] = inform_L[167][4];				l_cell_reg[175] = inform_L[175][4];				l_cell_reg[176] = inform_L[176][4];				l_cell_reg[177] = inform_L[184][4];				l_cell_reg[178] = inform_L[177][4];				l_cell_reg[179] = inform_L[185][4];				l_cell_reg[180] = inform_L[178][4];				l_cell_reg[181] = inform_L[186][4];				l_cell_reg[182] = inform_L[179][4];				l_cell_reg[183] = inform_L[187][4];				l_cell_reg[184] = inform_L[180][4];				l_cell_reg[185] = inform_L[188][4];				l_cell_reg[186] = inform_L[181][4];				l_cell_reg[187] = inform_L[189][4];				l_cell_reg[188] = inform_L[182][4];				l_cell_reg[189] = inform_L[190][4];				l_cell_reg[190] = inform_L[183][4];				l_cell_reg[191] = inform_L[191][4];				l_cell_reg[192] = inform_L[192][4];				l_cell_reg[193] = inform_L[200][4];				l_cell_reg[194] = inform_L[193][4];				l_cell_reg[195] = inform_L[201][4];				l_cell_reg[196] = inform_L[194][4];				l_cell_reg[197] = inform_L[202][4];				l_cell_reg[198] = inform_L[195][4];				l_cell_reg[199] = inform_L[203][4];				l_cell_reg[200] = inform_L[196][4];				l_cell_reg[201] = inform_L[204][4];				l_cell_reg[202] = inform_L[197][4];				l_cell_reg[203] = inform_L[205][4];				l_cell_reg[204] = inform_L[198][4];				l_cell_reg[205] = inform_L[206][4];				l_cell_reg[206] = inform_L[199][4];				l_cell_reg[207] = inform_L[207][4];				l_cell_reg[208] = inform_L[208][4];				l_cell_reg[209] = inform_L[216][4];				l_cell_reg[210] = inform_L[209][4];				l_cell_reg[211] = inform_L[217][4];				l_cell_reg[212] = inform_L[210][4];				l_cell_reg[213] = inform_L[218][4];				l_cell_reg[214] = inform_L[211][4];				l_cell_reg[215] = inform_L[219][4];				l_cell_reg[216] = inform_L[212][4];				l_cell_reg[217] = inform_L[220][4];				l_cell_reg[218] = inform_L[213][4];				l_cell_reg[219] = inform_L[221][4];				l_cell_reg[220] = inform_L[214][4];				l_cell_reg[221] = inform_L[222][4];				l_cell_reg[222] = inform_L[215][4];				l_cell_reg[223] = inform_L[223][4];				l_cell_reg[224] = inform_L[224][4];				l_cell_reg[225] = inform_L[232][4];				l_cell_reg[226] = inform_L[225][4];				l_cell_reg[227] = inform_L[233][4];				l_cell_reg[228] = inform_L[226][4];				l_cell_reg[229] = inform_L[234][4];				l_cell_reg[230] = inform_L[227][4];				l_cell_reg[231] = inform_L[235][4];				l_cell_reg[232] = inform_L[228][4];				l_cell_reg[233] = inform_L[236][4];				l_cell_reg[234] = inform_L[229][4];				l_cell_reg[235] = inform_L[237][4];				l_cell_reg[236] = inform_L[230][4];				l_cell_reg[237] = inform_L[238][4];				l_cell_reg[238] = inform_L[231][4];				l_cell_reg[239] = inform_L[239][4];				l_cell_reg[240] = inform_L[240][4];				l_cell_reg[241] = inform_L[248][4];				l_cell_reg[242] = inform_L[241][4];				l_cell_reg[243] = inform_L[249][4];				l_cell_reg[244] = inform_L[242][4];				l_cell_reg[245] = inform_L[250][4];				l_cell_reg[246] = inform_L[243][4];				l_cell_reg[247] = inform_L[251][4];				l_cell_reg[248] = inform_L[244][4];				l_cell_reg[249] = inform_L[252][4];				l_cell_reg[250] = inform_L[245][4];				l_cell_reg[251] = inform_L[253][4];				l_cell_reg[252] = inform_L[246][4];				l_cell_reg[253] = inform_L[254][4];				l_cell_reg[254] = inform_L[247][4];				l_cell_reg[255] = inform_L[255][4];				l_cell_reg[256] = inform_L[256][4];				l_cell_reg[257] = inform_L[264][4];				l_cell_reg[258] = inform_L[257][4];				l_cell_reg[259] = inform_L[265][4];				l_cell_reg[260] = inform_L[258][4];				l_cell_reg[261] = inform_L[266][4];				l_cell_reg[262] = inform_L[259][4];				l_cell_reg[263] = inform_L[267][4];				l_cell_reg[264] = inform_L[260][4];				l_cell_reg[265] = inform_L[268][4];				l_cell_reg[266] = inform_L[261][4];				l_cell_reg[267] = inform_L[269][4];				l_cell_reg[268] = inform_L[262][4];				l_cell_reg[269] = inform_L[270][4];				l_cell_reg[270] = inform_L[263][4];				l_cell_reg[271] = inform_L[271][4];				l_cell_reg[272] = inform_L[272][4];				l_cell_reg[273] = inform_L[280][4];				l_cell_reg[274] = inform_L[273][4];				l_cell_reg[275] = inform_L[281][4];				l_cell_reg[276] = inform_L[274][4];				l_cell_reg[277] = inform_L[282][4];				l_cell_reg[278] = inform_L[275][4];				l_cell_reg[279] = inform_L[283][4];				l_cell_reg[280] = inform_L[276][4];				l_cell_reg[281] = inform_L[284][4];				l_cell_reg[282] = inform_L[277][4];				l_cell_reg[283] = inform_L[285][4];				l_cell_reg[284] = inform_L[278][4];				l_cell_reg[285] = inform_L[286][4];				l_cell_reg[286] = inform_L[279][4];				l_cell_reg[287] = inform_L[287][4];				l_cell_reg[288] = inform_L[288][4];				l_cell_reg[289] = inform_L[296][4];				l_cell_reg[290] = inform_L[289][4];				l_cell_reg[291] = inform_L[297][4];				l_cell_reg[292] = inform_L[290][4];				l_cell_reg[293] = inform_L[298][4];				l_cell_reg[294] = inform_L[291][4];				l_cell_reg[295] = inform_L[299][4];				l_cell_reg[296] = inform_L[292][4];				l_cell_reg[297] = inform_L[300][4];				l_cell_reg[298] = inform_L[293][4];				l_cell_reg[299] = inform_L[301][4];				l_cell_reg[300] = inform_L[294][4];				l_cell_reg[301] = inform_L[302][4];				l_cell_reg[302] = inform_L[295][4];				l_cell_reg[303] = inform_L[303][4];				l_cell_reg[304] = inform_L[304][4];				l_cell_reg[305] = inform_L[312][4];				l_cell_reg[306] = inform_L[305][4];				l_cell_reg[307] = inform_L[313][4];				l_cell_reg[308] = inform_L[306][4];				l_cell_reg[309] = inform_L[314][4];				l_cell_reg[310] = inform_L[307][4];				l_cell_reg[311] = inform_L[315][4];				l_cell_reg[312] = inform_L[308][4];				l_cell_reg[313] = inform_L[316][4];				l_cell_reg[314] = inform_L[309][4];				l_cell_reg[315] = inform_L[317][4];				l_cell_reg[316] = inform_L[310][4];				l_cell_reg[317] = inform_L[318][4];				l_cell_reg[318] = inform_L[311][4];				l_cell_reg[319] = inform_L[319][4];				l_cell_reg[320] = inform_L[320][4];				l_cell_reg[321] = inform_L[328][4];				l_cell_reg[322] = inform_L[321][4];				l_cell_reg[323] = inform_L[329][4];				l_cell_reg[324] = inform_L[322][4];				l_cell_reg[325] = inform_L[330][4];				l_cell_reg[326] = inform_L[323][4];				l_cell_reg[327] = inform_L[331][4];				l_cell_reg[328] = inform_L[324][4];				l_cell_reg[329] = inform_L[332][4];				l_cell_reg[330] = inform_L[325][4];				l_cell_reg[331] = inform_L[333][4];				l_cell_reg[332] = inform_L[326][4];				l_cell_reg[333] = inform_L[334][4];				l_cell_reg[334] = inform_L[327][4];				l_cell_reg[335] = inform_L[335][4];				l_cell_reg[336] = inform_L[336][4];				l_cell_reg[337] = inform_L[344][4];				l_cell_reg[338] = inform_L[337][4];				l_cell_reg[339] = inform_L[345][4];				l_cell_reg[340] = inform_L[338][4];				l_cell_reg[341] = inform_L[346][4];				l_cell_reg[342] = inform_L[339][4];				l_cell_reg[343] = inform_L[347][4];				l_cell_reg[344] = inform_L[340][4];				l_cell_reg[345] = inform_L[348][4];				l_cell_reg[346] = inform_L[341][4];				l_cell_reg[347] = inform_L[349][4];				l_cell_reg[348] = inform_L[342][4];				l_cell_reg[349] = inform_L[350][4];				l_cell_reg[350] = inform_L[343][4];				l_cell_reg[351] = inform_L[351][4];				l_cell_reg[352] = inform_L[352][4];				l_cell_reg[353] = inform_L[360][4];				l_cell_reg[354] = inform_L[353][4];				l_cell_reg[355] = inform_L[361][4];				l_cell_reg[356] = inform_L[354][4];				l_cell_reg[357] = inform_L[362][4];				l_cell_reg[358] = inform_L[355][4];				l_cell_reg[359] = inform_L[363][4];				l_cell_reg[360] = inform_L[356][4];				l_cell_reg[361] = inform_L[364][4];				l_cell_reg[362] = inform_L[357][4];				l_cell_reg[363] = inform_L[365][4];				l_cell_reg[364] = inform_L[358][4];				l_cell_reg[365] = inform_L[366][4];				l_cell_reg[366] = inform_L[359][4];				l_cell_reg[367] = inform_L[367][4];				l_cell_reg[368] = inform_L[368][4];				l_cell_reg[369] = inform_L[376][4];				l_cell_reg[370] = inform_L[369][4];				l_cell_reg[371] = inform_L[377][4];				l_cell_reg[372] = inform_L[370][4];				l_cell_reg[373] = inform_L[378][4];				l_cell_reg[374] = inform_L[371][4];				l_cell_reg[375] = inform_L[379][4];				l_cell_reg[376] = inform_L[372][4];				l_cell_reg[377] = inform_L[380][4];				l_cell_reg[378] = inform_L[373][4];				l_cell_reg[379] = inform_L[381][4];				l_cell_reg[380] = inform_L[374][4];				l_cell_reg[381] = inform_L[382][4];				l_cell_reg[382] = inform_L[375][4];				l_cell_reg[383] = inform_L[383][4];				l_cell_reg[384] = inform_L[384][4];				l_cell_reg[385] = inform_L[392][4];				l_cell_reg[386] = inform_L[385][4];				l_cell_reg[387] = inform_L[393][4];				l_cell_reg[388] = inform_L[386][4];				l_cell_reg[389] = inform_L[394][4];				l_cell_reg[390] = inform_L[387][4];				l_cell_reg[391] = inform_L[395][4];				l_cell_reg[392] = inform_L[388][4];				l_cell_reg[393] = inform_L[396][4];				l_cell_reg[394] = inform_L[389][4];				l_cell_reg[395] = inform_L[397][4];				l_cell_reg[396] = inform_L[390][4];				l_cell_reg[397] = inform_L[398][4];				l_cell_reg[398] = inform_L[391][4];				l_cell_reg[399] = inform_L[399][4];				l_cell_reg[400] = inform_L[400][4];				l_cell_reg[401] = inform_L[408][4];				l_cell_reg[402] = inform_L[401][4];				l_cell_reg[403] = inform_L[409][4];				l_cell_reg[404] = inform_L[402][4];				l_cell_reg[405] = inform_L[410][4];				l_cell_reg[406] = inform_L[403][4];				l_cell_reg[407] = inform_L[411][4];				l_cell_reg[408] = inform_L[404][4];				l_cell_reg[409] = inform_L[412][4];				l_cell_reg[410] = inform_L[405][4];				l_cell_reg[411] = inform_L[413][4];				l_cell_reg[412] = inform_L[406][4];				l_cell_reg[413] = inform_L[414][4];				l_cell_reg[414] = inform_L[407][4];				l_cell_reg[415] = inform_L[415][4];				l_cell_reg[416] = inform_L[416][4];				l_cell_reg[417] = inform_L[424][4];				l_cell_reg[418] = inform_L[417][4];				l_cell_reg[419] = inform_L[425][4];				l_cell_reg[420] = inform_L[418][4];				l_cell_reg[421] = inform_L[426][4];				l_cell_reg[422] = inform_L[419][4];				l_cell_reg[423] = inform_L[427][4];				l_cell_reg[424] = inform_L[420][4];				l_cell_reg[425] = inform_L[428][4];				l_cell_reg[426] = inform_L[421][4];				l_cell_reg[427] = inform_L[429][4];				l_cell_reg[428] = inform_L[422][4];				l_cell_reg[429] = inform_L[430][4];				l_cell_reg[430] = inform_L[423][4];				l_cell_reg[431] = inform_L[431][4];				l_cell_reg[432] = inform_L[432][4];				l_cell_reg[433] = inform_L[440][4];				l_cell_reg[434] = inform_L[433][4];				l_cell_reg[435] = inform_L[441][4];				l_cell_reg[436] = inform_L[434][4];				l_cell_reg[437] = inform_L[442][4];				l_cell_reg[438] = inform_L[435][4];				l_cell_reg[439] = inform_L[443][4];				l_cell_reg[440] = inform_L[436][4];				l_cell_reg[441] = inform_L[444][4];				l_cell_reg[442] = inform_L[437][4];				l_cell_reg[443] = inform_L[445][4];				l_cell_reg[444] = inform_L[438][4];				l_cell_reg[445] = inform_L[446][4];				l_cell_reg[446] = inform_L[439][4];				l_cell_reg[447] = inform_L[447][4];				l_cell_reg[448] = inform_L[448][4];				l_cell_reg[449] = inform_L[456][4];				l_cell_reg[450] = inform_L[449][4];				l_cell_reg[451] = inform_L[457][4];				l_cell_reg[452] = inform_L[450][4];				l_cell_reg[453] = inform_L[458][4];				l_cell_reg[454] = inform_L[451][4];				l_cell_reg[455] = inform_L[459][4];				l_cell_reg[456] = inform_L[452][4];				l_cell_reg[457] = inform_L[460][4];				l_cell_reg[458] = inform_L[453][4];				l_cell_reg[459] = inform_L[461][4];				l_cell_reg[460] = inform_L[454][4];				l_cell_reg[461] = inform_L[462][4];				l_cell_reg[462] = inform_L[455][4];				l_cell_reg[463] = inform_L[463][4];				l_cell_reg[464] = inform_L[464][4];				l_cell_reg[465] = inform_L[472][4];				l_cell_reg[466] = inform_L[465][4];				l_cell_reg[467] = inform_L[473][4];				l_cell_reg[468] = inform_L[466][4];				l_cell_reg[469] = inform_L[474][4];				l_cell_reg[470] = inform_L[467][4];				l_cell_reg[471] = inform_L[475][4];				l_cell_reg[472] = inform_L[468][4];				l_cell_reg[473] = inform_L[476][4];				l_cell_reg[474] = inform_L[469][4];				l_cell_reg[475] = inform_L[477][4];				l_cell_reg[476] = inform_L[470][4];				l_cell_reg[477] = inform_L[478][4];				l_cell_reg[478] = inform_L[471][4];				l_cell_reg[479] = inform_L[479][4];				l_cell_reg[480] = inform_L[480][4];				l_cell_reg[481] = inform_L[488][4];				l_cell_reg[482] = inform_L[481][4];				l_cell_reg[483] = inform_L[489][4];				l_cell_reg[484] = inform_L[482][4];				l_cell_reg[485] = inform_L[490][4];				l_cell_reg[486] = inform_L[483][4];				l_cell_reg[487] = inform_L[491][4];				l_cell_reg[488] = inform_L[484][4];				l_cell_reg[489] = inform_L[492][4];				l_cell_reg[490] = inform_L[485][4];				l_cell_reg[491] = inform_L[493][4];				l_cell_reg[492] = inform_L[486][4];				l_cell_reg[493] = inform_L[494][4];				l_cell_reg[494] = inform_L[487][4];				l_cell_reg[495] = inform_L[495][4];				l_cell_reg[496] = inform_L[496][4];				l_cell_reg[497] = inform_L[504][4];				l_cell_reg[498] = inform_L[497][4];				l_cell_reg[499] = inform_L[505][4];				l_cell_reg[500] = inform_L[498][4];				l_cell_reg[501] = inform_L[506][4];				l_cell_reg[502] = inform_L[499][4];				l_cell_reg[503] = inform_L[507][4];				l_cell_reg[504] = inform_L[500][4];				l_cell_reg[505] = inform_L[508][4];				l_cell_reg[506] = inform_L[501][4];				l_cell_reg[507] = inform_L[509][4];				l_cell_reg[508] = inform_L[502][4];				l_cell_reg[509] = inform_L[510][4];				l_cell_reg[510] = inform_L[503][4];				l_cell_reg[511] = inform_L[511][4];				l_cell_reg[512] = inform_L[512][4];				l_cell_reg[513] = inform_L[520][4];				l_cell_reg[514] = inform_L[513][4];				l_cell_reg[515] = inform_L[521][4];				l_cell_reg[516] = inform_L[514][4];				l_cell_reg[517] = inform_L[522][4];				l_cell_reg[518] = inform_L[515][4];				l_cell_reg[519] = inform_L[523][4];				l_cell_reg[520] = inform_L[516][4];				l_cell_reg[521] = inform_L[524][4];				l_cell_reg[522] = inform_L[517][4];				l_cell_reg[523] = inform_L[525][4];				l_cell_reg[524] = inform_L[518][4];				l_cell_reg[525] = inform_L[526][4];				l_cell_reg[526] = inform_L[519][4];				l_cell_reg[527] = inform_L[527][4];				l_cell_reg[528] = inform_L[528][4];				l_cell_reg[529] = inform_L[536][4];				l_cell_reg[530] = inform_L[529][4];				l_cell_reg[531] = inform_L[537][4];				l_cell_reg[532] = inform_L[530][4];				l_cell_reg[533] = inform_L[538][4];				l_cell_reg[534] = inform_L[531][4];				l_cell_reg[535] = inform_L[539][4];				l_cell_reg[536] = inform_L[532][4];				l_cell_reg[537] = inform_L[540][4];				l_cell_reg[538] = inform_L[533][4];				l_cell_reg[539] = inform_L[541][4];				l_cell_reg[540] = inform_L[534][4];				l_cell_reg[541] = inform_L[542][4];				l_cell_reg[542] = inform_L[535][4];				l_cell_reg[543] = inform_L[543][4];				l_cell_reg[544] = inform_L[544][4];				l_cell_reg[545] = inform_L[552][4];				l_cell_reg[546] = inform_L[545][4];				l_cell_reg[547] = inform_L[553][4];				l_cell_reg[548] = inform_L[546][4];				l_cell_reg[549] = inform_L[554][4];				l_cell_reg[550] = inform_L[547][4];				l_cell_reg[551] = inform_L[555][4];				l_cell_reg[552] = inform_L[548][4];				l_cell_reg[553] = inform_L[556][4];				l_cell_reg[554] = inform_L[549][4];				l_cell_reg[555] = inform_L[557][4];				l_cell_reg[556] = inform_L[550][4];				l_cell_reg[557] = inform_L[558][4];				l_cell_reg[558] = inform_L[551][4];				l_cell_reg[559] = inform_L[559][4];				l_cell_reg[560] = inform_L[560][4];				l_cell_reg[561] = inform_L[568][4];				l_cell_reg[562] = inform_L[561][4];				l_cell_reg[563] = inform_L[569][4];				l_cell_reg[564] = inform_L[562][4];				l_cell_reg[565] = inform_L[570][4];				l_cell_reg[566] = inform_L[563][4];				l_cell_reg[567] = inform_L[571][4];				l_cell_reg[568] = inform_L[564][4];				l_cell_reg[569] = inform_L[572][4];				l_cell_reg[570] = inform_L[565][4];				l_cell_reg[571] = inform_L[573][4];				l_cell_reg[572] = inform_L[566][4];				l_cell_reg[573] = inform_L[574][4];				l_cell_reg[574] = inform_L[567][4];				l_cell_reg[575] = inform_L[575][4];				l_cell_reg[576] = inform_L[576][4];				l_cell_reg[577] = inform_L[584][4];				l_cell_reg[578] = inform_L[577][4];				l_cell_reg[579] = inform_L[585][4];				l_cell_reg[580] = inform_L[578][4];				l_cell_reg[581] = inform_L[586][4];				l_cell_reg[582] = inform_L[579][4];				l_cell_reg[583] = inform_L[587][4];				l_cell_reg[584] = inform_L[580][4];				l_cell_reg[585] = inform_L[588][4];				l_cell_reg[586] = inform_L[581][4];				l_cell_reg[587] = inform_L[589][4];				l_cell_reg[588] = inform_L[582][4];				l_cell_reg[589] = inform_L[590][4];				l_cell_reg[590] = inform_L[583][4];				l_cell_reg[591] = inform_L[591][4];				l_cell_reg[592] = inform_L[592][4];				l_cell_reg[593] = inform_L[600][4];				l_cell_reg[594] = inform_L[593][4];				l_cell_reg[595] = inform_L[601][4];				l_cell_reg[596] = inform_L[594][4];				l_cell_reg[597] = inform_L[602][4];				l_cell_reg[598] = inform_L[595][4];				l_cell_reg[599] = inform_L[603][4];				l_cell_reg[600] = inform_L[596][4];				l_cell_reg[601] = inform_L[604][4];				l_cell_reg[602] = inform_L[597][4];				l_cell_reg[603] = inform_L[605][4];				l_cell_reg[604] = inform_L[598][4];				l_cell_reg[605] = inform_L[606][4];				l_cell_reg[606] = inform_L[599][4];				l_cell_reg[607] = inform_L[607][4];				l_cell_reg[608] = inform_L[608][4];				l_cell_reg[609] = inform_L[616][4];				l_cell_reg[610] = inform_L[609][4];				l_cell_reg[611] = inform_L[617][4];				l_cell_reg[612] = inform_L[610][4];				l_cell_reg[613] = inform_L[618][4];				l_cell_reg[614] = inform_L[611][4];				l_cell_reg[615] = inform_L[619][4];				l_cell_reg[616] = inform_L[612][4];				l_cell_reg[617] = inform_L[620][4];				l_cell_reg[618] = inform_L[613][4];				l_cell_reg[619] = inform_L[621][4];				l_cell_reg[620] = inform_L[614][4];				l_cell_reg[621] = inform_L[622][4];				l_cell_reg[622] = inform_L[615][4];				l_cell_reg[623] = inform_L[623][4];				l_cell_reg[624] = inform_L[624][4];				l_cell_reg[625] = inform_L[632][4];				l_cell_reg[626] = inform_L[625][4];				l_cell_reg[627] = inform_L[633][4];				l_cell_reg[628] = inform_L[626][4];				l_cell_reg[629] = inform_L[634][4];				l_cell_reg[630] = inform_L[627][4];				l_cell_reg[631] = inform_L[635][4];				l_cell_reg[632] = inform_L[628][4];				l_cell_reg[633] = inform_L[636][4];				l_cell_reg[634] = inform_L[629][4];				l_cell_reg[635] = inform_L[637][4];				l_cell_reg[636] = inform_L[630][4];				l_cell_reg[637] = inform_L[638][4];				l_cell_reg[638] = inform_L[631][4];				l_cell_reg[639] = inform_L[639][4];				l_cell_reg[640] = inform_L[640][4];				l_cell_reg[641] = inform_L[648][4];				l_cell_reg[642] = inform_L[641][4];				l_cell_reg[643] = inform_L[649][4];				l_cell_reg[644] = inform_L[642][4];				l_cell_reg[645] = inform_L[650][4];				l_cell_reg[646] = inform_L[643][4];				l_cell_reg[647] = inform_L[651][4];				l_cell_reg[648] = inform_L[644][4];				l_cell_reg[649] = inform_L[652][4];				l_cell_reg[650] = inform_L[645][4];				l_cell_reg[651] = inform_L[653][4];				l_cell_reg[652] = inform_L[646][4];				l_cell_reg[653] = inform_L[654][4];				l_cell_reg[654] = inform_L[647][4];				l_cell_reg[655] = inform_L[655][4];				l_cell_reg[656] = inform_L[656][4];				l_cell_reg[657] = inform_L[664][4];				l_cell_reg[658] = inform_L[657][4];				l_cell_reg[659] = inform_L[665][4];				l_cell_reg[660] = inform_L[658][4];				l_cell_reg[661] = inform_L[666][4];				l_cell_reg[662] = inform_L[659][4];				l_cell_reg[663] = inform_L[667][4];				l_cell_reg[664] = inform_L[660][4];				l_cell_reg[665] = inform_L[668][4];				l_cell_reg[666] = inform_L[661][4];				l_cell_reg[667] = inform_L[669][4];				l_cell_reg[668] = inform_L[662][4];				l_cell_reg[669] = inform_L[670][4];				l_cell_reg[670] = inform_L[663][4];				l_cell_reg[671] = inform_L[671][4];				l_cell_reg[672] = inform_L[672][4];				l_cell_reg[673] = inform_L[680][4];				l_cell_reg[674] = inform_L[673][4];				l_cell_reg[675] = inform_L[681][4];				l_cell_reg[676] = inform_L[674][4];				l_cell_reg[677] = inform_L[682][4];				l_cell_reg[678] = inform_L[675][4];				l_cell_reg[679] = inform_L[683][4];				l_cell_reg[680] = inform_L[676][4];				l_cell_reg[681] = inform_L[684][4];				l_cell_reg[682] = inform_L[677][4];				l_cell_reg[683] = inform_L[685][4];				l_cell_reg[684] = inform_L[678][4];				l_cell_reg[685] = inform_L[686][4];				l_cell_reg[686] = inform_L[679][4];				l_cell_reg[687] = inform_L[687][4];				l_cell_reg[688] = inform_L[688][4];				l_cell_reg[689] = inform_L[696][4];				l_cell_reg[690] = inform_L[689][4];				l_cell_reg[691] = inform_L[697][4];				l_cell_reg[692] = inform_L[690][4];				l_cell_reg[693] = inform_L[698][4];				l_cell_reg[694] = inform_L[691][4];				l_cell_reg[695] = inform_L[699][4];				l_cell_reg[696] = inform_L[692][4];				l_cell_reg[697] = inform_L[700][4];				l_cell_reg[698] = inform_L[693][4];				l_cell_reg[699] = inform_L[701][4];				l_cell_reg[700] = inform_L[694][4];				l_cell_reg[701] = inform_L[702][4];				l_cell_reg[702] = inform_L[695][4];				l_cell_reg[703] = inform_L[703][4];				l_cell_reg[704] = inform_L[704][4];				l_cell_reg[705] = inform_L[712][4];				l_cell_reg[706] = inform_L[705][4];				l_cell_reg[707] = inform_L[713][4];				l_cell_reg[708] = inform_L[706][4];				l_cell_reg[709] = inform_L[714][4];				l_cell_reg[710] = inform_L[707][4];				l_cell_reg[711] = inform_L[715][4];				l_cell_reg[712] = inform_L[708][4];				l_cell_reg[713] = inform_L[716][4];				l_cell_reg[714] = inform_L[709][4];				l_cell_reg[715] = inform_L[717][4];				l_cell_reg[716] = inform_L[710][4];				l_cell_reg[717] = inform_L[718][4];				l_cell_reg[718] = inform_L[711][4];				l_cell_reg[719] = inform_L[719][4];				l_cell_reg[720] = inform_L[720][4];				l_cell_reg[721] = inform_L[728][4];				l_cell_reg[722] = inform_L[721][4];				l_cell_reg[723] = inform_L[729][4];				l_cell_reg[724] = inform_L[722][4];				l_cell_reg[725] = inform_L[730][4];				l_cell_reg[726] = inform_L[723][4];				l_cell_reg[727] = inform_L[731][4];				l_cell_reg[728] = inform_L[724][4];				l_cell_reg[729] = inform_L[732][4];				l_cell_reg[730] = inform_L[725][4];				l_cell_reg[731] = inform_L[733][4];				l_cell_reg[732] = inform_L[726][4];				l_cell_reg[733] = inform_L[734][4];				l_cell_reg[734] = inform_L[727][4];				l_cell_reg[735] = inform_L[735][4];				l_cell_reg[736] = inform_L[736][4];				l_cell_reg[737] = inform_L[744][4];				l_cell_reg[738] = inform_L[737][4];				l_cell_reg[739] = inform_L[745][4];				l_cell_reg[740] = inform_L[738][4];				l_cell_reg[741] = inform_L[746][4];				l_cell_reg[742] = inform_L[739][4];				l_cell_reg[743] = inform_L[747][4];				l_cell_reg[744] = inform_L[740][4];				l_cell_reg[745] = inform_L[748][4];				l_cell_reg[746] = inform_L[741][4];				l_cell_reg[747] = inform_L[749][4];				l_cell_reg[748] = inform_L[742][4];				l_cell_reg[749] = inform_L[750][4];				l_cell_reg[750] = inform_L[743][4];				l_cell_reg[751] = inform_L[751][4];				l_cell_reg[752] = inform_L[752][4];				l_cell_reg[753] = inform_L[760][4];				l_cell_reg[754] = inform_L[753][4];				l_cell_reg[755] = inform_L[761][4];				l_cell_reg[756] = inform_L[754][4];				l_cell_reg[757] = inform_L[762][4];				l_cell_reg[758] = inform_L[755][4];				l_cell_reg[759] = inform_L[763][4];				l_cell_reg[760] = inform_L[756][4];				l_cell_reg[761] = inform_L[764][4];				l_cell_reg[762] = inform_L[757][4];				l_cell_reg[763] = inform_L[765][4];				l_cell_reg[764] = inform_L[758][4];				l_cell_reg[765] = inform_L[766][4];				l_cell_reg[766] = inform_L[759][4];				l_cell_reg[767] = inform_L[767][4];				l_cell_reg[768] = inform_L[768][4];				l_cell_reg[769] = inform_L[776][4];				l_cell_reg[770] = inform_L[769][4];				l_cell_reg[771] = inform_L[777][4];				l_cell_reg[772] = inform_L[770][4];				l_cell_reg[773] = inform_L[778][4];				l_cell_reg[774] = inform_L[771][4];				l_cell_reg[775] = inform_L[779][4];				l_cell_reg[776] = inform_L[772][4];				l_cell_reg[777] = inform_L[780][4];				l_cell_reg[778] = inform_L[773][4];				l_cell_reg[779] = inform_L[781][4];				l_cell_reg[780] = inform_L[774][4];				l_cell_reg[781] = inform_L[782][4];				l_cell_reg[782] = inform_L[775][4];				l_cell_reg[783] = inform_L[783][4];				l_cell_reg[784] = inform_L[784][4];				l_cell_reg[785] = inform_L[792][4];				l_cell_reg[786] = inform_L[785][4];				l_cell_reg[787] = inform_L[793][4];				l_cell_reg[788] = inform_L[786][4];				l_cell_reg[789] = inform_L[794][4];				l_cell_reg[790] = inform_L[787][4];				l_cell_reg[791] = inform_L[795][4];				l_cell_reg[792] = inform_L[788][4];				l_cell_reg[793] = inform_L[796][4];				l_cell_reg[794] = inform_L[789][4];				l_cell_reg[795] = inform_L[797][4];				l_cell_reg[796] = inform_L[790][4];				l_cell_reg[797] = inform_L[798][4];				l_cell_reg[798] = inform_L[791][4];				l_cell_reg[799] = inform_L[799][4];				l_cell_reg[800] = inform_L[800][4];				l_cell_reg[801] = inform_L[808][4];				l_cell_reg[802] = inform_L[801][4];				l_cell_reg[803] = inform_L[809][4];				l_cell_reg[804] = inform_L[802][4];				l_cell_reg[805] = inform_L[810][4];				l_cell_reg[806] = inform_L[803][4];				l_cell_reg[807] = inform_L[811][4];				l_cell_reg[808] = inform_L[804][4];				l_cell_reg[809] = inform_L[812][4];				l_cell_reg[810] = inform_L[805][4];				l_cell_reg[811] = inform_L[813][4];				l_cell_reg[812] = inform_L[806][4];				l_cell_reg[813] = inform_L[814][4];				l_cell_reg[814] = inform_L[807][4];				l_cell_reg[815] = inform_L[815][4];				l_cell_reg[816] = inform_L[816][4];				l_cell_reg[817] = inform_L[824][4];				l_cell_reg[818] = inform_L[817][4];				l_cell_reg[819] = inform_L[825][4];				l_cell_reg[820] = inform_L[818][4];				l_cell_reg[821] = inform_L[826][4];				l_cell_reg[822] = inform_L[819][4];				l_cell_reg[823] = inform_L[827][4];				l_cell_reg[824] = inform_L[820][4];				l_cell_reg[825] = inform_L[828][4];				l_cell_reg[826] = inform_L[821][4];				l_cell_reg[827] = inform_L[829][4];				l_cell_reg[828] = inform_L[822][4];				l_cell_reg[829] = inform_L[830][4];				l_cell_reg[830] = inform_L[823][4];				l_cell_reg[831] = inform_L[831][4];				l_cell_reg[832] = inform_L[832][4];				l_cell_reg[833] = inform_L[840][4];				l_cell_reg[834] = inform_L[833][4];				l_cell_reg[835] = inform_L[841][4];				l_cell_reg[836] = inform_L[834][4];				l_cell_reg[837] = inform_L[842][4];				l_cell_reg[838] = inform_L[835][4];				l_cell_reg[839] = inform_L[843][4];				l_cell_reg[840] = inform_L[836][4];				l_cell_reg[841] = inform_L[844][4];				l_cell_reg[842] = inform_L[837][4];				l_cell_reg[843] = inform_L[845][4];				l_cell_reg[844] = inform_L[838][4];				l_cell_reg[845] = inform_L[846][4];				l_cell_reg[846] = inform_L[839][4];				l_cell_reg[847] = inform_L[847][4];				l_cell_reg[848] = inform_L[848][4];				l_cell_reg[849] = inform_L[856][4];				l_cell_reg[850] = inform_L[849][4];				l_cell_reg[851] = inform_L[857][4];				l_cell_reg[852] = inform_L[850][4];				l_cell_reg[853] = inform_L[858][4];				l_cell_reg[854] = inform_L[851][4];				l_cell_reg[855] = inform_L[859][4];				l_cell_reg[856] = inform_L[852][4];				l_cell_reg[857] = inform_L[860][4];				l_cell_reg[858] = inform_L[853][4];				l_cell_reg[859] = inform_L[861][4];				l_cell_reg[860] = inform_L[854][4];				l_cell_reg[861] = inform_L[862][4];				l_cell_reg[862] = inform_L[855][4];				l_cell_reg[863] = inform_L[863][4];				l_cell_reg[864] = inform_L[864][4];				l_cell_reg[865] = inform_L[872][4];				l_cell_reg[866] = inform_L[865][4];				l_cell_reg[867] = inform_L[873][4];				l_cell_reg[868] = inform_L[866][4];				l_cell_reg[869] = inform_L[874][4];				l_cell_reg[870] = inform_L[867][4];				l_cell_reg[871] = inform_L[875][4];				l_cell_reg[872] = inform_L[868][4];				l_cell_reg[873] = inform_L[876][4];				l_cell_reg[874] = inform_L[869][4];				l_cell_reg[875] = inform_L[877][4];				l_cell_reg[876] = inform_L[870][4];				l_cell_reg[877] = inform_L[878][4];				l_cell_reg[878] = inform_L[871][4];				l_cell_reg[879] = inform_L[879][4];				l_cell_reg[880] = inform_L[880][4];				l_cell_reg[881] = inform_L[888][4];				l_cell_reg[882] = inform_L[881][4];				l_cell_reg[883] = inform_L[889][4];				l_cell_reg[884] = inform_L[882][4];				l_cell_reg[885] = inform_L[890][4];				l_cell_reg[886] = inform_L[883][4];				l_cell_reg[887] = inform_L[891][4];				l_cell_reg[888] = inform_L[884][4];				l_cell_reg[889] = inform_L[892][4];				l_cell_reg[890] = inform_L[885][4];				l_cell_reg[891] = inform_L[893][4];				l_cell_reg[892] = inform_L[886][4];				l_cell_reg[893] = inform_L[894][4];				l_cell_reg[894] = inform_L[887][4];				l_cell_reg[895] = inform_L[895][4];				l_cell_reg[896] = inform_L[896][4];				l_cell_reg[897] = inform_L[904][4];				l_cell_reg[898] = inform_L[897][4];				l_cell_reg[899] = inform_L[905][4];				l_cell_reg[900] = inform_L[898][4];				l_cell_reg[901] = inform_L[906][4];				l_cell_reg[902] = inform_L[899][4];				l_cell_reg[903] = inform_L[907][4];				l_cell_reg[904] = inform_L[900][4];				l_cell_reg[905] = inform_L[908][4];				l_cell_reg[906] = inform_L[901][4];				l_cell_reg[907] = inform_L[909][4];				l_cell_reg[908] = inform_L[902][4];				l_cell_reg[909] = inform_L[910][4];				l_cell_reg[910] = inform_L[903][4];				l_cell_reg[911] = inform_L[911][4];				l_cell_reg[912] = inform_L[912][4];				l_cell_reg[913] = inform_L[920][4];				l_cell_reg[914] = inform_L[913][4];				l_cell_reg[915] = inform_L[921][4];				l_cell_reg[916] = inform_L[914][4];				l_cell_reg[917] = inform_L[922][4];				l_cell_reg[918] = inform_L[915][4];				l_cell_reg[919] = inform_L[923][4];				l_cell_reg[920] = inform_L[916][4];				l_cell_reg[921] = inform_L[924][4];				l_cell_reg[922] = inform_L[917][4];				l_cell_reg[923] = inform_L[925][4];				l_cell_reg[924] = inform_L[918][4];				l_cell_reg[925] = inform_L[926][4];				l_cell_reg[926] = inform_L[919][4];				l_cell_reg[927] = inform_L[927][4];				l_cell_reg[928] = inform_L[928][4];				l_cell_reg[929] = inform_L[936][4];				l_cell_reg[930] = inform_L[929][4];				l_cell_reg[931] = inform_L[937][4];				l_cell_reg[932] = inform_L[930][4];				l_cell_reg[933] = inform_L[938][4];				l_cell_reg[934] = inform_L[931][4];				l_cell_reg[935] = inform_L[939][4];				l_cell_reg[936] = inform_L[932][4];				l_cell_reg[937] = inform_L[940][4];				l_cell_reg[938] = inform_L[933][4];				l_cell_reg[939] = inform_L[941][4];				l_cell_reg[940] = inform_L[934][4];				l_cell_reg[941] = inform_L[942][4];				l_cell_reg[942] = inform_L[935][4];				l_cell_reg[943] = inform_L[943][4];				l_cell_reg[944] = inform_L[944][4];				l_cell_reg[945] = inform_L[952][4];				l_cell_reg[946] = inform_L[945][4];				l_cell_reg[947] = inform_L[953][4];				l_cell_reg[948] = inform_L[946][4];				l_cell_reg[949] = inform_L[954][4];				l_cell_reg[950] = inform_L[947][4];				l_cell_reg[951] = inform_L[955][4];				l_cell_reg[952] = inform_L[948][4];				l_cell_reg[953] = inform_L[956][4];				l_cell_reg[954] = inform_L[949][4];				l_cell_reg[955] = inform_L[957][4];				l_cell_reg[956] = inform_L[950][4];				l_cell_reg[957] = inform_L[958][4];				l_cell_reg[958] = inform_L[951][4];				l_cell_reg[959] = inform_L[959][4];				l_cell_reg[960] = inform_L[960][4];				l_cell_reg[961] = inform_L[968][4];				l_cell_reg[962] = inform_L[961][4];				l_cell_reg[963] = inform_L[969][4];				l_cell_reg[964] = inform_L[962][4];				l_cell_reg[965] = inform_L[970][4];				l_cell_reg[966] = inform_L[963][4];				l_cell_reg[967] = inform_L[971][4];				l_cell_reg[968] = inform_L[964][4];				l_cell_reg[969] = inform_L[972][4];				l_cell_reg[970] = inform_L[965][4];				l_cell_reg[971] = inform_L[973][4];				l_cell_reg[972] = inform_L[966][4];				l_cell_reg[973] = inform_L[974][4];				l_cell_reg[974] = inform_L[967][4];				l_cell_reg[975] = inform_L[975][4];				l_cell_reg[976] = inform_L[976][4];				l_cell_reg[977] = inform_L[984][4];				l_cell_reg[978] = inform_L[977][4];				l_cell_reg[979] = inform_L[985][4];				l_cell_reg[980] = inform_L[978][4];				l_cell_reg[981] = inform_L[986][4];				l_cell_reg[982] = inform_L[979][4];				l_cell_reg[983] = inform_L[987][4];				l_cell_reg[984] = inform_L[980][4];				l_cell_reg[985] = inform_L[988][4];				l_cell_reg[986] = inform_L[981][4];				l_cell_reg[987] = inform_L[989][4];				l_cell_reg[988] = inform_L[982][4];				l_cell_reg[989] = inform_L[990][4];				l_cell_reg[990] = inform_L[983][4];				l_cell_reg[991] = inform_L[991][4];				l_cell_reg[992] = inform_L[992][4];				l_cell_reg[993] = inform_L[1000][4];				l_cell_reg[994] = inform_L[993][4];				l_cell_reg[995] = inform_L[1001][4];				l_cell_reg[996] = inform_L[994][4];				l_cell_reg[997] = inform_L[1002][4];				l_cell_reg[998] = inform_L[995][4];				l_cell_reg[999] = inform_L[1003][4];				l_cell_reg[1000] = inform_L[996][4];				l_cell_reg[1001] = inform_L[1004][4];				l_cell_reg[1002] = inform_L[997][4];				l_cell_reg[1003] = inform_L[1005][4];				l_cell_reg[1004] = inform_L[998][4];				l_cell_reg[1005] = inform_L[1006][4];				l_cell_reg[1006] = inform_L[999][4];				l_cell_reg[1007] = inform_L[1007][4];				l_cell_reg[1008] = inform_L[1008][4];				l_cell_reg[1009] = inform_L[1016][4];				l_cell_reg[1010] = inform_L[1009][4];				l_cell_reg[1011] = inform_L[1017][4];				l_cell_reg[1012] = inform_L[1010][4];				l_cell_reg[1013] = inform_L[1018][4];				l_cell_reg[1014] = inform_L[1011][4];				l_cell_reg[1015] = inform_L[1019][4];				l_cell_reg[1016] = inform_L[1012][4];				l_cell_reg[1017] = inform_L[1020][4];				l_cell_reg[1018] = inform_L[1013][4];				l_cell_reg[1019] = inform_L[1021][4];				l_cell_reg[1020] = inform_L[1014][4];				l_cell_reg[1021] = inform_L[1022][4];				l_cell_reg[1022] = inform_L[1015][4];				l_cell_reg[1023] = inform_L[1023][4];			end
			5:			begin				r_cell_reg[0] = inform_R[0][4];				r_cell_reg[1] = inform_R[16][4];				r_cell_reg[2] = inform_R[1][4];				r_cell_reg[3] = inform_R[17][4];				r_cell_reg[4] = inform_R[2][4];				r_cell_reg[5] = inform_R[18][4];				r_cell_reg[6] = inform_R[3][4];				r_cell_reg[7] = inform_R[19][4];				r_cell_reg[8] = inform_R[4][4];				r_cell_reg[9] = inform_R[20][4];				r_cell_reg[10] = inform_R[5][4];				r_cell_reg[11] = inform_R[21][4];				r_cell_reg[12] = inform_R[6][4];				r_cell_reg[13] = inform_R[22][4];				r_cell_reg[14] = inform_R[7][4];				r_cell_reg[15] = inform_R[23][4];				r_cell_reg[16] = inform_R[8][4];				r_cell_reg[17] = inform_R[24][4];				r_cell_reg[18] = inform_R[9][4];				r_cell_reg[19] = inform_R[25][4];				r_cell_reg[20] = inform_R[10][4];				r_cell_reg[21] = inform_R[26][4];				r_cell_reg[22] = inform_R[11][4];				r_cell_reg[23] = inform_R[27][4];				r_cell_reg[24] = inform_R[12][4];				r_cell_reg[25] = inform_R[28][4];				r_cell_reg[26] = inform_R[13][4];				r_cell_reg[27] = inform_R[29][4];				r_cell_reg[28] = inform_R[14][4];				r_cell_reg[29] = inform_R[30][4];				r_cell_reg[30] = inform_R[15][4];				r_cell_reg[31] = inform_R[31][4];				r_cell_reg[32] = inform_R[32][4];				r_cell_reg[33] = inform_R[48][4];				r_cell_reg[34] = inform_R[33][4];				r_cell_reg[35] = inform_R[49][4];				r_cell_reg[36] = inform_R[34][4];				r_cell_reg[37] = inform_R[50][4];				r_cell_reg[38] = inform_R[35][4];				r_cell_reg[39] = inform_R[51][4];				r_cell_reg[40] = inform_R[36][4];				r_cell_reg[41] = inform_R[52][4];				r_cell_reg[42] = inform_R[37][4];				r_cell_reg[43] = inform_R[53][4];				r_cell_reg[44] = inform_R[38][4];				r_cell_reg[45] = inform_R[54][4];				r_cell_reg[46] = inform_R[39][4];				r_cell_reg[47] = inform_R[55][4];				r_cell_reg[48] = inform_R[40][4];				r_cell_reg[49] = inform_R[56][4];				r_cell_reg[50] = inform_R[41][4];				r_cell_reg[51] = inform_R[57][4];				r_cell_reg[52] = inform_R[42][4];				r_cell_reg[53] = inform_R[58][4];				r_cell_reg[54] = inform_R[43][4];				r_cell_reg[55] = inform_R[59][4];				r_cell_reg[56] = inform_R[44][4];				r_cell_reg[57] = inform_R[60][4];				r_cell_reg[58] = inform_R[45][4];				r_cell_reg[59] = inform_R[61][4];				r_cell_reg[60] = inform_R[46][4];				r_cell_reg[61] = inform_R[62][4];				r_cell_reg[62] = inform_R[47][4];				r_cell_reg[63] = inform_R[63][4];				r_cell_reg[64] = inform_R[64][4];				r_cell_reg[65] = inform_R[80][4];				r_cell_reg[66] = inform_R[65][4];				r_cell_reg[67] = inform_R[81][4];				r_cell_reg[68] = inform_R[66][4];				r_cell_reg[69] = inform_R[82][4];				r_cell_reg[70] = inform_R[67][4];				r_cell_reg[71] = inform_R[83][4];				r_cell_reg[72] = inform_R[68][4];				r_cell_reg[73] = inform_R[84][4];				r_cell_reg[74] = inform_R[69][4];				r_cell_reg[75] = inform_R[85][4];				r_cell_reg[76] = inform_R[70][4];				r_cell_reg[77] = inform_R[86][4];				r_cell_reg[78] = inform_R[71][4];				r_cell_reg[79] = inform_R[87][4];				r_cell_reg[80] = inform_R[72][4];				r_cell_reg[81] = inform_R[88][4];				r_cell_reg[82] = inform_R[73][4];				r_cell_reg[83] = inform_R[89][4];				r_cell_reg[84] = inform_R[74][4];				r_cell_reg[85] = inform_R[90][4];				r_cell_reg[86] = inform_R[75][4];				r_cell_reg[87] = inform_R[91][4];				r_cell_reg[88] = inform_R[76][4];				r_cell_reg[89] = inform_R[92][4];				r_cell_reg[90] = inform_R[77][4];				r_cell_reg[91] = inform_R[93][4];				r_cell_reg[92] = inform_R[78][4];				r_cell_reg[93] = inform_R[94][4];				r_cell_reg[94] = inform_R[79][4];				r_cell_reg[95] = inform_R[95][4];				r_cell_reg[96] = inform_R[96][4];				r_cell_reg[97] = inform_R[112][4];				r_cell_reg[98] = inform_R[97][4];				r_cell_reg[99] = inform_R[113][4];				r_cell_reg[100] = inform_R[98][4];				r_cell_reg[101] = inform_R[114][4];				r_cell_reg[102] = inform_R[99][4];				r_cell_reg[103] = inform_R[115][4];				r_cell_reg[104] = inform_R[100][4];				r_cell_reg[105] = inform_R[116][4];				r_cell_reg[106] = inform_R[101][4];				r_cell_reg[107] = inform_R[117][4];				r_cell_reg[108] = inform_R[102][4];				r_cell_reg[109] = inform_R[118][4];				r_cell_reg[110] = inform_R[103][4];				r_cell_reg[111] = inform_R[119][4];				r_cell_reg[112] = inform_R[104][4];				r_cell_reg[113] = inform_R[120][4];				r_cell_reg[114] = inform_R[105][4];				r_cell_reg[115] = inform_R[121][4];				r_cell_reg[116] = inform_R[106][4];				r_cell_reg[117] = inform_R[122][4];				r_cell_reg[118] = inform_R[107][4];				r_cell_reg[119] = inform_R[123][4];				r_cell_reg[120] = inform_R[108][4];				r_cell_reg[121] = inform_R[124][4];				r_cell_reg[122] = inform_R[109][4];				r_cell_reg[123] = inform_R[125][4];				r_cell_reg[124] = inform_R[110][4];				r_cell_reg[125] = inform_R[126][4];				r_cell_reg[126] = inform_R[111][4];				r_cell_reg[127] = inform_R[127][4];				r_cell_reg[128] = inform_R[128][4];				r_cell_reg[129] = inform_R[144][4];				r_cell_reg[130] = inform_R[129][4];				r_cell_reg[131] = inform_R[145][4];				r_cell_reg[132] = inform_R[130][4];				r_cell_reg[133] = inform_R[146][4];				r_cell_reg[134] = inform_R[131][4];				r_cell_reg[135] = inform_R[147][4];				r_cell_reg[136] = inform_R[132][4];				r_cell_reg[137] = inform_R[148][4];				r_cell_reg[138] = inform_R[133][4];				r_cell_reg[139] = inform_R[149][4];				r_cell_reg[140] = inform_R[134][4];				r_cell_reg[141] = inform_R[150][4];				r_cell_reg[142] = inform_R[135][4];				r_cell_reg[143] = inform_R[151][4];				r_cell_reg[144] = inform_R[136][4];				r_cell_reg[145] = inform_R[152][4];				r_cell_reg[146] = inform_R[137][4];				r_cell_reg[147] = inform_R[153][4];				r_cell_reg[148] = inform_R[138][4];				r_cell_reg[149] = inform_R[154][4];				r_cell_reg[150] = inform_R[139][4];				r_cell_reg[151] = inform_R[155][4];				r_cell_reg[152] = inform_R[140][4];				r_cell_reg[153] = inform_R[156][4];				r_cell_reg[154] = inform_R[141][4];				r_cell_reg[155] = inform_R[157][4];				r_cell_reg[156] = inform_R[142][4];				r_cell_reg[157] = inform_R[158][4];				r_cell_reg[158] = inform_R[143][4];				r_cell_reg[159] = inform_R[159][4];				r_cell_reg[160] = inform_R[160][4];				r_cell_reg[161] = inform_R[176][4];				r_cell_reg[162] = inform_R[161][4];				r_cell_reg[163] = inform_R[177][4];				r_cell_reg[164] = inform_R[162][4];				r_cell_reg[165] = inform_R[178][4];				r_cell_reg[166] = inform_R[163][4];				r_cell_reg[167] = inform_R[179][4];				r_cell_reg[168] = inform_R[164][4];				r_cell_reg[169] = inform_R[180][4];				r_cell_reg[170] = inform_R[165][4];				r_cell_reg[171] = inform_R[181][4];				r_cell_reg[172] = inform_R[166][4];				r_cell_reg[173] = inform_R[182][4];				r_cell_reg[174] = inform_R[167][4];				r_cell_reg[175] = inform_R[183][4];				r_cell_reg[176] = inform_R[168][4];				r_cell_reg[177] = inform_R[184][4];				r_cell_reg[178] = inform_R[169][4];				r_cell_reg[179] = inform_R[185][4];				r_cell_reg[180] = inform_R[170][4];				r_cell_reg[181] = inform_R[186][4];				r_cell_reg[182] = inform_R[171][4];				r_cell_reg[183] = inform_R[187][4];				r_cell_reg[184] = inform_R[172][4];				r_cell_reg[185] = inform_R[188][4];				r_cell_reg[186] = inform_R[173][4];				r_cell_reg[187] = inform_R[189][4];				r_cell_reg[188] = inform_R[174][4];				r_cell_reg[189] = inform_R[190][4];				r_cell_reg[190] = inform_R[175][4];				r_cell_reg[191] = inform_R[191][4];				r_cell_reg[192] = inform_R[192][4];				r_cell_reg[193] = inform_R[208][4];				r_cell_reg[194] = inform_R[193][4];				r_cell_reg[195] = inform_R[209][4];				r_cell_reg[196] = inform_R[194][4];				r_cell_reg[197] = inform_R[210][4];				r_cell_reg[198] = inform_R[195][4];				r_cell_reg[199] = inform_R[211][4];				r_cell_reg[200] = inform_R[196][4];				r_cell_reg[201] = inform_R[212][4];				r_cell_reg[202] = inform_R[197][4];				r_cell_reg[203] = inform_R[213][4];				r_cell_reg[204] = inform_R[198][4];				r_cell_reg[205] = inform_R[214][4];				r_cell_reg[206] = inform_R[199][4];				r_cell_reg[207] = inform_R[215][4];				r_cell_reg[208] = inform_R[200][4];				r_cell_reg[209] = inform_R[216][4];				r_cell_reg[210] = inform_R[201][4];				r_cell_reg[211] = inform_R[217][4];				r_cell_reg[212] = inform_R[202][4];				r_cell_reg[213] = inform_R[218][4];				r_cell_reg[214] = inform_R[203][4];				r_cell_reg[215] = inform_R[219][4];				r_cell_reg[216] = inform_R[204][4];				r_cell_reg[217] = inform_R[220][4];				r_cell_reg[218] = inform_R[205][4];				r_cell_reg[219] = inform_R[221][4];				r_cell_reg[220] = inform_R[206][4];				r_cell_reg[221] = inform_R[222][4];				r_cell_reg[222] = inform_R[207][4];				r_cell_reg[223] = inform_R[223][4];				r_cell_reg[224] = inform_R[224][4];				r_cell_reg[225] = inform_R[240][4];				r_cell_reg[226] = inform_R[225][4];				r_cell_reg[227] = inform_R[241][4];				r_cell_reg[228] = inform_R[226][4];				r_cell_reg[229] = inform_R[242][4];				r_cell_reg[230] = inform_R[227][4];				r_cell_reg[231] = inform_R[243][4];				r_cell_reg[232] = inform_R[228][4];				r_cell_reg[233] = inform_R[244][4];				r_cell_reg[234] = inform_R[229][4];				r_cell_reg[235] = inform_R[245][4];				r_cell_reg[236] = inform_R[230][4];				r_cell_reg[237] = inform_R[246][4];				r_cell_reg[238] = inform_R[231][4];				r_cell_reg[239] = inform_R[247][4];				r_cell_reg[240] = inform_R[232][4];				r_cell_reg[241] = inform_R[248][4];				r_cell_reg[242] = inform_R[233][4];				r_cell_reg[243] = inform_R[249][4];				r_cell_reg[244] = inform_R[234][4];				r_cell_reg[245] = inform_R[250][4];				r_cell_reg[246] = inform_R[235][4];				r_cell_reg[247] = inform_R[251][4];				r_cell_reg[248] = inform_R[236][4];				r_cell_reg[249] = inform_R[252][4];				r_cell_reg[250] = inform_R[237][4];				r_cell_reg[251] = inform_R[253][4];				r_cell_reg[252] = inform_R[238][4];				r_cell_reg[253] = inform_R[254][4];				r_cell_reg[254] = inform_R[239][4];				r_cell_reg[255] = inform_R[255][4];				r_cell_reg[256] = inform_R[256][4];				r_cell_reg[257] = inform_R[272][4];				r_cell_reg[258] = inform_R[257][4];				r_cell_reg[259] = inform_R[273][4];				r_cell_reg[260] = inform_R[258][4];				r_cell_reg[261] = inform_R[274][4];				r_cell_reg[262] = inform_R[259][4];				r_cell_reg[263] = inform_R[275][4];				r_cell_reg[264] = inform_R[260][4];				r_cell_reg[265] = inform_R[276][4];				r_cell_reg[266] = inform_R[261][4];				r_cell_reg[267] = inform_R[277][4];				r_cell_reg[268] = inform_R[262][4];				r_cell_reg[269] = inform_R[278][4];				r_cell_reg[270] = inform_R[263][4];				r_cell_reg[271] = inform_R[279][4];				r_cell_reg[272] = inform_R[264][4];				r_cell_reg[273] = inform_R[280][4];				r_cell_reg[274] = inform_R[265][4];				r_cell_reg[275] = inform_R[281][4];				r_cell_reg[276] = inform_R[266][4];				r_cell_reg[277] = inform_R[282][4];				r_cell_reg[278] = inform_R[267][4];				r_cell_reg[279] = inform_R[283][4];				r_cell_reg[280] = inform_R[268][4];				r_cell_reg[281] = inform_R[284][4];				r_cell_reg[282] = inform_R[269][4];				r_cell_reg[283] = inform_R[285][4];				r_cell_reg[284] = inform_R[270][4];				r_cell_reg[285] = inform_R[286][4];				r_cell_reg[286] = inform_R[271][4];				r_cell_reg[287] = inform_R[287][4];				r_cell_reg[288] = inform_R[288][4];				r_cell_reg[289] = inform_R[304][4];				r_cell_reg[290] = inform_R[289][4];				r_cell_reg[291] = inform_R[305][4];				r_cell_reg[292] = inform_R[290][4];				r_cell_reg[293] = inform_R[306][4];				r_cell_reg[294] = inform_R[291][4];				r_cell_reg[295] = inform_R[307][4];				r_cell_reg[296] = inform_R[292][4];				r_cell_reg[297] = inform_R[308][4];				r_cell_reg[298] = inform_R[293][4];				r_cell_reg[299] = inform_R[309][4];				r_cell_reg[300] = inform_R[294][4];				r_cell_reg[301] = inform_R[310][4];				r_cell_reg[302] = inform_R[295][4];				r_cell_reg[303] = inform_R[311][4];				r_cell_reg[304] = inform_R[296][4];				r_cell_reg[305] = inform_R[312][4];				r_cell_reg[306] = inform_R[297][4];				r_cell_reg[307] = inform_R[313][4];				r_cell_reg[308] = inform_R[298][4];				r_cell_reg[309] = inform_R[314][4];				r_cell_reg[310] = inform_R[299][4];				r_cell_reg[311] = inform_R[315][4];				r_cell_reg[312] = inform_R[300][4];				r_cell_reg[313] = inform_R[316][4];				r_cell_reg[314] = inform_R[301][4];				r_cell_reg[315] = inform_R[317][4];				r_cell_reg[316] = inform_R[302][4];				r_cell_reg[317] = inform_R[318][4];				r_cell_reg[318] = inform_R[303][4];				r_cell_reg[319] = inform_R[319][4];				r_cell_reg[320] = inform_R[320][4];				r_cell_reg[321] = inform_R[336][4];				r_cell_reg[322] = inform_R[321][4];				r_cell_reg[323] = inform_R[337][4];				r_cell_reg[324] = inform_R[322][4];				r_cell_reg[325] = inform_R[338][4];				r_cell_reg[326] = inform_R[323][4];				r_cell_reg[327] = inform_R[339][4];				r_cell_reg[328] = inform_R[324][4];				r_cell_reg[329] = inform_R[340][4];				r_cell_reg[330] = inform_R[325][4];				r_cell_reg[331] = inform_R[341][4];				r_cell_reg[332] = inform_R[326][4];				r_cell_reg[333] = inform_R[342][4];				r_cell_reg[334] = inform_R[327][4];				r_cell_reg[335] = inform_R[343][4];				r_cell_reg[336] = inform_R[328][4];				r_cell_reg[337] = inform_R[344][4];				r_cell_reg[338] = inform_R[329][4];				r_cell_reg[339] = inform_R[345][4];				r_cell_reg[340] = inform_R[330][4];				r_cell_reg[341] = inform_R[346][4];				r_cell_reg[342] = inform_R[331][4];				r_cell_reg[343] = inform_R[347][4];				r_cell_reg[344] = inform_R[332][4];				r_cell_reg[345] = inform_R[348][4];				r_cell_reg[346] = inform_R[333][4];				r_cell_reg[347] = inform_R[349][4];				r_cell_reg[348] = inform_R[334][4];				r_cell_reg[349] = inform_R[350][4];				r_cell_reg[350] = inform_R[335][4];				r_cell_reg[351] = inform_R[351][4];				r_cell_reg[352] = inform_R[352][4];				r_cell_reg[353] = inform_R[368][4];				r_cell_reg[354] = inform_R[353][4];				r_cell_reg[355] = inform_R[369][4];				r_cell_reg[356] = inform_R[354][4];				r_cell_reg[357] = inform_R[370][4];				r_cell_reg[358] = inform_R[355][4];				r_cell_reg[359] = inform_R[371][4];				r_cell_reg[360] = inform_R[356][4];				r_cell_reg[361] = inform_R[372][4];				r_cell_reg[362] = inform_R[357][4];				r_cell_reg[363] = inform_R[373][4];				r_cell_reg[364] = inform_R[358][4];				r_cell_reg[365] = inform_R[374][4];				r_cell_reg[366] = inform_R[359][4];				r_cell_reg[367] = inform_R[375][4];				r_cell_reg[368] = inform_R[360][4];				r_cell_reg[369] = inform_R[376][4];				r_cell_reg[370] = inform_R[361][4];				r_cell_reg[371] = inform_R[377][4];				r_cell_reg[372] = inform_R[362][4];				r_cell_reg[373] = inform_R[378][4];				r_cell_reg[374] = inform_R[363][4];				r_cell_reg[375] = inform_R[379][4];				r_cell_reg[376] = inform_R[364][4];				r_cell_reg[377] = inform_R[380][4];				r_cell_reg[378] = inform_R[365][4];				r_cell_reg[379] = inform_R[381][4];				r_cell_reg[380] = inform_R[366][4];				r_cell_reg[381] = inform_R[382][4];				r_cell_reg[382] = inform_R[367][4];				r_cell_reg[383] = inform_R[383][4];				r_cell_reg[384] = inform_R[384][4];				r_cell_reg[385] = inform_R[400][4];				r_cell_reg[386] = inform_R[385][4];				r_cell_reg[387] = inform_R[401][4];				r_cell_reg[388] = inform_R[386][4];				r_cell_reg[389] = inform_R[402][4];				r_cell_reg[390] = inform_R[387][4];				r_cell_reg[391] = inform_R[403][4];				r_cell_reg[392] = inform_R[388][4];				r_cell_reg[393] = inform_R[404][4];				r_cell_reg[394] = inform_R[389][4];				r_cell_reg[395] = inform_R[405][4];				r_cell_reg[396] = inform_R[390][4];				r_cell_reg[397] = inform_R[406][4];				r_cell_reg[398] = inform_R[391][4];				r_cell_reg[399] = inform_R[407][4];				r_cell_reg[400] = inform_R[392][4];				r_cell_reg[401] = inform_R[408][4];				r_cell_reg[402] = inform_R[393][4];				r_cell_reg[403] = inform_R[409][4];				r_cell_reg[404] = inform_R[394][4];				r_cell_reg[405] = inform_R[410][4];				r_cell_reg[406] = inform_R[395][4];				r_cell_reg[407] = inform_R[411][4];				r_cell_reg[408] = inform_R[396][4];				r_cell_reg[409] = inform_R[412][4];				r_cell_reg[410] = inform_R[397][4];				r_cell_reg[411] = inform_R[413][4];				r_cell_reg[412] = inform_R[398][4];				r_cell_reg[413] = inform_R[414][4];				r_cell_reg[414] = inform_R[399][4];				r_cell_reg[415] = inform_R[415][4];				r_cell_reg[416] = inform_R[416][4];				r_cell_reg[417] = inform_R[432][4];				r_cell_reg[418] = inform_R[417][4];				r_cell_reg[419] = inform_R[433][4];				r_cell_reg[420] = inform_R[418][4];				r_cell_reg[421] = inform_R[434][4];				r_cell_reg[422] = inform_R[419][4];				r_cell_reg[423] = inform_R[435][4];				r_cell_reg[424] = inform_R[420][4];				r_cell_reg[425] = inform_R[436][4];				r_cell_reg[426] = inform_R[421][4];				r_cell_reg[427] = inform_R[437][4];				r_cell_reg[428] = inform_R[422][4];				r_cell_reg[429] = inform_R[438][4];				r_cell_reg[430] = inform_R[423][4];				r_cell_reg[431] = inform_R[439][4];				r_cell_reg[432] = inform_R[424][4];				r_cell_reg[433] = inform_R[440][4];				r_cell_reg[434] = inform_R[425][4];				r_cell_reg[435] = inform_R[441][4];				r_cell_reg[436] = inform_R[426][4];				r_cell_reg[437] = inform_R[442][4];				r_cell_reg[438] = inform_R[427][4];				r_cell_reg[439] = inform_R[443][4];				r_cell_reg[440] = inform_R[428][4];				r_cell_reg[441] = inform_R[444][4];				r_cell_reg[442] = inform_R[429][4];				r_cell_reg[443] = inform_R[445][4];				r_cell_reg[444] = inform_R[430][4];				r_cell_reg[445] = inform_R[446][4];				r_cell_reg[446] = inform_R[431][4];				r_cell_reg[447] = inform_R[447][4];				r_cell_reg[448] = inform_R[448][4];				r_cell_reg[449] = inform_R[464][4];				r_cell_reg[450] = inform_R[449][4];				r_cell_reg[451] = inform_R[465][4];				r_cell_reg[452] = inform_R[450][4];				r_cell_reg[453] = inform_R[466][4];				r_cell_reg[454] = inform_R[451][4];				r_cell_reg[455] = inform_R[467][4];				r_cell_reg[456] = inform_R[452][4];				r_cell_reg[457] = inform_R[468][4];				r_cell_reg[458] = inform_R[453][4];				r_cell_reg[459] = inform_R[469][4];				r_cell_reg[460] = inform_R[454][4];				r_cell_reg[461] = inform_R[470][4];				r_cell_reg[462] = inform_R[455][4];				r_cell_reg[463] = inform_R[471][4];				r_cell_reg[464] = inform_R[456][4];				r_cell_reg[465] = inform_R[472][4];				r_cell_reg[466] = inform_R[457][4];				r_cell_reg[467] = inform_R[473][4];				r_cell_reg[468] = inform_R[458][4];				r_cell_reg[469] = inform_R[474][4];				r_cell_reg[470] = inform_R[459][4];				r_cell_reg[471] = inform_R[475][4];				r_cell_reg[472] = inform_R[460][4];				r_cell_reg[473] = inform_R[476][4];				r_cell_reg[474] = inform_R[461][4];				r_cell_reg[475] = inform_R[477][4];				r_cell_reg[476] = inform_R[462][4];				r_cell_reg[477] = inform_R[478][4];				r_cell_reg[478] = inform_R[463][4];				r_cell_reg[479] = inform_R[479][4];				r_cell_reg[480] = inform_R[480][4];				r_cell_reg[481] = inform_R[496][4];				r_cell_reg[482] = inform_R[481][4];				r_cell_reg[483] = inform_R[497][4];				r_cell_reg[484] = inform_R[482][4];				r_cell_reg[485] = inform_R[498][4];				r_cell_reg[486] = inform_R[483][4];				r_cell_reg[487] = inform_R[499][4];				r_cell_reg[488] = inform_R[484][4];				r_cell_reg[489] = inform_R[500][4];				r_cell_reg[490] = inform_R[485][4];				r_cell_reg[491] = inform_R[501][4];				r_cell_reg[492] = inform_R[486][4];				r_cell_reg[493] = inform_R[502][4];				r_cell_reg[494] = inform_R[487][4];				r_cell_reg[495] = inform_R[503][4];				r_cell_reg[496] = inform_R[488][4];				r_cell_reg[497] = inform_R[504][4];				r_cell_reg[498] = inform_R[489][4];				r_cell_reg[499] = inform_R[505][4];				r_cell_reg[500] = inform_R[490][4];				r_cell_reg[501] = inform_R[506][4];				r_cell_reg[502] = inform_R[491][4];				r_cell_reg[503] = inform_R[507][4];				r_cell_reg[504] = inform_R[492][4];				r_cell_reg[505] = inform_R[508][4];				r_cell_reg[506] = inform_R[493][4];				r_cell_reg[507] = inform_R[509][4];				r_cell_reg[508] = inform_R[494][4];				r_cell_reg[509] = inform_R[510][4];				r_cell_reg[510] = inform_R[495][4];				r_cell_reg[511] = inform_R[511][4];				r_cell_reg[512] = inform_R[512][4];				r_cell_reg[513] = inform_R[528][4];				r_cell_reg[514] = inform_R[513][4];				r_cell_reg[515] = inform_R[529][4];				r_cell_reg[516] = inform_R[514][4];				r_cell_reg[517] = inform_R[530][4];				r_cell_reg[518] = inform_R[515][4];				r_cell_reg[519] = inform_R[531][4];				r_cell_reg[520] = inform_R[516][4];				r_cell_reg[521] = inform_R[532][4];				r_cell_reg[522] = inform_R[517][4];				r_cell_reg[523] = inform_R[533][4];				r_cell_reg[524] = inform_R[518][4];				r_cell_reg[525] = inform_R[534][4];				r_cell_reg[526] = inform_R[519][4];				r_cell_reg[527] = inform_R[535][4];				r_cell_reg[528] = inform_R[520][4];				r_cell_reg[529] = inform_R[536][4];				r_cell_reg[530] = inform_R[521][4];				r_cell_reg[531] = inform_R[537][4];				r_cell_reg[532] = inform_R[522][4];				r_cell_reg[533] = inform_R[538][4];				r_cell_reg[534] = inform_R[523][4];				r_cell_reg[535] = inform_R[539][4];				r_cell_reg[536] = inform_R[524][4];				r_cell_reg[537] = inform_R[540][4];				r_cell_reg[538] = inform_R[525][4];				r_cell_reg[539] = inform_R[541][4];				r_cell_reg[540] = inform_R[526][4];				r_cell_reg[541] = inform_R[542][4];				r_cell_reg[542] = inform_R[527][4];				r_cell_reg[543] = inform_R[543][4];				r_cell_reg[544] = inform_R[544][4];				r_cell_reg[545] = inform_R[560][4];				r_cell_reg[546] = inform_R[545][4];				r_cell_reg[547] = inform_R[561][4];				r_cell_reg[548] = inform_R[546][4];				r_cell_reg[549] = inform_R[562][4];				r_cell_reg[550] = inform_R[547][4];				r_cell_reg[551] = inform_R[563][4];				r_cell_reg[552] = inform_R[548][4];				r_cell_reg[553] = inform_R[564][4];				r_cell_reg[554] = inform_R[549][4];				r_cell_reg[555] = inform_R[565][4];				r_cell_reg[556] = inform_R[550][4];				r_cell_reg[557] = inform_R[566][4];				r_cell_reg[558] = inform_R[551][4];				r_cell_reg[559] = inform_R[567][4];				r_cell_reg[560] = inform_R[552][4];				r_cell_reg[561] = inform_R[568][4];				r_cell_reg[562] = inform_R[553][4];				r_cell_reg[563] = inform_R[569][4];				r_cell_reg[564] = inform_R[554][4];				r_cell_reg[565] = inform_R[570][4];				r_cell_reg[566] = inform_R[555][4];				r_cell_reg[567] = inform_R[571][4];				r_cell_reg[568] = inform_R[556][4];				r_cell_reg[569] = inform_R[572][4];				r_cell_reg[570] = inform_R[557][4];				r_cell_reg[571] = inform_R[573][4];				r_cell_reg[572] = inform_R[558][4];				r_cell_reg[573] = inform_R[574][4];				r_cell_reg[574] = inform_R[559][4];				r_cell_reg[575] = inform_R[575][4];				r_cell_reg[576] = inform_R[576][4];				r_cell_reg[577] = inform_R[592][4];				r_cell_reg[578] = inform_R[577][4];				r_cell_reg[579] = inform_R[593][4];				r_cell_reg[580] = inform_R[578][4];				r_cell_reg[581] = inform_R[594][4];				r_cell_reg[582] = inform_R[579][4];				r_cell_reg[583] = inform_R[595][4];				r_cell_reg[584] = inform_R[580][4];				r_cell_reg[585] = inform_R[596][4];				r_cell_reg[586] = inform_R[581][4];				r_cell_reg[587] = inform_R[597][4];				r_cell_reg[588] = inform_R[582][4];				r_cell_reg[589] = inform_R[598][4];				r_cell_reg[590] = inform_R[583][4];				r_cell_reg[591] = inform_R[599][4];				r_cell_reg[592] = inform_R[584][4];				r_cell_reg[593] = inform_R[600][4];				r_cell_reg[594] = inform_R[585][4];				r_cell_reg[595] = inform_R[601][4];				r_cell_reg[596] = inform_R[586][4];				r_cell_reg[597] = inform_R[602][4];				r_cell_reg[598] = inform_R[587][4];				r_cell_reg[599] = inform_R[603][4];				r_cell_reg[600] = inform_R[588][4];				r_cell_reg[601] = inform_R[604][4];				r_cell_reg[602] = inform_R[589][4];				r_cell_reg[603] = inform_R[605][4];				r_cell_reg[604] = inform_R[590][4];				r_cell_reg[605] = inform_R[606][4];				r_cell_reg[606] = inform_R[591][4];				r_cell_reg[607] = inform_R[607][4];				r_cell_reg[608] = inform_R[608][4];				r_cell_reg[609] = inform_R[624][4];				r_cell_reg[610] = inform_R[609][4];				r_cell_reg[611] = inform_R[625][4];				r_cell_reg[612] = inform_R[610][4];				r_cell_reg[613] = inform_R[626][4];				r_cell_reg[614] = inform_R[611][4];				r_cell_reg[615] = inform_R[627][4];				r_cell_reg[616] = inform_R[612][4];				r_cell_reg[617] = inform_R[628][4];				r_cell_reg[618] = inform_R[613][4];				r_cell_reg[619] = inform_R[629][4];				r_cell_reg[620] = inform_R[614][4];				r_cell_reg[621] = inform_R[630][4];				r_cell_reg[622] = inform_R[615][4];				r_cell_reg[623] = inform_R[631][4];				r_cell_reg[624] = inform_R[616][4];				r_cell_reg[625] = inform_R[632][4];				r_cell_reg[626] = inform_R[617][4];				r_cell_reg[627] = inform_R[633][4];				r_cell_reg[628] = inform_R[618][4];				r_cell_reg[629] = inform_R[634][4];				r_cell_reg[630] = inform_R[619][4];				r_cell_reg[631] = inform_R[635][4];				r_cell_reg[632] = inform_R[620][4];				r_cell_reg[633] = inform_R[636][4];				r_cell_reg[634] = inform_R[621][4];				r_cell_reg[635] = inform_R[637][4];				r_cell_reg[636] = inform_R[622][4];				r_cell_reg[637] = inform_R[638][4];				r_cell_reg[638] = inform_R[623][4];				r_cell_reg[639] = inform_R[639][4];				r_cell_reg[640] = inform_R[640][4];				r_cell_reg[641] = inform_R[656][4];				r_cell_reg[642] = inform_R[641][4];				r_cell_reg[643] = inform_R[657][4];				r_cell_reg[644] = inform_R[642][4];				r_cell_reg[645] = inform_R[658][4];				r_cell_reg[646] = inform_R[643][4];				r_cell_reg[647] = inform_R[659][4];				r_cell_reg[648] = inform_R[644][4];				r_cell_reg[649] = inform_R[660][4];				r_cell_reg[650] = inform_R[645][4];				r_cell_reg[651] = inform_R[661][4];				r_cell_reg[652] = inform_R[646][4];				r_cell_reg[653] = inform_R[662][4];				r_cell_reg[654] = inform_R[647][4];				r_cell_reg[655] = inform_R[663][4];				r_cell_reg[656] = inform_R[648][4];				r_cell_reg[657] = inform_R[664][4];				r_cell_reg[658] = inform_R[649][4];				r_cell_reg[659] = inform_R[665][4];				r_cell_reg[660] = inform_R[650][4];				r_cell_reg[661] = inform_R[666][4];				r_cell_reg[662] = inform_R[651][4];				r_cell_reg[663] = inform_R[667][4];				r_cell_reg[664] = inform_R[652][4];				r_cell_reg[665] = inform_R[668][4];				r_cell_reg[666] = inform_R[653][4];				r_cell_reg[667] = inform_R[669][4];				r_cell_reg[668] = inform_R[654][4];				r_cell_reg[669] = inform_R[670][4];				r_cell_reg[670] = inform_R[655][4];				r_cell_reg[671] = inform_R[671][4];				r_cell_reg[672] = inform_R[672][4];				r_cell_reg[673] = inform_R[688][4];				r_cell_reg[674] = inform_R[673][4];				r_cell_reg[675] = inform_R[689][4];				r_cell_reg[676] = inform_R[674][4];				r_cell_reg[677] = inform_R[690][4];				r_cell_reg[678] = inform_R[675][4];				r_cell_reg[679] = inform_R[691][4];				r_cell_reg[680] = inform_R[676][4];				r_cell_reg[681] = inform_R[692][4];				r_cell_reg[682] = inform_R[677][4];				r_cell_reg[683] = inform_R[693][4];				r_cell_reg[684] = inform_R[678][4];				r_cell_reg[685] = inform_R[694][4];				r_cell_reg[686] = inform_R[679][4];				r_cell_reg[687] = inform_R[695][4];				r_cell_reg[688] = inform_R[680][4];				r_cell_reg[689] = inform_R[696][4];				r_cell_reg[690] = inform_R[681][4];				r_cell_reg[691] = inform_R[697][4];				r_cell_reg[692] = inform_R[682][4];				r_cell_reg[693] = inform_R[698][4];				r_cell_reg[694] = inform_R[683][4];				r_cell_reg[695] = inform_R[699][4];				r_cell_reg[696] = inform_R[684][4];				r_cell_reg[697] = inform_R[700][4];				r_cell_reg[698] = inform_R[685][4];				r_cell_reg[699] = inform_R[701][4];				r_cell_reg[700] = inform_R[686][4];				r_cell_reg[701] = inform_R[702][4];				r_cell_reg[702] = inform_R[687][4];				r_cell_reg[703] = inform_R[703][4];				r_cell_reg[704] = inform_R[704][4];				r_cell_reg[705] = inform_R[720][4];				r_cell_reg[706] = inform_R[705][4];				r_cell_reg[707] = inform_R[721][4];				r_cell_reg[708] = inform_R[706][4];				r_cell_reg[709] = inform_R[722][4];				r_cell_reg[710] = inform_R[707][4];				r_cell_reg[711] = inform_R[723][4];				r_cell_reg[712] = inform_R[708][4];				r_cell_reg[713] = inform_R[724][4];				r_cell_reg[714] = inform_R[709][4];				r_cell_reg[715] = inform_R[725][4];				r_cell_reg[716] = inform_R[710][4];				r_cell_reg[717] = inform_R[726][4];				r_cell_reg[718] = inform_R[711][4];				r_cell_reg[719] = inform_R[727][4];				r_cell_reg[720] = inform_R[712][4];				r_cell_reg[721] = inform_R[728][4];				r_cell_reg[722] = inform_R[713][4];				r_cell_reg[723] = inform_R[729][4];				r_cell_reg[724] = inform_R[714][4];				r_cell_reg[725] = inform_R[730][4];				r_cell_reg[726] = inform_R[715][4];				r_cell_reg[727] = inform_R[731][4];				r_cell_reg[728] = inform_R[716][4];				r_cell_reg[729] = inform_R[732][4];				r_cell_reg[730] = inform_R[717][4];				r_cell_reg[731] = inform_R[733][4];				r_cell_reg[732] = inform_R[718][4];				r_cell_reg[733] = inform_R[734][4];				r_cell_reg[734] = inform_R[719][4];				r_cell_reg[735] = inform_R[735][4];				r_cell_reg[736] = inform_R[736][4];				r_cell_reg[737] = inform_R[752][4];				r_cell_reg[738] = inform_R[737][4];				r_cell_reg[739] = inform_R[753][4];				r_cell_reg[740] = inform_R[738][4];				r_cell_reg[741] = inform_R[754][4];				r_cell_reg[742] = inform_R[739][4];				r_cell_reg[743] = inform_R[755][4];				r_cell_reg[744] = inform_R[740][4];				r_cell_reg[745] = inform_R[756][4];				r_cell_reg[746] = inform_R[741][4];				r_cell_reg[747] = inform_R[757][4];				r_cell_reg[748] = inform_R[742][4];				r_cell_reg[749] = inform_R[758][4];				r_cell_reg[750] = inform_R[743][4];				r_cell_reg[751] = inform_R[759][4];				r_cell_reg[752] = inform_R[744][4];				r_cell_reg[753] = inform_R[760][4];				r_cell_reg[754] = inform_R[745][4];				r_cell_reg[755] = inform_R[761][4];				r_cell_reg[756] = inform_R[746][4];				r_cell_reg[757] = inform_R[762][4];				r_cell_reg[758] = inform_R[747][4];				r_cell_reg[759] = inform_R[763][4];				r_cell_reg[760] = inform_R[748][4];				r_cell_reg[761] = inform_R[764][4];				r_cell_reg[762] = inform_R[749][4];				r_cell_reg[763] = inform_R[765][4];				r_cell_reg[764] = inform_R[750][4];				r_cell_reg[765] = inform_R[766][4];				r_cell_reg[766] = inform_R[751][4];				r_cell_reg[767] = inform_R[767][4];				r_cell_reg[768] = inform_R[768][4];				r_cell_reg[769] = inform_R[784][4];				r_cell_reg[770] = inform_R[769][4];				r_cell_reg[771] = inform_R[785][4];				r_cell_reg[772] = inform_R[770][4];				r_cell_reg[773] = inform_R[786][4];				r_cell_reg[774] = inform_R[771][4];				r_cell_reg[775] = inform_R[787][4];				r_cell_reg[776] = inform_R[772][4];				r_cell_reg[777] = inform_R[788][4];				r_cell_reg[778] = inform_R[773][4];				r_cell_reg[779] = inform_R[789][4];				r_cell_reg[780] = inform_R[774][4];				r_cell_reg[781] = inform_R[790][4];				r_cell_reg[782] = inform_R[775][4];				r_cell_reg[783] = inform_R[791][4];				r_cell_reg[784] = inform_R[776][4];				r_cell_reg[785] = inform_R[792][4];				r_cell_reg[786] = inform_R[777][4];				r_cell_reg[787] = inform_R[793][4];				r_cell_reg[788] = inform_R[778][4];				r_cell_reg[789] = inform_R[794][4];				r_cell_reg[790] = inform_R[779][4];				r_cell_reg[791] = inform_R[795][4];				r_cell_reg[792] = inform_R[780][4];				r_cell_reg[793] = inform_R[796][4];				r_cell_reg[794] = inform_R[781][4];				r_cell_reg[795] = inform_R[797][4];				r_cell_reg[796] = inform_R[782][4];				r_cell_reg[797] = inform_R[798][4];				r_cell_reg[798] = inform_R[783][4];				r_cell_reg[799] = inform_R[799][4];				r_cell_reg[800] = inform_R[800][4];				r_cell_reg[801] = inform_R[816][4];				r_cell_reg[802] = inform_R[801][4];				r_cell_reg[803] = inform_R[817][4];				r_cell_reg[804] = inform_R[802][4];				r_cell_reg[805] = inform_R[818][4];				r_cell_reg[806] = inform_R[803][4];				r_cell_reg[807] = inform_R[819][4];				r_cell_reg[808] = inform_R[804][4];				r_cell_reg[809] = inform_R[820][4];				r_cell_reg[810] = inform_R[805][4];				r_cell_reg[811] = inform_R[821][4];				r_cell_reg[812] = inform_R[806][4];				r_cell_reg[813] = inform_R[822][4];				r_cell_reg[814] = inform_R[807][4];				r_cell_reg[815] = inform_R[823][4];				r_cell_reg[816] = inform_R[808][4];				r_cell_reg[817] = inform_R[824][4];				r_cell_reg[818] = inform_R[809][4];				r_cell_reg[819] = inform_R[825][4];				r_cell_reg[820] = inform_R[810][4];				r_cell_reg[821] = inform_R[826][4];				r_cell_reg[822] = inform_R[811][4];				r_cell_reg[823] = inform_R[827][4];				r_cell_reg[824] = inform_R[812][4];				r_cell_reg[825] = inform_R[828][4];				r_cell_reg[826] = inform_R[813][4];				r_cell_reg[827] = inform_R[829][4];				r_cell_reg[828] = inform_R[814][4];				r_cell_reg[829] = inform_R[830][4];				r_cell_reg[830] = inform_R[815][4];				r_cell_reg[831] = inform_R[831][4];				r_cell_reg[832] = inform_R[832][4];				r_cell_reg[833] = inform_R[848][4];				r_cell_reg[834] = inform_R[833][4];				r_cell_reg[835] = inform_R[849][4];				r_cell_reg[836] = inform_R[834][4];				r_cell_reg[837] = inform_R[850][4];				r_cell_reg[838] = inform_R[835][4];				r_cell_reg[839] = inform_R[851][4];				r_cell_reg[840] = inform_R[836][4];				r_cell_reg[841] = inform_R[852][4];				r_cell_reg[842] = inform_R[837][4];				r_cell_reg[843] = inform_R[853][4];				r_cell_reg[844] = inform_R[838][4];				r_cell_reg[845] = inform_R[854][4];				r_cell_reg[846] = inform_R[839][4];				r_cell_reg[847] = inform_R[855][4];				r_cell_reg[848] = inform_R[840][4];				r_cell_reg[849] = inform_R[856][4];				r_cell_reg[850] = inform_R[841][4];				r_cell_reg[851] = inform_R[857][4];				r_cell_reg[852] = inform_R[842][4];				r_cell_reg[853] = inform_R[858][4];				r_cell_reg[854] = inform_R[843][4];				r_cell_reg[855] = inform_R[859][4];				r_cell_reg[856] = inform_R[844][4];				r_cell_reg[857] = inform_R[860][4];				r_cell_reg[858] = inform_R[845][4];				r_cell_reg[859] = inform_R[861][4];				r_cell_reg[860] = inform_R[846][4];				r_cell_reg[861] = inform_R[862][4];				r_cell_reg[862] = inform_R[847][4];				r_cell_reg[863] = inform_R[863][4];				r_cell_reg[864] = inform_R[864][4];				r_cell_reg[865] = inform_R[880][4];				r_cell_reg[866] = inform_R[865][4];				r_cell_reg[867] = inform_R[881][4];				r_cell_reg[868] = inform_R[866][4];				r_cell_reg[869] = inform_R[882][4];				r_cell_reg[870] = inform_R[867][4];				r_cell_reg[871] = inform_R[883][4];				r_cell_reg[872] = inform_R[868][4];				r_cell_reg[873] = inform_R[884][4];				r_cell_reg[874] = inform_R[869][4];				r_cell_reg[875] = inform_R[885][4];				r_cell_reg[876] = inform_R[870][4];				r_cell_reg[877] = inform_R[886][4];				r_cell_reg[878] = inform_R[871][4];				r_cell_reg[879] = inform_R[887][4];				r_cell_reg[880] = inform_R[872][4];				r_cell_reg[881] = inform_R[888][4];				r_cell_reg[882] = inform_R[873][4];				r_cell_reg[883] = inform_R[889][4];				r_cell_reg[884] = inform_R[874][4];				r_cell_reg[885] = inform_R[890][4];				r_cell_reg[886] = inform_R[875][4];				r_cell_reg[887] = inform_R[891][4];				r_cell_reg[888] = inform_R[876][4];				r_cell_reg[889] = inform_R[892][4];				r_cell_reg[890] = inform_R[877][4];				r_cell_reg[891] = inform_R[893][4];				r_cell_reg[892] = inform_R[878][4];				r_cell_reg[893] = inform_R[894][4];				r_cell_reg[894] = inform_R[879][4];				r_cell_reg[895] = inform_R[895][4];				r_cell_reg[896] = inform_R[896][4];				r_cell_reg[897] = inform_R[912][4];				r_cell_reg[898] = inform_R[897][4];				r_cell_reg[899] = inform_R[913][4];				r_cell_reg[900] = inform_R[898][4];				r_cell_reg[901] = inform_R[914][4];				r_cell_reg[902] = inform_R[899][4];				r_cell_reg[903] = inform_R[915][4];				r_cell_reg[904] = inform_R[900][4];				r_cell_reg[905] = inform_R[916][4];				r_cell_reg[906] = inform_R[901][4];				r_cell_reg[907] = inform_R[917][4];				r_cell_reg[908] = inform_R[902][4];				r_cell_reg[909] = inform_R[918][4];				r_cell_reg[910] = inform_R[903][4];				r_cell_reg[911] = inform_R[919][4];				r_cell_reg[912] = inform_R[904][4];				r_cell_reg[913] = inform_R[920][4];				r_cell_reg[914] = inform_R[905][4];				r_cell_reg[915] = inform_R[921][4];				r_cell_reg[916] = inform_R[906][4];				r_cell_reg[917] = inform_R[922][4];				r_cell_reg[918] = inform_R[907][4];				r_cell_reg[919] = inform_R[923][4];				r_cell_reg[920] = inform_R[908][4];				r_cell_reg[921] = inform_R[924][4];				r_cell_reg[922] = inform_R[909][4];				r_cell_reg[923] = inform_R[925][4];				r_cell_reg[924] = inform_R[910][4];				r_cell_reg[925] = inform_R[926][4];				r_cell_reg[926] = inform_R[911][4];				r_cell_reg[927] = inform_R[927][4];				r_cell_reg[928] = inform_R[928][4];				r_cell_reg[929] = inform_R[944][4];				r_cell_reg[930] = inform_R[929][4];				r_cell_reg[931] = inform_R[945][4];				r_cell_reg[932] = inform_R[930][4];				r_cell_reg[933] = inform_R[946][4];				r_cell_reg[934] = inform_R[931][4];				r_cell_reg[935] = inform_R[947][4];				r_cell_reg[936] = inform_R[932][4];				r_cell_reg[937] = inform_R[948][4];				r_cell_reg[938] = inform_R[933][4];				r_cell_reg[939] = inform_R[949][4];				r_cell_reg[940] = inform_R[934][4];				r_cell_reg[941] = inform_R[950][4];				r_cell_reg[942] = inform_R[935][4];				r_cell_reg[943] = inform_R[951][4];				r_cell_reg[944] = inform_R[936][4];				r_cell_reg[945] = inform_R[952][4];				r_cell_reg[946] = inform_R[937][4];				r_cell_reg[947] = inform_R[953][4];				r_cell_reg[948] = inform_R[938][4];				r_cell_reg[949] = inform_R[954][4];				r_cell_reg[950] = inform_R[939][4];				r_cell_reg[951] = inform_R[955][4];				r_cell_reg[952] = inform_R[940][4];				r_cell_reg[953] = inform_R[956][4];				r_cell_reg[954] = inform_R[941][4];				r_cell_reg[955] = inform_R[957][4];				r_cell_reg[956] = inform_R[942][4];				r_cell_reg[957] = inform_R[958][4];				r_cell_reg[958] = inform_R[943][4];				r_cell_reg[959] = inform_R[959][4];				r_cell_reg[960] = inform_R[960][4];				r_cell_reg[961] = inform_R[976][4];				r_cell_reg[962] = inform_R[961][4];				r_cell_reg[963] = inform_R[977][4];				r_cell_reg[964] = inform_R[962][4];				r_cell_reg[965] = inform_R[978][4];				r_cell_reg[966] = inform_R[963][4];				r_cell_reg[967] = inform_R[979][4];				r_cell_reg[968] = inform_R[964][4];				r_cell_reg[969] = inform_R[980][4];				r_cell_reg[970] = inform_R[965][4];				r_cell_reg[971] = inform_R[981][4];				r_cell_reg[972] = inform_R[966][4];				r_cell_reg[973] = inform_R[982][4];				r_cell_reg[974] = inform_R[967][4];				r_cell_reg[975] = inform_R[983][4];				r_cell_reg[976] = inform_R[968][4];				r_cell_reg[977] = inform_R[984][4];				r_cell_reg[978] = inform_R[969][4];				r_cell_reg[979] = inform_R[985][4];				r_cell_reg[980] = inform_R[970][4];				r_cell_reg[981] = inform_R[986][4];				r_cell_reg[982] = inform_R[971][4];				r_cell_reg[983] = inform_R[987][4];				r_cell_reg[984] = inform_R[972][4];				r_cell_reg[985] = inform_R[988][4];				r_cell_reg[986] = inform_R[973][4];				r_cell_reg[987] = inform_R[989][4];				r_cell_reg[988] = inform_R[974][4];				r_cell_reg[989] = inform_R[990][4];				r_cell_reg[990] = inform_R[975][4];				r_cell_reg[991] = inform_R[991][4];				r_cell_reg[992] = inform_R[992][4];				r_cell_reg[993] = inform_R[1008][4];				r_cell_reg[994] = inform_R[993][4];				r_cell_reg[995] = inform_R[1009][4];				r_cell_reg[996] = inform_R[994][4];				r_cell_reg[997] = inform_R[1010][4];				r_cell_reg[998] = inform_R[995][4];				r_cell_reg[999] = inform_R[1011][4];				r_cell_reg[1000] = inform_R[996][4];				r_cell_reg[1001] = inform_R[1012][4];				r_cell_reg[1002] = inform_R[997][4];				r_cell_reg[1003] = inform_R[1013][4];				r_cell_reg[1004] = inform_R[998][4];				r_cell_reg[1005] = inform_R[1014][4];				r_cell_reg[1006] = inform_R[999][4];				r_cell_reg[1007] = inform_R[1015][4];				r_cell_reg[1008] = inform_R[1000][4];				r_cell_reg[1009] = inform_R[1016][4];				r_cell_reg[1010] = inform_R[1001][4];				r_cell_reg[1011] = inform_R[1017][4];				r_cell_reg[1012] = inform_R[1002][4];				r_cell_reg[1013] = inform_R[1018][4];				r_cell_reg[1014] = inform_R[1003][4];				r_cell_reg[1015] = inform_R[1019][4];				r_cell_reg[1016] = inform_R[1004][4];				r_cell_reg[1017] = inform_R[1020][4];				r_cell_reg[1018] = inform_R[1005][4];				r_cell_reg[1019] = inform_R[1021][4];				r_cell_reg[1020] = inform_R[1006][4];				r_cell_reg[1021] = inform_R[1022][4];				r_cell_reg[1022] = inform_R[1007][4];				r_cell_reg[1023] = inform_R[1023][4];				l_cell_reg[0] = inform_L[0][5];				l_cell_reg[1] = inform_L[16][5];				l_cell_reg[2] = inform_L[1][5];				l_cell_reg[3] = inform_L[17][5];				l_cell_reg[4] = inform_L[2][5];				l_cell_reg[5] = inform_L[18][5];				l_cell_reg[6] = inform_L[3][5];				l_cell_reg[7] = inform_L[19][5];				l_cell_reg[8] = inform_L[4][5];				l_cell_reg[9] = inform_L[20][5];				l_cell_reg[10] = inform_L[5][5];				l_cell_reg[11] = inform_L[21][5];				l_cell_reg[12] = inform_L[6][5];				l_cell_reg[13] = inform_L[22][5];				l_cell_reg[14] = inform_L[7][5];				l_cell_reg[15] = inform_L[23][5];				l_cell_reg[16] = inform_L[8][5];				l_cell_reg[17] = inform_L[24][5];				l_cell_reg[18] = inform_L[9][5];				l_cell_reg[19] = inform_L[25][5];				l_cell_reg[20] = inform_L[10][5];				l_cell_reg[21] = inform_L[26][5];				l_cell_reg[22] = inform_L[11][5];				l_cell_reg[23] = inform_L[27][5];				l_cell_reg[24] = inform_L[12][5];				l_cell_reg[25] = inform_L[28][5];				l_cell_reg[26] = inform_L[13][5];				l_cell_reg[27] = inform_L[29][5];				l_cell_reg[28] = inform_L[14][5];				l_cell_reg[29] = inform_L[30][5];				l_cell_reg[30] = inform_L[15][5];				l_cell_reg[31] = inform_L[31][5];				l_cell_reg[32] = inform_L[32][5];				l_cell_reg[33] = inform_L[48][5];				l_cell_reg[34] = inform_L[33][5];				l_cell_reg[35] = inform_L[49][5];				l_cell_reg[36] = inform_L[34][5];				l_cell_reg[37] = inform_L[50][5];				l_cell_reg[38] = inform_L[35][5];				l_cell_reg[39] = inform_L[51][5];				l_cell_reg[40] = inform_L[36][5];				l_cell_reg[41] = inform_L[52][5];				l_cell_reg[42] = inform_L[37][5];				l_cell_reg[43] = inform_L[53][5];				l_cell_reg[44] = inform_L[38][5];				l_cell_reg[45] = inform_L[54][5];				l_cell_reg[46] = inform_L[39][5];				l_cell_reg[47] = inform_L[55][5];				l_cell_reg[48] = inform_L[40][5];				l_cell_reg[49] = inform_L[56][5];				l_cell_reg[50] = inform_L[41][5];				l_cell_reg[51] = inform_L[57][5];				l_cell_reg[52] = inform_L[42][5];				l_cell_reg[53] = inform_L[58][5];				l_cell_reg[54] = inform_L[43][5];				l_cell_reg[55] = inform_L[59][5];				l_cell_reg[56] = inform_L[44][5];				l_cell_reg[57] = inform_L[60][5];				l_cell_reg[58] = inform_L[45][5];				l_cell_reg[59] = inform_L[61][5];				l_cell_reg[60] = inform_L[46][5];				l_cell_reg[61] = inform_L[62][5];				l_cell_reg[62] = inform_L[47][5];				l_cell_reg[63] = inform_L[63][5];				l_cell_reg[64] = inform_L[64][5];				l_cell_reg[65] = inform_L[80][5];				l_cell_reg[66] = inform_L[65][5];				l_cell_reg[67] = inform_L[81][5];				l_cell_reg[68] = inform_L[66][5];				l_cell_reg[69] = inform_L[82][5];				l_cell_reg[70] = inform_L[67][5];				l_cell_reg[71] = inform_L[83][5];				l_cell_reg[72] = inform_L[68][5];				l_cell_reg[73] = inform_L[84][5];				l_cell_reg[74] = inform_L[69][5];				l_cell_reg[75] = inform_L[85][5];				l_cell_reg[76] = inform_L[70][5];				l_cell_reg[77] = inform_L[86][5];				l_cell_reg[78] = inform_L[71][5];				l_cell_reg[79] = inform_L[87][5];				l_cell_reg[80] = inform_L[72][5];				l_cell_reg[81] = inform_L[88][5];				l_cell_reg[82] = inform_L[73][5];				l_cell_reg[83] = inform_L[89][5];				l_cell_reg[84] = inform_L[74][5];				l_cell_reg[85] = inform_L[90][5];				l_cell_reg[86] = inform_L[75][5];				l_cell_reg[87] = inform_L[91][5];				l_cell_reg[88] = inform_L[76][5];				l_cell_reg[89] = inform_L[92][5];				l_cell_reg[90] = inform_L[77][5];				l_cell_reg[91] = inform_L[93][5];				l_cell_reg[92] = inform_L[78][5];				l_cell_reg[93] = inform_L[94][5];				l_cell_reg[94] = inform_L[79][5];				l_cell_reg[95] = inform_L[95][5];				l_cell_reg[96] = inform_L[96][5];				l_cell_reg[97] = inform_L[112][5];				l_cell_reg[98] = inform_L[97][5];				l_cell_reg[99] = inform_L[113][5];				l_cell_reg[100] = inform_L[98][5];				l_cell_reg[101] = inform_L[114][5];				l_cell_reg[102] = inform_L[99][5];				l_cell_reg[103] = inform_L[115][5];				l_cell_reg[104] = inform_L[100][5];				l_cell_reg[105] = inform_L[116][5];				l_cell_reg[106] = inform_L[101][5];				l_cell_reg[107] = inform_L[117][5];				l_cell_reg[108] = inform_L[102][5];				l_cell_reg[109] = inform_L[118][5];				l_cell_reg[110] = inform_L[103][5];				l_cell_reg[111] = inform_L[119][5];				l_cell_reg[112] = inform_L[104][5];				l_cell_reg[113] = inform_L[120][5];				l_cell_reg[114] = inform_L[105][5];				l_cell_reg[115] = inform_L[121][5];				l_cell_reg[116] = inform_L[106][5];				l_cell_reg[117] = inform_L[122][5];				l_cell_reg[118] = inform_L[107][5];				l_cell_reg[119] = inform_L[123][5];				l_cell_reg[120] = inform_L[108][5];				l_cell_reg[121] = inform_L[124][5];				l_cell_reg[122] = inform_L[109][5];				l_cell_reg[123] = inform_L[125][5];				l_cell_reg[124] = inform_L[110][5];				l_cell_reg[125] = inform_L[126][5];				l_cell_reg[126] = inform_L[111][5];				l_cell_reg[127] = inform_L[127][5];				l_cell_reg[128] = inform_L[128][5];				l_cell_reg[129] = inform_L[144][5];				l_cell_reg[130] = inform_L[129][5];				l_cell_reg[131] = inform_L[145][5];				l_cell_reg[132] = inform_L[130][5];				l_cell_reg[133] = inform_L[146][5];				l_cell_reg[134] = inform_L[131][5];				l_cell_reg[135] = inform_L[147][5];				l_cell_reg[136] = inform_L[132][5];				l_cell_reg[137] = inform_L[148][5];				l_cell_reg[138] = inform_L[133][5];				l_cell_reg[139] = inform_L[149][5];				l_cell_reg[140] = inform_L[134][5];				l_cell_reg[141] = inform_L[150][5];				l_cell_reg[142] = inform_L[135][5];				l_cell_reg[143] = inform_L[151][5];				l_cell_reg[144] = inform_L[136][5];				l_cell_reg[145] = inform_L[152][5];				l_cell_reg[146] = inform_L[137][5];				l_cell_reg[147] = inform_L[153][5];				l_cell_reg[148] = inform_L[138][5];				l_cell_reg[149] = inform_L[154][5];				l_cell_reg[150] = inform_L[139][5];				l_cell_reg[151] = inform_L[155][5];				l_cell_reg[152] = inform_L[140][5];				l_cell_reg[153] = inform_L[156][5];				l_cell_reg[154] = inform_L[141][5];				l_cell_reg[155] = inform_L[157][5];				l_cell_reg[156] = inform_L[142][5];				l_cell_reg[157] = inform_L[158][5];				l_cell_reg[158] = inform_L[143][5];				l_cell_reg[159] = inform_L[159][5];				l_cell_reg[160] = inform_L[160][5];				l_cell_reg[161] = inform_L[176][5];				l_cell_reg[162] = inform_L[161][5];				l_cell_reg[163] = inform_L[177][5];				l_cell_reg[164] = inform_L[162][5];				l_cell_reg[165] = inform_L[178][5];				l_cell_reg[166] = inform_L[163][5];				l_cell_reg[167] = inform_L[179][5];				l_cell_reg[168] = inform_L[164][5];				l_cell_reg[169] = inform_L[180][5];				l_cell_reg[170] = inform_L[165][5];				l_cell_reg[171] = inform_L[181][5];				l_cell_reg[172] = inform_L[166][5];				l_cell_reg[173] = inform_L[182][5];				l_cell_reg[174] = inform_L[167][5];				l_cell_reg[175] = inform_L[183][5];				l_cell_reg[176] = inform_L[168][5];				l_cell_reg[177] = inform_L[184][5];				l_cell_reg[178] = inform_L[169][5];				l_cell_reg[179] = inform_L[185][5];				l_cell_reg[180] = inform_L[170][5];				l_cell_reg[181] = inform_L[186][5];				l_cell_reg[182] = inform_L[171][5];				l_cell_reg[183] = inform_L[187][5];				l_cell_reg[184] = inform_L[172][5];				l_cell_reg[185] = inform_L[188][5];				l_cell_reg[186] = inform_L[173][5];				l_cell_reg[187] = inform_L[189][5];				l_cell_reg[188] = inform_L[174][5];				l_cell_reg[189] = inform_L[190][5];				l_cell_reg[190] = inform_L[175][5];				l_cell_reg[191] = inform_L[191][5];				l_cell_reg[192] = inform_L[192][5];				l_cell_reg[193] = inform_L[208][5];				l_cell_reg[194] = inform_L[193][5];				l_cell_reg[195] = inform_L[209][5];				l_cell_reg[196] = inform_L[194][5];				l_cell_reg[197] = inform_L[210][5];				l_cell_reg[198] = inform_L[195][5];				l_cell_reg[199] = inform_L[211][5];				l_cell_reg[200] = inform_L[196][5];				l_cell_reg[201] = inform_L[212][5];				l_cell_reg[202] = inform_L[197][5];				l_cell_reg[203] = inform_L[213][5];				l_cell_reg[204] = inform_L[198][5];				l_cell_reg[205] = inform_L[214][5];				l_cell_reg[206] = inform_L[199][5];				l_cell_reg[207] = inform_L[215][5];				l_cell_reg[208] = inform_L[200][5];				l_cell_reg[209] = inform_L[216][5];				l_cell_reg[210] = inform_L[201][5];				l_cell_reg[211] = inform_L[217][5];				l_cell_reg[212] = inform_L[202][5];				l_cell_reg[213] = inform_L[218][5];				l_cell_reg[214] = inform_L[203][5];				l_cell_reg[215] = inform_L[219][5];				l_cell_reg[216] = inform_L[204][5];				l_cell_reg[217] = inform_L[220][5];				l_cell_reg[218] = inform_L[205][5];				l_cell_reg[219] = inform_L[221][5];				l_cell_reg[220] = inform_L[206][5];				l_cell_reg[221] = inform_L[222][5];				l_cell_reg[222] = inform_L[207][5];				l_cell_reg[223] = inform_L[223][5];				l_cell_reg[224] = inform_L[224][5];				l_cell_reg[225] = inform_L[240][5];				l_cell_reg[226] = inform_L[225][5];				l_cell_reg[227] = inform_L[241][5];				l_cell_reg[228] = inform_L[226][5];				l_cell_reg[229] = inform_L[242][5];				l_cell_reg[230] = inform_L[227][5];				l_cell_reg[231] = inform_L[243][5];				l_cell_reg[232] = inform_L[228][5];				l_cell_reg[233] = inform_L[244][5];				l_cell_reg[234] = inform_L[229][5];				l_cell_reg[235] = inform_L[245][5];				l_cell_reg[236] = inform_L[230][5];				l_cell_reg[237] = inform_L[246][5];				l_cell_reg[238] = inform_L[231][5];				l_cell_reg[239] = inform_L[247][5];				l_cell_reg[240] = inform_L[232][5];				l_cell_reg[241] = inform_L[248][5];				l_cell_reg[242] = inform_L[233][5];				l_cell_reg[243] = inform_L[249][5];				l_cell_reg[244] = inform_L[234][5];				l_cell_reg[245] = inform_L[250][5];				l_cell_reg[246] = inform_L[235][5];				l_cell_reg[247] = inform_L[251][5];				l_cell_reg[248] = inform_L[236][5];				l_cell_reg[249] = inform_L[252][5];				l_cell_reg[250] = inform_L[237][5];				l_cell_reg[251] = inform_L[253][5];				l_cell_reg[252] = inform_L[238][5];				l_cell_reg[253] = inform_L[254][5];				l_cell_reg[254] = inform_L[239][5];				l_cell_reg[255] = inform_L[255][5];				l_cell_reg[256] = inform_L[256][5];				l_cell_reg[257] = inform_L[272][5];				l_cell_reg[258] = inform_L[257][5];				l_cell_reg[259] = inform_L[273][5];				l_cell_reg[260] = inform_L[258][5];				l_cell_reg[261] = inform_L[274][5];				l_cell_reg[262] = inform_L[259][5];				l_cell_reg[263] = inform_L[275][5];				l_cell_reg[264] = inform_L[260][5];				l_cell_reg[265] = inform_L[276][5];				l_cell_reg[266] = inform_L[261][5];				l_cell_reg[267] = inform_L[277][5];				l_cell_reg[268] = inform_L[262][5];				l_cell_reg[269] = inform_L[278][5];				l_cell_reg[270] = inform_L[263][5];				l_cell_reg[271] = inform_L[279][5];				l_cell_reg[272] = inform_L[264][5];				l_cell_reg[273] = inform_L[280][5];				l_cell_reg[274] = inform_L[265][5];				l_cell_reg[275] = inform_L[281][5];				l_cell_reg[276] = inform_L[266][5];				l_cell_reg[277] = inform_L[282][5];				l_cell_reg[278] = inform_L[267][5];				l_cell_reg[279] = inform_L[283][5];				l_cell_reg[280] = inform_L[268][5];				l_cell_reg[281] = inform_L[284][5];				l_cell_reg[282] = inform_L[269][5];				l_cell_reg[283] = inform_L[285][5];				l_cell_reg[284] = inform_L[270][5];				l_cell_reg[285] = inform_L[286][5];				l_cell_reg[286] = inform_L[271][5];				l_cell_reg[287] = inform_L[287][5];				l_cell_reg[288] = inform_L[288][5];				l_cell_reg[289] = inform_L[304][5];				l_cell_reg[290] = inform_L[289][5];				l_cell_reg[291] = inform_L[305][5];				l_cell_reg[292] = inform_L[290][5];				l_cell_reg[293] = inform_L[306][5];				l_cell_reg[294] = inform_L[291][5];				l_cell_reg[295] = inform_L[307][5];				l_cell_reg[296] = inform_L[292][5];				l_cell_reg[297] = inform_L[308][5];				l_cell_reg[298] = inform_L[293][5];				l_cell_reg[299] = inform_L[309][5];				l_cell_reg[300] = inform_L[294][5];				l_cell_reg[301] = inform_L[310][5];				l_cell_reg[302] = inform_L[295][5];				l_cell_reg[303] = inform_L[311][5];				l_cell_reg[304] = inform_L[296][5];				l_cell_reg[305] = inform_L[312][5];				l_cell_reg[306] = inform_L[297][5];				l_cell_reg[307] = inform_L[313][5];				l_cell_reg[308] = inform_L[298][5];				l_cell_reg[309] = inform_L[314][5];				l_cell_reg[310] = inform_L[299][5];				l_cell_reg[311] = inform_L[315][5];				l_cell_reg[312] = inform_L[300][5];				l_cell_reg[313] = inform_L[316][5];				l_cell_reg[314] = inform_L[301][5];				l_cell_reg[315] = inform_L[317][5];				l_cell_reg[316] = inform_L[302][5];				l_cell_reg[317] = inform_L[318][5];				l_cell_reg[318] = inform_L[303][5];				l_cell_reg[319] = inform_L[319][5];				l_cell_reg[320] = inform_L[320][5];				l_cell_reg[321] = inform_L[336][5];				l_cell_reg[322] = inform_L[321][5];				l_cell_reg[323] = inform_L[337][5];				l_cell_reg[324] = inform_L[322][5];				l_cell_reg[325] = inform_L[338][5];				l_cell_reg[326] = inform_L[323][5];				l_cell_reg[327] = inform_L[339][5];				l_cell_reg[328] = inform_L[324][5];				l_cell_reg[329] = inform_L[340][5];				l_cell_reg[330] = inform_L[325][5];				l_cell_reg[331] = inform_L[341][5];				l_cell_reg[332] = inform_L[326][5];				l_cell_reg[333] = inform_L[342][5];				l_cell_reg[334] = inform_L[327][5];				l_cell_reg[335] = inform_L[343][5];				l_cell_reg[336] = inform_L[328][5];				l_cell_reg[337] = inform_L[344][5];				l_cell_reg[338] = inform_L[329][5];				l_cell_reg[339] = inform_L[345][5];				l_cell_reg[340] = inform_L[330][5];				l_cell_reg[341] = inform_L[346][5];				l_cell_reg[342] = inform_L[331][5];				l_cell_reg[343] = inform_L[347][5];				l_cell_reg[344] = inform_L[332][5];				l_cell_reg[345] = inform_L[348][5];				l_cell_reg[346] = inform_L[333][5];				l_cell_reg[347] = inform_L[349][5];				l_cell_reg[348] = inform_L[334][5];				l_cell_reg[349] = inform_L[350][5];				l_cell_reg[350] = inform_L[335][5];				l_cell_reg[351] = inform_L[351][5];				l_cell_reg[352] = inform_L[352][5];				l_cell_reg[353] = inform_L[368][5];				l_cell_reg[354] = inform_L[353][5];				l_cell_reg[355] = inform_L[369][5];				l_cell_reg[356] = inform_L[354][5];				l_cell_reg[357] = inform_L[370][5];				l_cell_reg[358] = inform_L[355][5];				l_cell_reg[359] = inform_L[371][5];				l_cell_reg[360] = inform_L[356][5];				l_cell_reg[361] = inform_L[372][5];				l_cell_reg[362] = inform_L[357][5];				l_cell_reg[363] = inform_L[373][5];				l_cell_reg[364] = inform_L[358][5];				l_cell_reg[365] = inform_L[374][5];				l_cell_reg[366] = inform_L[359][5];				l_cell_reg[367] = inform_L[375][5];				l_cell_reg[368] = inform_L[360][5];				l_cell_reg[369] = inform_L[376][5];				l_cell_reg[370] = inform_L[361][5];				l_cell_reg[371] = inform_L[377][5];				l_cell_reg[372] = inform_L[362][5];				l_cell_reg[373] = inform_L[378][5];				l_cell_reg[374] = inform_L[363][5];				l_cell_reg[375] = inform_L[379][5];				l_cell_reg[376] = inform_L[364][5];				l_cell_reg[377] = inform_L[380][5];				l_cell_reg[378] = inform_L[365][5];				l_cell_reg[379] = inform_L[381][5];				l_cell_reg[380] = inform_L[366][5];				l_cell_reg[381] = inform_L[382][5];				l_cell_reg[382] = inform_L[367][5];				l_cell_reg[383] = inform_L[383][5];				l_cell_reg[384] = inform_L[384][5];				l_cell_reg[385] = inform_L[400][5];				l_cell_reg[386] = inform_L[385][5];				l_cell_reg[387] = inform_L[401][5];				l_cell_reg[388] = inform_L[386][5];				l_cell_reg[389] = inform_L[402][5];				l_cell_reg[390] = inform_L[387][5];				l_cell_reg[391] = inform_L[403][5];				l_cell_reg[392] = inform_L[388][5];				l_cell_reg[393] = inform_L[404][5];				l_cell_reg[394] = inform_L[389][5];				l_cell_reg[395] = inform_L[405][5];				l_cell_reg[396] = inform_L[390][5];				l_cell_reg[397] = inform_L[406][5];				l_cell_reg[398] = inform_L[391][5];				l_cell_reg[399] = inform_L[407][5];				l_cell_reg[400] = inform_L[392][5];				l_cell_reg[401] = inform_L[408][5];				l_cell_reg[402] = inform_L[393][5];				l_cell_reg[403] = inform_L[409][5];				l_cell_reg[404] = inform_L[394][5];				l_cell_reg[405] = inform_L[410][5];				l_cell_reg[406] = inform_L[395][5];				l_cell_reg[407] = inform_L[411][5];				l_cell_reg[408] = inform_L[396][5];				l_cell_reg[409] = inform_L[412][5];				l_cell_reg[410] = inform_L[397][5];				l_cell_reg[411] = inform_L[413][5];				l_cell_reg[412] = inform_L[398][5];				l_cell_reg[413] = inform_L[414][5];				l_cell_reg[414] = inform_L[399][5];				l_cell_reg[415] = inform_L[415][5];				l_cell_reg[416] = inform_L[416][5];				l_cell_reg[417] = inform_L[432][5];				l_cell_reg[418] = inform_L[417][5];				l_cell_reg[419] = inform_L[433][5];				l_cell_reg[420] = inform_L[418][5];				l_cell_reg[421] = inform_L[434][5];				l_cell_reg[422] = inform_L[419][5];				l_cell_reg[423] = inform_L[435][5];				l_cell_reg[424] = inform_L[420][5];				l_cell_reg[425] = inform_L[436][5];				l_cell_reg[426] = inform_L[421][5];				l_cell_reg[427] = inform_L[437][5];				l_cell_reg[428] = inform_L[422][5];				l_cell_reg[429] = inform_L[438][5];				l_cell_reg[430] = inform_L[423][5];				l_cell_reg[431] = inform_L[439][5];				l_cell_reg[432] = inform_L[424][5];				l_cell_reg[433] = inform_L[440][5];				l_cell_reg[434] = inform_L[425][5];				l_cell_reg[435] = inform_L[441][5];				l_cell_reg[436] = inform_L[426][5];				l_cell_reg[437] = inform_L[442][5];				l_cell_reg[438] = inform_L[427][5];				l_cell_reg[439] = inform_L[443][5];				l_cell_reg[440] = inform_L[428][5];				l_cell_reg[441] = inform_L[444][5];				l_cell_reg[442] = inform_L[429][5];				l_cell_reg[443] = inform_L[445][5];				l_cell_reg[444] = inform_L[430][5];				l_cell_reg[445] = inform_L[446][5];				l_cell_reg[446] = inform_L[431][5];				l_cell_reg[447] = inform_L[447][5];				l_cell_reg[448] = inform_L[448][5];				l_cell_reg[449] = inform_L[464][5];				l_cell_reg[450] = inform_L[449][5];				l_cell_reg[451] = inform_L[465][5];				l_cell_reg[452] = inform_L[450][5];				l_cell_reg[453] = inform_L[466][5];				l_cell_reg[454] = inform_L[451][5];				l_cell_reg[455] = inform_L[467][5];				l_cell_reg[456] = inform_L[452][5];				l_cell_reg[457] = inform_L[468][5];				l_cell_reg[458] = inform_L[453][5];				l_cell_reg[459] = inform_L[469][5];				l_cell_reg[460] = inform_L[454][5];				l_cell_reg[461] = inform_L[470][5];				l_cell_reg[462] = inform_L[455][5];				l_cell_reg[463] = inform_L[471][5];				l_cell_reg[464] = inform_L[456][5];				l_cell_reg[465] = inform_L[472][5];				l_cell_reg[466] = inform_L[457][5];				l_cell_reg[467] = inform_L[473][5];				l_cell_reg[468] = inform_L[458][5];				l_cell_reg[469] = inform_L[474][5];				l_cell_reg[470] = inform_L[459][5];				l_cell_reg[471] = inform_L[475][5];				l_cell_reg[472] = inform_L[460][5];				l_cell_reg[473] = inform_L[476][5];				l_cell_reg[474] = inform_L[461][5];				l_cell_reg[475] = inform_L[477][5];				l_cell_reg[476] = inform_L[462][5];				l_cell_reg[477] = inform_L[478][5];				l_cell_reg[478] = inform_L[463][5];				l_cell_reg[479] = inform_L[479][5];				l_cell_reg[480] = inform_L[480][5];				l_cell_reg[481] = inform_L[496][5];				l_cell_reg[482] = inform_L[481][5];				l_cell_reg[483] = inform_L[497][5];				l_cell_reg[484] = inform_L[482][5];				l_cell_reg[485] = inform_L[498][5];				l_cell_reg[486] = inform_L[483][5];				l_cell_reg[487] = inform_L[499][5];				l_cell_reg[488] = inform_L[484][5];				l_cell_reg[489] = inform_L[500][5];				l_cell_reg[490] = inform_L[485][5];				l_cell_reg[491] = inform_L[501][5];				l_cell_reg[492] = inform_L[486][5];				l_cell_reg[493] = inform_L[502][5];				l_cell_reg[494] = inform_L[487][5];				l_cell_reg[495] = inform_L[503][5];				l_cell_reg[496] = inform_L[488][5];				l_cell_reg[497] = inform_L[504][5];				l_cell_reg[498] = inform_L[489][5];				l_cell_reg[499] = inform_L[505][5];				l_cell_reg[500] = inform_L[490][5];				l_cell_reg[501] = inform_L[506][5];				l_cell_reg[502] = inform_L[491][5];				l_cell_reg[503] = inform_L[507][5];				l_cell_reg[504] = inform_L[492][5];				l_cell_reg[505] = inform_L[508][5];				l_cell_reg[506] = inform_L[493][5];				l_cell_reg[507] = inform_L[509][5];				l_cell_reg[508] = inform_L[494][5];				l_cell_reg[509] = inform_L[510][5];				l_cell_reg[510] = inform_L[495][5];				l_cell_reg[511] = inform_L[511][5];				l_cell_reg[512] = inform_L[512][5];				l_cell_reg[513] = inform_L[528][5];				l_cell_reg[514] = inform_L[513][5];				l_cell_reg[515] = inform_L[529][5];				l_cell_reg[516] = inform_L[514][5];				l_cell_reg[517] = inform_L[530][5];				l_cell_reg[518] = inform_L[515][5];				l_cell_reg[519] = inform_L[531][5];				l_cell_reg[520] = inform_L[516][5];				l_cell_reg[521] = inform_L[532][5];				l_cell_reg[522] = inform_L[517][5];				l_cell_reg[523] = inform_L[533][5];				l_cell_reg[524] = inform_L[518][5];				l_cell_reg[525] = inform_L[534][5];				l_cell_reg[526] = inform_L[519][5];				l_cell_reg[527] = inform_L[535][5];				l_cell_reg[528] = inform_L[520][5];				l_cell_reg[529] = inform_L[536][5];				l_cell_reg[530] = inform_L[521][5];				l_cell_reg[531] = inform_L[537][5];				l_cell_reg[532] = inform_L[522][5];				l_cell_reg[533] = inform_L[538][5];				l_cell_reg[534] = inform_L[523][5];				l_cell_reg[535] = inform_L[539][5];				l_cell_reg[536] = inform_L[524][5];				l_cell_reg[537] = inform_L[540][5];				l_cell_reg[538] = inform_L[525][5];				l_cell_reg[539] = inform_L[541][5];				l_cell_reg[540] = inform_L[526][5];				l_cell_reg[541] = inform_L[542][5];				l_cell_reg[542] = inform_L[527][5];				l_cell_reg[543] = inform_L[543][5];				l_cell_reg[544] = inform_L[544][5];				l_cell_reg[545] = inform_L[560][5];				l_cell_reg[546] = inform_L[545][5];				l_cell_reg[547] = inform_L[561][5];				l_cell_reg[548] = inform_L[546][5];				l_cell_reg[549] = inform_L[562][5];				l_cell_reg[550] = inform_L[547][5];				l_cell_reg[551] = inform_L[563][5];				l_cell_reg[552] = inform_L[548][5];				l_cell_reg[553] = inform_L[564][5];				l_cell_reg[554] = inform_L[549][5];				l_cell_reg[555] = inform_L[565][5];				l_cell_reg[556] = inform_L[550][5];				l_cell_reg[557] = inform_L[566][5];				l_cell_reg[558] = inform_L[551][5];				l_cell_reg[559] = inform_L[567][5];				l_cell_reg[560] = inform_L[552][5];				l_cell_reg[561] = inform_L[568][5];				l_cell_reg[562] = inform_L[553][5];				l_cell_reg[563] = inform_L[569][5];				l_cell_reg[564] = inform_L[554][5];				l_cell_reg[565] = inform_L[570][5];				l_cell_reg[566] = inform_L[555][5];				l_cell_reg[567] = inform_L[571][5];				l_cell_reg[568] = inform_L[556][5];				l_cell_reg[569] = inform_L[572][5];				l_cell_reg[570] = inform_L[557][5];				l_cell_reg[571] = inform_L[573][5];				l_cell_reg[572] = inform_L[558][5];				l_cell_reg[573] = inform_L[574][5];				l_cell_reg[574] = inform_L[559][5];				l_cell_reg[575] = inform_L[575][5];				l_cell_reg[576] = inform_L[576][5];				l_cell_reg[577] = inform_L[592][5];				l_cell_reg[578] = inform_L[577][5];				l_cell_reg[579] = inform_L[593][5];				l_cell_reg[580] = inform_L[578][5];				l_cell_reg[581] = inform_L[594][5];				l_cell_reg[582] = inform_L[579][5];				l_cell_reg[583] = inform_L[595][5];				l_cell_reg[584] = inform_L[580][5];				l_cell_reg[585] = inform_L[596][5];				l_cell_reg[586] = inform_L[581][5];				l_cell_reg[587] = inform_L[597][5];				l_cell_reg[588] = inform_L[582][5];				l_cell_reg[589] = inform_L[598][5];				l_cell_reg[590] = inform_L[583][5];				l_cell_reg[591] = inform_L[599][5];				l_cell_reg[592] = inform_L[584][5];				l_cell_reg[593] = inform_L[600][5];				l_cell_reg[594] = inform_L[585][5];				l_cell_reg[595] = inform_L[601][5];				l_cell_reg[596] = inform_L[586][5];				l_cell_reg[597] = inform_L[602][5];				l_cell_reg[598] = inform_L[587][5];				l_cell_reg[599] = inform_L[603][5];				l_cell_reg[600] = inform_L[588][5];				l_cell_reg[601] = inform_L[604][5];				l_cell_reg[602] = inform_L[589][5];				l_cell_reg[603] = inform_L[605][5];				l_cell_reg[604] = inform_L[590][5];				l_cell_reg[605] = inform_L[606][5];				l_cell_reg[606] = inform_L[591][5];				l_cell_reg[607] = inform_L[607][5];				l_cell_reg[608] = inform_L[608][5];				l_cell_reg[609] = inform_L[624][5];				l_cell_reg[610] = inform_L[609][5];				l_cell_reg[611] = inform_L[625][5];				l_cell_reg[612] = inform_L[610][5];				l_cell_reg[613] = inform_L[626][5];				l_cell_reg[614] = inform_L[611][5];				l_cell_reg[615] = inform_L[627][5];				l_cell_reg[616] = inform_L[612][5];				l_cell_reg[617] = inform_L[628][5];				l_cell_reg[618] = inform_L[613][5];				l_cell_reg[619] = inform_L[629][5];				l_cell_reg[620] = inform_L[614][5];				l_cell_reg[621] = inform_L[630][5];				l_cell_reg[622] = inform_L[615][5];				l_cell_reg[623] = inform_L[631][5];				l_cell_reg[624] = inform_L[616][5];				l_cell_reg[625] = inform_L[632][5];				l_cell_reg[626] = inform_L[617][5];				l_cell_reg[627] = inform_L[633][5];				l_cell_reg[628] = inform_L[618][5];				l_cell_reg[629] = inform_L[634][5];				l_cell_reg[630] = inform_L[619][5];				l_cell_reg[631] = inform_L[635][5];				l_cell_reg[632] = inform_L[620][5];				l_cell_reg[633] = inform_L[636][5];				l_cell_reg[634] = inform_L[621][5];				l_cell_reg[635] = inform_L[637][5];				l_cell_reg[636] = inform_L[622][5];				l_cell_reg[637] = inform_L[638][5];				l_cell_reg[638] = inform_L[623][5];				l_cell_reg[639] = inform_L[639][5];				l_cell_reg[640] = inform_L[640][5];				l_cell_reg[641] = inform_L[656][5];				l_cell_reg[642] = inform_L[641][5];				l_cell_reg[643] = inform_L[657][5];				l_cell_reg[644] = inform_L[642][5];				l_cell_reg[645] = inform_L[658][5];				l_cell_reg[646] = inform_L[643][5];				l_cell_reg[647] = inform_L[659][5];				l_cell_reg[648] = inform_L[644][5];				l_cell_reg[649] = inform_L[660][5];				l_cell_reg[650] = inform_L[645][5];				l_cell_reg[651] = inform_L[661][5];				l_cell_reg[652] = inform_L[646][5];				l_cell_reg[653] = inform_L[662][5];				l_cell_reg[654] = inform_L[647][5];				l_cell_reg[655] = inform_L[663][5];				l_cell_reg[656] = inform_L[648][5];				l_cell_reg[657] = inform_L[664][5];				l_cell_reg[658] = inform_L[649][5];				l_cell_reg[659] = inform_L[665][5];				l_cell_reg[660] = inform_L[650][5];				l_cell_reg[661] = inform_L[666][5];				l_cell_reg[662] = inform_L[651][5];				l_cell_reg[663] = inform_L[667][5];				l_cell_reg[664] = inform_L[652][5];				l_cell_reg[665] = inform_L[668][5];				l_cell_reg[666] = inform_L[653][5];				l_cell_reg[667] = inform_L[669][5];				l_cell_reg[668] = inform_L[654][5];				l_cell_reg[669] = inform_L[670][5];				l_cell_reg[670] = inform_L[655][5];				l_cell_reg[671] = inform_L[671][5];				l_cell_reg[672] = inform_L[672][5];				l_cell_reg[673] = inform_L[688][5];				l_cell_reg[674] = inform_L[673][5];				l_cell_reg[675] = inform_L[689][5];				l_cell_reg[676] = inform_L[674][5];				l_cell_reg[677] = inform_L[690][5];				l_cell_reg[678] = inform_L[675][5];				l_cell_reg[679] = inform_L[691][5];				l_cell_reg[680] = inform_L[676][5];				l_cell_reg[681] = inform_L[692][5];				l_cell_reg[682] = inform_L[677][5];				l_cell_reg[683] = inform_L[693][5];				l_cell_reg[684] = inform_L[678][5];				l_cell_reg[685] = inform_L[694][5];				l_cell_reg[686] = inform_L[679][5];				l_cell_reg[687] = inform_L[695][5];				l_cell_reg[688] = inform_L[680][5];				l_cell_reg[689] = inform_L[696][5];				l_cell_reg[690] = inform_L[681][5];				l_cell_reg[691] = inform_L[697][5];				l_cell_reg[692] = inform_L[682][5];				l_cell_reg[693] = inform_L[698][5];				l_cell_reg[694] = inform_L[683][5];				l_cell_reg[695] = inform_L[699][5];				l_cell_reg[696] = inform_L[684][5];				l_cell_reg[697] = inform_L[700][5];				l_cell_reg[698] = inform_L[685][5];				l_cell_reg[699] = inform_L[701][5];				l_cell_reg[700] = inform_L[686][5];				l_cell_reg[701] = inform_L[702][5];				l_cell_reg[702] = inform_L[687][5];				l_cell_reg[703] = inform_L[703][5];				l_cell_reg[704] = inform_L[704][5];				l_cell_reg[705] = inform_L[720][5];				l_cell_reg[706] = inform_L[705][5];				l_cell_reg[707] = inform_L[721][5];				l_cell_reg[708] = inform_L[706][5];				l_cell_reg[709] = inform_L[722][5];				l_cell_reg[710] = inform_L[707][5];				l_cell_reg[711] = inform_L[723][5];				l_cell_reg[712] = inform_L[708][5];				l_cell_reg[713] = inform_L[724][5];				l_cell_reg[714] = inform_L[709][5];				l_cell_reg[715] = inform_L[725][5];				l_cell_reg[716] = inform_L[710][5];				l_cell_reg[717] = inform_L[726][5];				l_cell_reg[718] = inform_L[711][5];				l_cell_reg[719] = inform_L[727][5];				l_cell_reg[720] = inform_L[712][5];				l_cell_reg[721] = inform_L[728][5];				l_cell_reg[722] = inform_L[713][5];				l_cell_reg[723] = inform_L[729][5];				l_cell_reg[724] = inform_L[714][5];				l_cell_reg[725] = inform_L[730][5];				l_cell_reg[726] = inform_L[715][5];				l_cell_reg[727] = inform_L[731][5];				l_cell_reg[728] = inform_L[716][5];				l_cell_reg[729] = inform_L[732][5];				l_cell_reg[730] = inform_L[717][5];				l_cell_reg[731] = inform_L[733][5];				l_cell_reg[732] = inform_L[718][5];				l_cell_reg[733] = inform_L[734][5];				l_cell_reg[734] = inform_L[719][5];				l_cell_reg[735] = inform_L[735][5];				l_cell_reg[736] = inform_L[736][5];				l_cell_reg[737] = inform_L[752][5];				l_cell_reg[738] = inform_L[737][5];				l_cell_reg[739] = inform_L[753][5];				l_cell_reg[740] = inform_L[738][5];				l_cell_reg[741] = inform_L[754][5];				l_cell_reg[742] = inform_L[739][5];				l_cell_reg[743] = inform_L[755][5];				l_cell_reg[744] = inform_L[740][5];				l_cell_reg[745] = inform_L[756][5];				l_cell_reg[746] = inform_L[741][5];				l_cell_reg[747] = inform_L[757][5];				l_cell_reg[748] = inform_L[742][5];				l_cell_reg[749] = inform_L[758][5];				l_cell_reg[750] = inform_L[743][5];				l_cell_reg[751] = inform_L[759][5];				l_cell_reg[752] = inform_L[744][5];				l_cell_reg[753] = inform_L[760][5];				l_cell_reg[754] = inform_L[745][5];				l_cell_reg[755] = inform_L[761][5];				l_cell_reg[756] = inform_L[746][5];				l_cell_reg[757] = inform_L[762][5];				l_cell_reg[758] = inform_L[747][5];				l_cell_reg[759] = inform_L[763][5];				l_cell_reg[760] = inform_L[748][5];				l_cell_reg[761] = inform_L[764][5];				l_cell_reg[762] = inform_L[749][5];				l_cell_reg[763] = inform_L[765][5];				l_cell_reg[764] = inform_L[750][5];				l_cell_reg[765] = inform_L[766][5];				l_cell_reg[766] = inform_L[751][5];				l_cell_reg[767] = inform_L[767][5];				l_cell_reg[768] = inform_L[768][5];				l_cell_reg[769] = inform_L[784][5];				l_cell_reg[770] = inform_L[769][5];				l_cell_reg[771] = inform_L[785][5];				l_cell_reg[772] = inform_L[770][5];				l_cell_reg[773] = inform_L[786][5];				l_cell_reg[774] = inform_L[771][5];				l_cell_reg[775] = inform_L[787][5];				l_cell_reg[776] = inform_L[772][5];				l_cell_reg[777] = inform_L[788][5];				l_cell_reg[778] = inform_L[773][5];				l_cell_reg[779] = inform_L[789][5];				l_cell_reg[780] = inform_L[774][5];				l_cell_reg[781] = inform_L[790][5];				l_cell_reg[782] = inform_L[775][5];				l_cell_reg[783] = inform_L[791][5];				l_cell_reg[784] = inform_L[776][5];				l_cell_reg[785] = inform_L[792][5];				l_cell_reg[786] = inform_L[777][5];				l_cell_reg[787] = inform_L[793][5];				l_cell_reg[788] = inform_L[778][5];				l_cell_reg[789] = inform_L[794][5];				l_cell_reg[790] = inform_L[779][5];				l_cell_reg[791] = inform_L[795][5];				l_cell_reg[792] = inform_L[780][5];				l_cell_reg[793] = inform_L[796][5];				l_cell_reg[794] = inform_L[781][5];				l_cell_reg[795] = inform_L[797][5];				l_cell_reg[796] = inform_L[782][5];				l_cell_reg[797] = inform_L[798][5];				l_cell_reg[798] = inform_L[783][5];				l_cell_reg[799] = inform_L[799][5];				l_cell_reg[800] = inform_L[800][5];				l_cell_reg[801] = inform_L[816][5];				l_cell_reg[802] = inform_L[801][5];				l_cell_reg[803] = inform_L[817][5];				l_cell_reg[804] = inform_L[802][5];				l_cell_reg[805] = inform_L[818][5];				l_cell_reg[806] = inform_L[803][5];				l_cell_reg[807] = inform_L[819][5];				l_cell_reg[808] = inform_L[804][5];				l_cell_reg[809] = inform_L[820][5];				l_cell_reg[810] = inform_L[805][5];				l_cell_reg[811] = inform_L[821][5];				l_cell_reg[812] = inform_L[806][5];				l_cell_reg[813] = inform_L[822][5];				l_cell_reg[814] = inform_L[807][5];				l_cell_reg[815] = inform_L[823][5];				l_cell_reg[816] = inform_L[808][5];				l_cell_reg[817] = inform_L[824][5];				l_cell_reg[818] = inform_L[809][5];				l_cell_reg[819] = inform_L[825][5];				l_cell_reg[820] = inform_L[810][5];				l_cell_reg[821] = inform_L[826][5];				l_cell_reg[822] = inform_L[811][5];				l_cell_reg[823] = inform_L[827][5];				l_cell_reg[824] = inform_L[812][5];				l_cell_reg[825] = inform_L[828][5];				l_cell_reg[826] = inform_L[813][5];				l_cell_reg[827] = inform_L[829][5];				l_cell_reg[828] = inform_L[814][5];				l_cell_reg[829] = inform_L[830][5];				l_cell_reg[830] = inform_L[815][5];				l_cell_reg[831] = inform_L[831][5];				l_cell_reg[832] = inform_L[832][5];				l_cell_reg[833] = inform_L[848][5];				l_cell_reg[834] = inform_L[833][5];				l_cell_reg[835] = inform_L[849][5];				l_cell_reg[836] = inform_L[834][5];				l_cell_reg[837] = inform_L[850][5];				l_cell_reg[838] = inform_L[835][5];				l_cell_reg[839] = inform_L[851][5];				l_cell_reg[840] = inform_L[836][5];				l_cell_reg[841] = inform_L[852][5];				l_cell_reg[842] = inform_L[837][5];				l_cell_reg[843] = inform_L[853][5];				l_cell_reg[844] = inform_L[838][5];				l_cell_reg[845] = inform_L[854][5];				l_cell_reg[846] = inform_L[839][5];				l_cell_reg[847] = inform_L[855][5];				l_cell_reg[848] = inform_L[840][5];				l_cell_reg[849] = inform_L[856][5];				l_cell_reg[850] = inform_L[841][5];				l_cell_reg[851] = inform_L[857][5];				l_cell_reg[852] = inform_L[842][5];				l_cell_reg[853] = inform_L[858][5];				l_cell_reg[854] = inform_L[843][5];				l_cell_reg[855] = inform_L[859][5];				l_cell_reg[856] = inform_L[844][5];				l_cell_reg[857] = inform_L[860][5];				l_cell_reg[858] = inform_L[845][5];				l_cell_reg[859] = inform_L[861][5];				l_cell_reg[860] = inform_L[846][5];				l_cell_reg[861] = inform_L[862][5];				l_cell_reg[862] = inform_L[847][5];				l_cell_reg[863] = inform_L[863][5];				l_cell_reg[864] = inform_L[864][5];				l_cell_reg[865] = inform_L[880][5];				l_cell_reg[866] = inform_L[865][5];				l_cell_reg[867] = inform_L[881][5];				l_cell_reg[868] = inform_L[866][5];				l_cell_reg[869] = inform_L[882][5];				l_cell_reg[870] = inform_L[867][5];				l_cell_reg[871] = inform_L[883][5];				l_cell_reg[872] = inform_L[868][5];				l_cell_reg[873] = inform_L[884][5];				l_cell_reg[874] = inform_L[869][5];				l_cell_reg[875] = inform_L[885][5];				l_cell_reg[876] = inform_L[870][5];				l_cell_reg[877] = inform_L[886][5];				l_cell_reg[878] = inform_L[871][5];				l_cell_reg[879] = inform_L[887][5];				l_cell_reg[880] = inform_L[872][5];				l_cell_reg[881] = inform_L[888][5];				l_cell_reg[882] = inform_L[873][5];				l_cell_reg[883] = inform_L[889][5];				l_cell_reg[884] = inform_L[874][5];				l_cell_reg[885] = inform_L[890][5];				l_cell_reg[886] = inform_L[875][5];				l_cell_reg[887] = inform_L[891][5];				l_cell_reg[888] = inform_L[876][5];				l_cell_reg[889] = inform_L[892][5];				l_cell_reg[890] = inform_L[877][5];				l_cell_reg[891] = inform_L[893][5];				l_cell_reg[892] = inform_L[878][5];				l_cell_reg[893] = inform_L[894][5];				l_cell_reg[894] = inform_L[879][5];				l_cell_reg[895] = inform_L[895][5];				l_cell_reg[896] = inform_L[896][5];				l_cell_reg[897] = inform_L[912][5];				l_cell_reg[898] = inform_L[897][5];				l_cell_reg[899] = inform_L[913][5];				l_cell_reg[900] = inform_L[898][5];				l_cell_reg[901] = inform_L[914][5];				l_cell_reg[902] = inform_L[899][5];				l_cell_reg[903] = inform_L[915][5];				l_cell_reg[904] = inform_L[900][5];				l_cell_reg[905] = inform_L[916][5];				l_cell_reg[906] = inform_L[901][5];				l_cell_reg[907] = inform_L[917][5];				l_cell_reg[908] = inform_L[902][5];				l_cell_reg[909] = inform_L[918][5];				l_cell_reg[910] = inform_L[903][5];				l_cell_reg[911] = inform_L[919][5];				l_cell_reg[912] = inform_L[904][5];				l_cell_reg[913] = inform_L[920][5];				l_cell_reg[914] = inform_L[905][5];				l_cell_reg[915] = inform_L[921][5];				l_cell_reg[916] = inform_L[906][5];				l_cell_reg[917] = inform_L[922][5];				l_cell_reg[918] = inform_L[907][5];				l_cell_reg[919] = inform_L[923][5];				l_cell_reg[920] = inform_L[908][5];				l_cell_reg[921] = inform_L[924][5];				l_cell_reg[922] = inform_L[909][5];				l_cell_reg[923] = inform_L[925][5];				l_cell_reg[924] = inform_L[910][5];				l_cell_reg[925] = inform_L[926][5];				l_cell_reg[926] = inform_L[911][5];				l_cell_reg[927] = inform_L[927][5];				l_cell_reg[928] = inform_L[928][5];				l_cell_reg[929] = inform_L[944][5];				l_cell_reg[930] = inform_L[929][5];				l_cell_reg[931] = inform_L[945][5];				l_cell_reg[932] = inform_L[930][5];				l_cell_reg[933] = inform_L[946][5];				l_cell_reg[934] = inform_L[931][5];				l_cell_reg[935] = inform_L[947][5];				l_cell_reg[936] = inform_L[932][5];				l_cell_reg[937] = inform_L[948][5];				l_cell_reg[938] = inform_L[933][5];				l_cell_reg[939] = inform_L[949][5];				l_cell_reg[940] = inform_L[934][5];				l_cell_reg[941] = inform_L[950][5];				l_cell_reg[942] = inform_L[935][5];				l_cell_reg[943] = inform_L[951][5];				l_cell_reg[944] = inform_L[936][5];				l_cell_reg[945] = inform_L[952][5];				l_cell_reg[946] = inform_L[937][5];				l_cell_reg[947] = inform_L[953][5];				l_cell_reg[948] = inform_L[938][5];				l_cell_reg[949] = inform_L[954][5];				l_cell_reg[950] = inform_L[939][5];				l_cell_reg[951] = inform_L[955][5];				l_cell_reg[952] = inform_L[940][5];				l_cell_reg[953] = inform_L[956][5];				l_cell_reg[954] = inform_L[941][5];				l_cell_reg[955] = inform_L[957][5];				l_cell_reg[956] = inform_L[942][5];				l_cell_reg[957] = inform_L[958][5];				l_cell_reg[958] = inform_L[943][5];				l_cell_reg[959] = inform_L[959][5];				l_cell_reg[960] = inform_L[960][5];				l_cell_reg[961] = inform_L[976][5];				l_cell_reg[962] = inform_L[961][5];				l_cell_reg[963] = inform_L[977][5];				l_cell_reg[964] = inform_L[962][5];				l_cell_reg[965] = inform_L[978][5];				l_cell_reg[966] = inform_L[963][5];				l_cell_reg[967] = inform_L[979][5];				l_cell_reg[968] = inform_L[964][5];				l_cell_reg[969] = inform_L[980][5];				l_cell_reg[970] = inform_L[965][5];				l_cell_reg[971] = inform_L[981][5];				l_cell_reg[972] = inform_L[966][5];				l_cell_reg[973] = inform_L[982][5];				l_cell_reg[974] = inform_L[967][5];				l_cell_reg[975] = inform_L[983][5];				l_cell_reg[976] = inform_L[968][5];				l_cell_reg[977] = inform_L[984][5];				l_cell_reg[978] = inform_L[969][5];				l_cell_reg[979] = inform_L[985][5];				l_cell_reg[980] = inform_L[970][5];				l_cell_reg[981] = inform_L[986][5];				l_cell_reg[982] = inform_L[971][5];				l_cell_reg[983] = inform_L[987][5];				l_cell_reg[984] = inform_L[972][5];				l_cell_reg[985] = inform_L[988][5];				l_cell_reg[986] = inform_L[973][5];				l_cell_reg[987] = inform_L[989][5];				l_cell_reg[988] = inform_L[974][5];				l_cell_reg[989] = inform_L[990][5];				l_cell_reg[990] = inform_L[975][5];				l_cell_reg[991] = inform_L[991][5];				l_cell_reg[992] = inform_L[992][5];				l_cell_reg[993] = inform_L[1008][5];				l_cell_reg[994] = inform_L[993][5];				l_cell_reg[995] = inform_L[1009][5];				l_cell_reg[996] = inform_L[994][5];				l_cell_reg[997] = inform_L[1010][5];				l_cell_reg[998] = inform_L[995][5];				l_cell_reg[999] = inform_L[1011][5];				l_cell_reg[1000] = inform_L[996][5];				l_cell_reg[1001] = inform_L[1012][5];				l_cell_reg[1002] = inform_L[997][5];				l_cell_reg[1003] = inform_L[1013][5];				l_cell_reg[1004] = inform_L[998][5];				l_cell_reg[1005] = inform_L[1014][5];				l_cell_reg[1006] = inform_L[999][5];				l_cell_reg[1007] = inform_L[1015][5];				l_cell_reg[1008] = inform_L[1000][5];				l_cell_reg[1009] = inform_L[1016][5];				l_cell_reg[1010] = inform_L[1001][5];				l_cell_reg[1011] = inform_L[1017][5];				l_cell_reg[1012] = inform_L[1002][5];				l_cell_reg[1013] = inform_L[1018][5];				l_cell_reg[1014] = inform_L[1003][5];				l_cell_reg[1015] = inform_L[1019][5];				l_cell_reg[1016] = inform_L[1004][5];				l_cell_reg[1017] = inform_L[1020][5];				l_cell_reg[1018] = inform_L[1005][5];				l_cell_reg[1019] = inform_L[1021][5];				l_cell_reg[1020] = inform_L[1006][5];				l_cell_reg[1021] = inform_L[1022][5];				l_cell_reg[1022] = inform_L[1007][5];				l_cell_reg[1023] = inform_L[1023][5];			end
			6:			begin				r_cell_reg[0] = inform_R[0][5];				r_cell_reg[1] = inform_R[32][5];				r_cell_reg[2] = inform_R[1][5];				r_cell_reg[3] = inform_R[33][5];				r_cell_reg[4] = inform_R[2][5];				r_cell_reg[5] = inform_R[34][5];				r_cell_reg[6] = inform_R[3][5];				r_cell_reg[7] = inform_R[35][5];				r_cell_reg[8] = inform_R[4][5];				r_cell_reg[9] = inform_R[36][5];				r_cell_reg[10] = inform_R[5][5];				r_cell_reg[11] = inform_R[37][5];				r_cell_reg[12] = inform_R[6][5];				r_cell_reg[13] = inform_R[38][5];				r_cell_reg[14] = inform_R[7][5];				r_cell_reg[15] = inform_R[39][5];				r_cell_reg[16] = inform_R[8][5];				r_cell_reg[17] = inform_R[40][5];				r_cell_reg[18] = inform_R[9][5];				r_cell_reg[19] = inform_R[41][5];				r_cell_reg[20] = inform_R[10][5];				r_cell_reg[21] = inform_R[42][5];				r_cell_reg[22] = inform_R[11][5];				r_cell_reg[23] = inform_R[43][5];				r_cell_reg[24] = inform_R[12][5];				r_cell_reg[25] = inform_R[44][5];				r_cell_reg[26] = inform_R[13][5];				r_cell_reg[27] = inform_R[45][5];				r_cell_reg[28] = inform_R[14][5];				r_cell_reg[29] = inform_R[46][5];				r_cell_reg[30] = inform_R[15][5];				r_cell_reg[31] = inform_R[47][5];				r_cell_reg[32] = inform_R[16][5];				r_cell_reg[33] = inform_R[48][5];				r_cell_reg[34] = inform_R[17][5];				r_cell_reg[35] = inform_R[49][5];				r_cell_reg[36] = inform_R[18][5];				r_cell_reg[37] = inform_R[50][5];				r_cell_reg[38] = inform_R[19][5];				r_cell_reg[39] = inform_R[51][5];				r_cell_reg[40] = inform_R[20][5];				r_cell_reg[41] = inform_R[52][5];				r_cell_reg[42] = inform_R[21][5];				r_cell_reg[43] = inform_R[53][5];				r_cell_reg[44] = inform_R[22][5];				r_cell_reg[45] = inform_R[54][5];				r_cell_reg[46] = inform_R[23][5];				r_cell_reg[47] = inform_R[55][5];				r_cell_reg[48] = inform_R[24][5];				r_cell_reg[49] = inform_R[56][5];				r_cell_reg[50] = inform_R[25][5];				r_cell_reg[51] = inform_R[57][5];				r_cell_reg[52] = inform_R[26][5];				r_cell_reg[53] = inform_R[58][5];				r_cell_reg[54] = inform_R[27][5];				r_cell_reg[55] = inform_R[59][5];				r_cell_reg[56] = inform_R[28][5];				r_cell_reg[57] = inform_R[60][5];				r_cell_reg[58] = inform_R[29][5];				r_cell_reg[59] = inform_R[61][5];				r_cell_reg[60] = inform_R[30][5];				r_cell_reg[61] = inform_R[62][5];				r_cell_reg[62] = inform_R[31][5];				r_cell_reg[63] = inform_R[63][5];				r_cell_reg[64] = inform_R[64][5];				r_cell_reg[65] = inform_R[96][5];				r_cell_reg[66] = inform_R[65][5];				r_cell_reg[67] = inform_R[97][5];				r_cell_reg[68] = inform_R[66][5];				r_cell_reg[69] = inform_R[98][5];				r_cell_reg[70] = inform_R[67][5];				r_cell_reg[71] = inform_R[99][5];				r_cell_reg[72] = inform_R[68][5];				r_cell_reg[73] = inform_R[100][5];				r_cell_reg[74] = inform_R[69][5];				r_cell_reg[75] = inform_R[101][5];				r_cell_reg[76] = inform_R[70][5];				r_cell_reg[77] = inform_R[102][5];				r_cell_reg[78] = inform_R[71][5];				r_cell_reg[79] = inform_R[103][5];				r_cell_reg[80] = inform_R[72][5];				r_cell_reg[81] = inform_R[104][5];				r_cell_reg[82] = inform_R[73][5];				r_cell_reg[83] = inform_R[105][5];				r_cell_reg[84] = inform_R[74][5];				r_cell_reg[85] = inform_R[106][5];				r_cell_reg[86] = inform_R[75][5];				r_cell_reg[87] = inform_R[107][5];				r_cell_reg[88] = inform_R[76][5];				r_cell_reg[89] = inform_R[108][5];				r_cell_reg[90] = inform_R[77][5];				r_cell_reg[91] = inform_R[109][5];				r_cell_reg[92] = inform_R[78][5];				r_cell_reg[93] = inform_R[110][5];				r_cell_reg[94] = inform_R[79][5];				r_cell_reg[95] = inform_R[111][5];				r_cell_reg[96] = inform_R[80][5];				r_cell_reg[97] = inform_R[112][5];				r_cell_reg[98] = inform_R[81][5];				r_cell_reg[99] = inform_R[113][5];				r_cell_reg[100] = inform_R[82][5];				r_cell_reg[101] = inform_R[114][5];				r_cell_reg[102] = inform_R[83][5];				r_cell_reg[103] = inform_R[115][5];				r_cell_reg[104] = inform_R[84][5];				r_cell_reg[105] = inform_R[116][5];				r_cell_reg[106] = inform_R[85][5];				r_cell_reg[107] = inform_R[117][5];				r_cell_reg[108] = inform_R[86][5];				r_cell_reg[109] = inform_R[118][5];				r_cell_reg[110] = inform_R[87][5];				r_cell_reg[111] = inform_R[119][5];				r_cell_reg[112] = inform_R[88][5];				r_cell_reg[113] = inform_R[120][5];				r_cell_reg[114] = inform_R[89][5];				r_cell_reg[115] = inform_R[121][5];				r_cell_reg[116] = inform_R[90][5];				r_cell_reg[117] = inform_R[122][5];				r_cell_reg[118] = inform_R[91][5];				r_cell_reg[119] = inform_R[123][5];				r_cell_reg[120] = inform_R[92][5];				r_cell_reg[121] = inform_R[124][5];				r_cell_reg[122] = inform_R[93][5];				r_cell_reg[123] = inform_R[125][5];				r_cell_reg[124] = inform_R[94][5];				r_cell_reg[125] = inform_R[126][5];				r_cell_reg[126] = inform_R[95][5];				r_cell_reg[127] = inform_R[127][5];				r_cell_reg[128] = inform_R[128][5];				r_cell_reg[129] = inform_R[160][5];				r_cell_reg[130] = inform_R[129][5];				r_cell_reg[131] = inform_R[161][5];				r_cell_reg[132] = inform_R[130][5];				r_cell_reg[133] = inform_R[162][5];				r_cell_reg[134] = inform_R[131][5];				r_cell_reg[135] = inform_R[163][5];				r_cell_reg[136] = inform_R[132][5];				r_cell_reg[137] = inform_R[164][5];				r_cell_reg[138] = inform_R[133][5];				r_cell_reg[139] = inform_R[165][5];				r_cell_reg[140] = inform_R[134][5];				r_cell_reg[141] = inform_R[166][5];				r_cell_reg[142] = inform_R[135][5];				r_cell_reg[143] = inform_R[167][5];				r_cell_reg[144] = inform_R[136][5];				r_cell_reg[145] = inform_R[168][5];				r_cell_reg[146] = inform_R[137][5];				r_cell_reg[147] = inform_R[169][5];				r_cell_reg[148] = inform_R[138][5];				r_cell_reg[149] = inform_R[170][5];				r_cell_reg[150] = inform_R[139][5];				r_cell_reg[151] = inform_R[171][5];				r_cell_reg[152] = inform_R[140][5];				r_cell_reg[153] = inform_R[172][5];				r_cell_reg[154] = inform_R[141][5];				r_cell_reg[155] = inform_R[173][5];				r_cell_reg[156] = inform_R[142][5];				r_cell_reg[157] = inform_R[174][5];				r_cell_reg[158] = inform_R[143][5];				r_cell_reg[159] = inform_R[175][5];				r_cell_reg[160] = inform_R[144][5];				r_cell_reg[161] = inform_R[176][5];				r_cell_reg[162] = inform_R[145][5];				r_cell_reg[163] = inform_R[177][5];				r_cell_reg[164] = inform_R[146][5];				r_cell_reg[165] = inform_R[178][5];				r_cell_reg[166] = inform_R[147][5];				r_cell_reg[167] = inform_R[179][5];				r_cell_reg[168] = inform_R[148][5];				r_cell_reg[169] = inform_R[180][5];				r_cell_reg[170] = inform_R[149][5];				r_cell_reg[171] = inform_R[181][5];				r_cell_reg[172] = inform_R[150][5];				r_cell_reg[173] = inform_R[182][5];				r_cell_reg[174] = inform_R[151][5];				r_cell_reg[175] = inform_R[183][5];				r_cell_reg[176] = inform_R[152][5];				r_cell_reg[177] = inform_R[184][5];				r_cell_reg[178] = inform_R[153][5];				r_cell_reg[179] = inform_R[185][5];				r_cell_reg[180] = inform_R[154][5];				r_cell_reg[181] = inform_R[186][5];				r_cell_reg[182] = inform_R[155][5];				r_cell_reg[183] = inform_R[187][5];				r_cell_reg[184] = inform_R[156][5];				r_cell_reg[185] = inform_R[188][5];				r_cell_reg[186] = inform_R[157][5];				r_cell_reg[187] = inform_R[189][5];				r_cell_reg[188] = inform_R[158][5];				r_cell_reg[189] = inform_R[190][5];				r_cell_reg[190] = inform_R[159][5];				r_cell_reg[191] = inform_R[191][5];				r_cell_reg[192] = inform_R[192][5];				r_cell_reg[193] = inform_R[224][5];				r_cell_reg[194] = inform_R[193][5];				r_cell_reg[195] = inform_R[225][5];				r_cell_reg[196] = inform_R[194][5];				r_cell_reg[197] = inform_R[226][5];				r_cell_reg[198] = inform_R[195][5];				r_cell_reg[199] = inform_R[227][5];				r_cell_reg[200] = inform_R[196][5];				r_cell_reg[201] = inform_R[228][5];				r_cell_reg[202] = inform_R[197][5];				r_cell_reg[203] = inform_R[229][5];				r_cell_reg[204] = inform_R[198][5];				r_cell_reg[205] = inform_R[230][5];				r_cell_reg[206] = inform_R[199][5];				r_cell_reg[207] = inform_R[231][5];				r_cell_reg[208] = inform_R[200][5];				r_cell_reg[209] = inform_R[232][5];				r_cell_reg[210] = inform_R[201][5];				r_cell_reg[211] = inform_R[233][5];				r_cell_reg[212] = inform_R[202][5];				r_cell_reg[213] = inform_R[234][5];				r_cell_reg[214] = inform_R[203][5];				r_cell_reg[215] = inform_R[235][5];				r_cell_reg[216] = inform_R[204][5];				r_cell_reg[217] = inform_R[236][5];				r_cell_reg[218] = inform_R[205][5];				r_cell_reg[219] = inform_R[237][5];				r_cell_reg[220] = inform_R[206][5];				r_cell_reg[221] = inform_R[238][5];				r_cell_reg[222] = inform_R[207][5];				r_cell_reg[223] = inform_R[239][5];				r_cell_reg[224] = inform_R[208][5];				r_cell_reg[225] = inform_R[240][5];				r_cell_reg[226] = inform_R[209][5];				r_cell_reg[227] = inform_R[241][5];				r_cell_reg[228] = inform_R[210][5];				r_cell_reg[229] = inform_R[242][5];				r_cell_reg[230] = inform_R[211][5];				r_cell_reg[231] = inform_R[243][5];				r_cell_reg[232] = inform_R[212][5];				r_cell_reg[233] = inform_R[244][5];				r_cell_reg[234] = inform_R[213][5];				r_cell_reg[235] = inform_R[245][5];				r_cell_reg[236] = inform_R[214][5];				r_cell_reg[237] = inform_R[246][5];				r_cell_reg[238] = inform_R[215][5];				r_cell_reg[239] = inform_R[247][5];				r_cell_reg[240] = inform_R[216][5];				r_cell_reg[241] = inform_R[248][5];				r_cell_reg[242] = inform_R[217][5];				r_cell_reg[243] = inform_R[249][5];				r_cell_reg[244] = inform_R[218][5];				r_cell_reg[245] = inform_R[250][5];				r_cell_reg[246] = inform_R[219][5];				r_cell_reg[247] = inform_R[251][5];				r_cell_reg[248] = inform_R[220][5];				r_cell_reg[249] = inform_R[252][5];				r_cell_reg[250] = inform_R[221][5];				r_cell_reg[251] = inform_R[253][5];				r_cell_reg[252] = inform_R[222][5];				r_cell_reg[253] = inform_R[254][5];				r_cell_reg[254] = inform_R[223][5];				r_cell_reg[255] = inform_R[255][5];				r_cell_reg[256] = inform_R[256][5];				r_cell_reg[257] = inform_R[288][5];				r_cell_reg[258] = inform_R[257][5];				r_cell_reg[259] = inform_R[289][5];				r_cell_reg[260] = inform_R[258][5];				r_cell_reg[261] = inform_R[290][5];				r_cell_reg[262] = inform_R[259][5];				r_cell_reg[263] = inform_R[291][5];				r_cell_reg[264] = inform_R[260][5];				r_cell_reg[265] = inform_R[292][5];				r_cell_reg[266] = inform_R[261][5];				r_cell_reg[267] = inform_R[293][5];				r_cell_reg[268] = inform_R[262][5];				r_cell_reg[269] = inform_R[294][5];				r_cell_reg[270] = inform_R[263][5];				r_cell_reg[271] = inform_R[295][5];				r_cell_reg[272] = inform_R[264][5];				r_cell_reg[273] = inform_R[296][5];				r_cell_reg[274] = inform_R[265][5];				r_cell_reg[275] = inform_R[297][5];				r_cell_reg[276] = inform_R[266][5];				r_cell_reg[277] = inform_R[298][5];				r_cell_reg[278] = inform_R[267][5];				r_cell_reg[279] = inform_R[299][5];				r_cell_reg[280] = inform_R[268][5];				r_cell_reg[281] = inform_R[300][5];				r_cell_reg[282] = inform_R[269][5];				r_cell_reg[283] = inform_R[301][5];				r_cell_reg[284] = inform_R[270][5];				r_cell_reg[285] = inform_R[302][5];				r_cell_reg[286] = inform_R[271][5];				r_cell_reg[287] = inform_R[303][5];				r_cell_reg[288] = inform_R[272][5];				r_cell_reg[289] = inform_R[304][5];				r_cell_reg[290] = inform_R[273][5];				r_cell_reg[291] = inform_R[305][5];				r_cell_reg[292] = inform_R[274][5];				r_cell_reg[293] = inform_R[306][5];				r_cell_reg[294] = inform_R[275][5];				r_cell_reg[295] = inform_R[307][5];				r_cell_reg[296] = inform_R[276][5];				r_cell_reg[297] = inform_R[308][5];				r_cell_reg[298] = inform_R[277][5];				r_cell_reg[299] = inform_R[309][5];				r_cell_reg[300] = inform_R[278][5];				r_cell_reg[301] = inform_R[310][5];				r_cell_reg[302] = inform_R[279][5];				r_cell_reg[303] = inform_R[311][5];				r_cell_reg[304] = inform_R[280][5];				r_cell_reg[305] = inform_R[312][5];				r_cell_reg[306] = inform_R[281][5];				r_cell_reg[307] = inform_R[313][5];				r_cell_reg[308] = inform_R[282][5];				r_cell_reg[309] = inform_R[314][5];				r_cell_reg[310] = inform_R[283][5];				r_cell_reg[311] = inform_R[315][5];				r_cell_reg[312] = inform_R[284][5];				r_cell_reg[313] = inform_R[316][5];				r_cell_reg[314] = inform_R[285][5];				r_cell_reg[315] = inform_R[317][5];				r_cell_reg[316] = inform_R[286][5];				r_cell_reg[317] = inform_R[318][5];				r_cell_reg[318] = inform_R[287][5];				r_cell_reg[319] = inform_R[319][5];				r_cell_reg[320] = inform_R[320][5];				r_cell_reg[321] = inform_R[352][5];				r_cell_reg[322] = inform_R[321][5];				r_cell_reg[323] = inform_R[353][5];				r_cell_reg[324] = inform_R[322][5];				r_cell_reg[325] = inform_R[354][5];				r_cell_reg[326] = inform_R[323][5];				r_cell_reg[327] = inform_R[355][5];				r_cell_reg[328] = inform_R[324][5];				r_cell_reg[329] = inform_R[356][5];				r_cell_reg[330] = inform_R[325][5];				r_cell_reg[331] = inform_R[357][5];				r_cell_reg[332] = inform_R[326][5];				r_cell_reg[333] = inform_R[358][5];				r_cell_reg[334] = inform_R[327][5];				r_cell_reg[335] = inform_R[359][5];				r_cell_reg[336] = inform_R[328][5];				r_cell_reg[337] = inform_R[360][5];				r_cell_reg[338] = inform_R[329][5];				r_cell_reg[339] = inform_R[361][5];				r_cell_reg[340] = inform_R[330][5];				r_cell_reg[341] = inform_R[362][5];				r_cell_reg[342] = inform_R[331][5];				r_cell_reg[343] = inform_R[363][5];				r_cell_reg[344] = inform_R[332][5];				r_cell_reg[345] = inform_R[364][5];				r_cell_reg[346] = inform_R[333][5];				r_cell_reg[347] = inform_R[365][5];				r_cell_reg[348] = inform_R[334][5];				r_cell_reg[349] = inform_R[366][5];				r_cell_reg[350] = inform_R[335][5];				r_cell_reg[351] = inform_R[367][5];				r_cell_reg[352] = inform_R[336][5];				r_cell_reg[353] = inform_R[368][5];				r_cell_reg[354] = inform_R[337][5];				r_cell_reg[355] = inform_R[369][5];				r_cell_reg[356] = inform_R[338][5];				r_cell_reg[357] = inform_R[370][5];				r_cell_reg[358] = inform_R[339][5];				r_cell_reg[359] = inform_R[371][5];				r_cell_reg[360] = inform_R[340][5];				r_cell_reg[361] = inform_R[372][5];				r_cell_reg[362] = inform_R[341][5];				r_cell_reg[363] = inform_R[373][5];				r_cell_reg[364] = inform_R[342][5];				r_cell_reg[365] = inform_R[374][5];				r_cell_reg[366] = inform_R[343][5];				r_cell_reg[367] = inform_R[375][5];				r_cell_reg[368] = inform_R[344][5];				r_cell_reg[369] = inform_R[376][5];				r_cell_reg[370] = inform_R[345][5];				r_cell_reg[371] = inform_R[377][5];				r_cell_reg[372] = inform_R[346][5];				r_cell_reg[373] = inform_R[378][5];				r_cell_reg[374] = inform_R[347][5];				r_cell_reg[375] = inform_R[379][5];				r_cell_reg[376] = inform_R[348][5];				r_cell_reg[377] = inform_R[380][5];				r_cell_reg[378] = inform_R[349][5];				r_cell_reg[379] = inform_R[381][5];				r_cell_reg[380] = inform_R[350][5];				r_cell_reg[381] = inform_R[382][5];				r_cell_reg[382] = inform_R[351][5];				r_cell_reg[383] = inform_R[383][5];				r_cell_reg[384] = inform_R[384][5];				r_cell_reg[385] = inform_R[416][5];				r_cell_reg[386] = inform_R[385][5];				r_cell_reg[387] = inform_R[417][5];				r_cell_reg[388] = inform_R[386][5];				r_cell_reg[389] = inform_R[418][5];				r_cell_reg[390] = inform_R[387][5];				r_cell_reg[391] = inform_R[419][5];				r_cell_reg[392] = inform_R[388][5];				r_cell_reg[393] = inform_R[420][5];				r_cell_reg[394] = inform_R[389][5];				r_cell_reg[395] = inform_R[421][5];				r_cell_reg[396] = inform_R[390][5];				r_cell_reg[397] = inform_R[422][5];				r_cell_reg[398] = inform_R[391][5];				r_cell_reg[399] = inform_R[423][5];				r_cell_reg[400] = inform_R[392][5];				r_cell_reg[401] = inform_R[424][5];				r_cell_reg[402] = inform_R[393][5];				r_cell_reg[403] = inform_R[425][5];				r_cell_reg[404] = inform_R[394][5];				r_cell_reg[405] = inform_R[426][5];				r_cell_reg[406] = inform_R[395][5];				r_cell_reg[407] = inform_R[427][5];				r_cell_reg[408] = inform_R[396][5];				r_cell_reg[409] = inform_R[428][5];				r_cell_reg[410] = inform_R[397][5];				r_cell_reg[411] = inform_R[429][5];				r_cell_reg[412] = inform_R[398][5];				r_cell_reg[413] = inform_R[430][5];				r_cell_reg[414] = inform_R[399][5];				r_cell_reg[415] = inform_R[431][5];				r_cell_reg[416] = inform_R[400][5];				r_cell_reg[417] = inform_R[432][5];				r_cell_reg[418] = inform_R[401][5];				r_cell_reg[419] = inform_R[433][5];				r_cell_reg[420] = inform_R[402][5];				r_cell_reg[421] = inform_R[434][5];				r_cell_reg[422] = inform_R[403][5];				r_cell_reg[423] = inform_R[435][5];				r_cell_reg[424] = inform_R[404][5];				r_cell_reg[425] = inform_R[436][5];				r_cell_reg[426] = inform_R[405][5];				r_cell_reg[427] = inform_R[437][5];				r_cell_reg[428] = inform_R[406][5];				r_cell_reg[429] = inform_R[438][5];				r_cell_reg[430] = inform_R[407][5];				r_cell_reg[431] = inform_R[439][5];				r_cell_reg[432] = inform_R[408][5];				r_cell_reg[433] = inform_R[440][5];				r_cell_reg[434] = inform_R[409][5];				r_cell_reg[435] = inform_R[441][5];				r_cell_reg[436] = inform_R[410][5];				r_cell_reg[437] = inform_R[442][5];				r_cell_reg[438] = inform_R[411][5];				r_cell_reg[439] = inform_R[443][5];				r_cell_reg[440] = inform_R[412][5];				r_cell_reg[441] = inform_R[444][5];				r_cell_reg[442] = inform_R[413][5];				r_cell_reg[443] = inform_R[445][5];				r_cell_reg[444] = inform_R[414][5];				r_cell_reg[445] = inform_R[446][5];				r_cell_reg[446] = inform_R[415][5];				r_cell_reg[447] = inform_R[447][5];				r_cell_reg[448] = inform_R[448][5];				r_cell_reg[449] = inform_R[480][5];				r_cell_reg[450] = inform_R[449][5];				r_cell_reg[451] = inform_R[481][5];				r_cell_reg[452] = inform_R[450][5];				r_cell_reg[453] = inform_R[482][5];				r_cell_reg[454] = inform_R[451][5];				r_cell_reg[455] = inform_R[483][5];				r_cell_reg[456] = inform_R[452][5];				r_cell_reg[457] = inform_R[484][5];				r_cell_reg[458] = inform_R[453][5];				r_cell_reg[459] = inform_R[485][5];				r_cell_reg[460] = inform_R[454][5];				r_cell_reg[461] = inform_R[486][5];				r_cell_reg[462] = inform_R[455][5];				r_cell_reg[463] = inform_R[487][5];				r_cell_reg[464] = inform_R[456][5];				r_cell_reg[465] = inform_R[488][5];				r_cell_reg[466] = inform_R[457][5];				r_cell_reg[467] = inform_R[489][5];				r_cell_reg[468] = inform_R[458][5];				r_cell_reg[469] = inform_R[490][5];				r_cell_reg[470] = inform_R[459][5];				r_cell_reg[471] = inform_R[491][5];				r_cell_reg[472] = inform_R[460][5];				r_cell_reg[473] = inform_R[492][5];				r_cell_reg[474] = inform_R[461][5];				r_cell_reg[475] = inform_R[493][5];				r_cell_reg[476] = inform_R[462][5];				r_cell_reg[477] = inform_R[494][5];				r_cell_reg[478] = inform_R[463][5];				r_cell_reg[479] = inform_R[495][5];				r_cell_reg[480] = inform_R[464][5];				r_cell_reg[481] = inform_R[496][5];				r_cell_reg[482] = inform_R[465][5];				r_cell_reg[483] = inform_R[497][5];				r_cell_reg[484] = inform_R[466][5];				r_cell_reg[485] = inform_R[498][5];				r_cell_reg[486] = inform_R[467][5];				r_cell_reg[487] = inform_R[499][5];				r_cell_reg[488] = inform_R[468][5];				r_cell_reg[489] = inform_R[500][5];				r_cell_reg[490] = inform_R[469][5];				r_cell_reg[491] = inform_R[501][5];				r_cell_reg[492] = inform_R[470][5];				r_cell_reg[493] = inform_R[502][5];				r_cell_reg[494] = inform_R[471][5];				r_cell_reg[495] = inform_R[503][5];				r_cell_reg[496] = inform_R[472][5];				r_cell_reg[497] = inform_R[504][5];				r_cell_reg[498] = inform_R[473][5];				r_cell_reg[499] = inform_R[505][5];				r_cell_reg[500] = inform_R[474][5];				r_cell_reg[501] = inform_R[506][5];				r_cell_reg[502] = inform_R[475][5];				r_cell_reg[503] = inform_R[507][5];				r_cell_reg[504] = inform_R[476][5];				r_cell_reg[505] = inform_R[508][5];				r_cell_reg[506] = inform_R[477][5];				r_cell_reg[507] = inform_R[509][5];				r_cell_reg[508] = inform_R[478][5];				r_cell_reg[509] = inform_R[510][5];				r_cell_reg[510] = inform_R[479][5];				r_cell_reg[511] = inform_R[511][5];				r_cell_reg[512] = inform_R[512][5];				r_cell_reg[513] = inform_R[544][5];				r_cell_reg[514] = inform_R[513][5];				r_cell_reg[515] = inform_R[545][5];				r_cell_reg[516] = inform_R[514][5];				r_cell_reg[517] = inform_R[546][5];				r_cell_reg[518] = inform_R[515][5];				r_cell_reg[519] = inform_R[547][5];				r_cell_reg[520] = inform_R[516][5];				r_cell_reg[521] = inform_R[548][5];				r_cell_reg[522] = inform_R[517][5];				r_cell_reg[523] = inform_R[549][5];				r_cell_reg[524] = inform_R[518][5];				r_cell_reg[525] = inform_R[550][5];				r_cell_reg[526] = inform_R[519][5];				r_cell_reg[527] = inform_R[551][5];				r_cell_reg[528] = inform_R[520][5];				r_cell_reg[529] = inform_R[552][5];				r_cell_reg[530] = inform_R[521][5];				r_cell_reg[531] = inform_R[553][5];				r_cell_reg[532] = inform_R[522][5];				r_cell_reg[533] = inform_R[554][5];				r_cell_reg[534] = inform_R[523][5];				r_cell_reg[535] = inform_R[555][5];				r_cell_reg[536] = inform_R[524][5];				r_cell_reg[537] = inform_R[556][5];				r_cell_reg[538] = inform_R[525][5];				r_cell_reg[539] = inform_R[557][5];				r_cell_reg[540] = inform_R[526][5];				r_cell_reg[541] = inform_R[558][5];				r_cell_reg[542] = inform_R[527][5];				r_cell_reg[543] = inform_R[559][5];				r_cell_reg[544] = inform_R[528][5];				r_cell_reg[545] = inform_R[560][5];				r_cell_reg[546] = inform_R[529][5];				r_cell_reg[547] = inform_R[561][5];				r_cell_reg[548] = inform_R[530][5];				r_cell_reg[549] = inform_R[562][5];				r_cell_reg[550] = inform_R[531][5];				r_cell_reg[551] = inform_R[563][5];				r_cell_reg[552] = inform_R[532][5];				r_cell_reg[553] = inform_R[564][5];				r_cell_reg[554] = inform_R[533][5];				r_cell_reg[555] = inform_R[565][5];				r_cell_reg[556] = inform_R[534][5];				r_cell_reg[557] = inform_R[566][5];				r_cell_reg[558] = inform_R[535][5];				r_cell_reg[559] = inform_R[567][5];				r_cell_reg[560] = inform_R[536][5];				r_cell_reg[561] = inform_R[568][5];				r_cell_reg[562] = inform_R[537][5];				r_cell_reg[563] = inform_R[569][5];				r_cell_reg[564] = inform_R[538][5];				r_cell_reg[565] = inform_R[570][5];				r_cell_reg[566] = inform_R[539][5];				r_cell_reg[567] = inform_R[571][5];				r_cell_reg[568] = inform_R[540][5];				r_cell_reg[569] = inform_R[572][5];				r_cell_reg[570] = inform_R[541][5];				r_cell_reg[571] = inform_R[573][5];				r_cell_reg[572] = inform_R[542][5];				r_cell_reg[573] = inform_R[574][5];				r_cell_reg[574] = inform_R[543][5];				r_cell_reg[575] = inform_R[575][5];				r_cell_reg[576] = inform_R[576][5];				r_cell_reg[577] = inform_R[608][5];				r_cell_reg[578] = inform_R[577][5];				r_cell_reg[579] = inform_R[609][5];				r_cell_reg[580] = inform_R[578][5];				r_cell_reg[581] = inform_R[610][5];				r_cell_reg[582] = inform_R[579][5];				r_cell_reg[583] = inform_R[611][5];				r_cell_reg[584] = inform_R[580][5];				r_cell_reg[585] = inform_R[612][5];				r_cell_reg[586] = inform_R[581][5];				r_cell_reg[587] = inform_R[613][5];				r_cell_reg[588] = inform_R[582][5];				r_cell_reg[589] = inform_R[614][5];				r_cell_reg[590] = inform_R[583][5];				r_cell_reg[591] = inform_R[615][5];				r_cell_reg[592] = inform_R[584][5];				r_cell_reg[593] = inform_R[616][5];				r_cell_reg[594] = inform_R[585][5];				r_cell_reg[595] = inform_R[617][5];				r_cell_reg[596] = inform_R[586][5];				r_cell_reg[597] = inform_R[618][5];				r_cell_reg[598] = inform_R[587][5];				r_cell_reg[599] = inform_R[619][5];				r_cell_reg[600] = inform_R[588][5];				r_cell_reg[601] = inform_R[620][5];				r_cell_reg[602] = inform_R[589][5];				r_cell_reg[603] = inform_R[621][5];				r_cell_reg[604] = inform_R[590][5];				r_cell_reg[605] = inform_R[622][5];				r_cell_reg[606] = inform_R[591][5];				r_cell_reg[607] = inform_R[623][5];				r_cell_reg[608] = inform_R[592][5];				r_cell_reg[609] = inform_R[624][5];				r_cell_reg[610] = inform_R[593][5];				r_cell_reg[611] = inform_R[625][5];				r_cell_reg[612] = inform_R[594][5];				r_cell_reg[613] = inform_R[626][5];				r_cell_reg[614] = inform_R[595][5];				r_cell_reg[615] = inform_R[627][5];				r_cell_reg[616] = inform_R[596][5];				r_cell_reg[617] = inform_R[628][5];				r_cell_reg[618] = inform_R[597][5];				r_cell_reg[619] = inform_R[629][5];				r_cell_reg[620] = inform_R[598][5];				r_cell_reg[621] = inform_R[630][5];				r_cell_reg[622] = inform_R[599][5];				r_cell_reg[623] = inform_R[631][5];				r_cell_reg[624] = inform_R[600][5];				r_cell_reg[625] = inform_R[632][5];				r_cell_reg[626] = inform_R[601][5];				r_cell_reg[627] = inform_R[633][5];				r_cell_reg[628] = inform_R[602][5];				r_cell_reg[629] = inform_R[634][5];				r_cell_reg[630] = inform_R[603][5];				r_cell_reg[631] = inform_R[635][5];				r_cell_reg[632] = inform_R[604][5];				r_cell_reg[633] = inform_R[636][5];				r_cell_reg[634] = inform_R[605][5];				r_cell_reg[635] = inform_R[637][5];				r_cell_reg[636] = inform_R[606][5];				r_cell_reg[637] = inform_R[638][5];				r_cell_reg[638] = inform_R[607][5];				r_cell_reg[639] = inform_R[639][5];				r_cell_reg[640] = inform_R[640][5];				r_cell_reg[641] = inform_R[672][5];				r_cell_reg[642] = inform_R[641][5];				r_cell_reg[643] = inform_R[673][5];				r_cell_reg[644] = inform_R[642][5];				r_cell_reg[645] = inform_R[674][5];				r_cell_reg[646] = inform_R[643][5];				r_cell_reg[647] = inform_R[675][5];				r_cell_reg[648] = inform_R[644][5];				r_cell_reg[649] = inform_R[676][5];				r_cell_reg[650] = inform_R[645][5];				r_cell_reg[651] = inform_R[677][5];				r_cell_reg[652] = inform_R[646][5];				r_cell_reg[653] = inform_R[678][5];				r_cell_reg[654] = inform_R[647][5];				r_cell_reg[655] = inform_R[679][5];				r_cell_reg[656] = inform_R[648][5];				r_cell_reg[657] = inform_R[680][5];				r_cell_reg[658] = inform_R[649][5];				r_cell_reg[659] = inform_R[681][5];				r_cell_reg[660] = inform_R[650][5];				r_cell_reg[661] = inform_R[682][5];				r_cell_reg[662] = inform_R[651][5];				r_cell_reg[663] = inform_R[683][5];				r_cell_reg[664] = inform_R[652][5];				r_cell_reg[665] = inform_R[684][5];				r_cell_reg[666] = inform_R[653][5];				r_cell_reg[667] = inform_R[685][5];				r_cell_reg[668] = inform_R[654][5];				r_cell_reg[669] = inform_R[686][5];				r_cell_reg[670] = inform_R[655][5];				r_cell_reg[671] = inform_R[687][5];				r_cell_reg[672] = inform_R[656][5];				r_cell_reg[673] = inform_R[688][5];				r_cell_reg[674] = inform_R[657][5];				r_cell_reg[675] = inform_R[689][5];				r_cell_reg[676] = inform_R[658][5];				r_cell_reg[677] = inform_R[690][5];				r_cell_reg[678] = inform_R[659][5];				r_cell_reg[679] = inform_R[691][5];				r_cell_reg[680] = inform_R[660][5];				r_cell_reg[681] = inform_R[692][5];				r_cell_reg[682] = inform_R[661][5];				r_cell_reg[683] = inform_R[693][5];				r_cell_reg[684] = inform_R[662][5];				r_cell_reg[685] = inform_R[694][5];				r_cell_reg[686] = inform_R[663][5];				r_cell_reg[687] = inform_R[695][5];				r_cell_reg[688] = inform_R[664][5];				r_cell_reg[689] = inform_R[696][5];				r_cell_reg[690] = inform_R[665][5];				r_cell_reg[691] = inform_R[697][5];				r_cell_reg[692] = inform_R[666][5];				r_cell_reg[693] = inform_R[698][5];				r_cell_reg[694] = inform_R[667][5];				r_cell_reg[695] = inform_R[699][5];				r_cell_reg[696] = inform_R[668][5];				r_cell_reg[697] = inform_R[700][5];				r_cell_reg[698] = inform_R[669][5];				r_cell_reg[699] = inform_R[701][5];				r_cell_reg[700] = inform_R[670][5];				r_cell_reg[701] = inform_R[702][5];				r_cell_reg[702] = inform_R[671][5];				r_cell_reg[703] = inform_R[703][5];				r_cell_reg[704] = inform_R[704][5];				r_cell_reg[705] = inform_R[736][5];				r_cell_reg[706] = inform_R[705][5];				r_cell_reg[707] = inform_R[737][5];				r_cell_reg[708] = inform_R[706][5];				r_cell_reg[709] = inform_R[738][5];				r_cell_reg[710] = inform_R[707][5];				r_cell_reg[711] = inform_R[739][5];				r_cell_reg[712] = inform_R[708][5];				r_cell_reg[713] = inform_R[740][5];				r_cell_reg[714] = inform_R[709][5];				r_cell_reg[715] = inform_R[741][5];				r_cell_reg[716] = inform_R[710][5];				r_cell_reg[717] = inform_R[742][5];				r_cell_reg[718] = inform_R[711][5];				r_cell_reg[719] = inform_R[743][5];				r_cell_reg[720] = inform_R[712][5];				r_cell_reg[721] = inform_R[744][5];				r_cell_reg[722] = inform_R[713][5];				r_cell_reg[723] = inform_R[745][5];				r_cell_reg[724] = inform_R[714][5];				r_cell_reg[725] = inform_R[746][5];				r_cell_reg[726] = inform_R[715][5];				r_cell_reg[727] = inform_R[747][5];				r_cell_reg[728] = inform_R[716][5];				r_cell_reg[729] = inform_R[748][5];				r_cell_reg[730] = inform_R[717][5];				r_cell_reg[731] = inform_R[749][5];				r_cell_reg[732] = inform_R[718][5];				r_cell_reg[733] = inform_R[750][5];				r_cell_reg[734] = inform_R[719][5];				r_cell_reg[735] = inform_R[751][5];				r_cell_reg[736] = inform_R[720][5];				r_cell_reg[737] = inform_R[752][5];				r_cell_reg[738] = inform_R[721][5];				r_cell_reg[739] = inform_R[753][5];				r_cell_reg[740] = inform_R[722][5];				r_cell_reg[741] = inform_R[754][5];				r_cell_reg[742] = inform_R[723][5];				r_cell_reg[743] = inform_R[755][5];				r_cell_reg[744] = inform_R[724][5];				r_cell_reg[745] = inform_R[756][5];				r_cell_reg[746] = inform_R[725][5];				r_cell_reg[747] = inform_R[757][5];				r_cell_reg[748] = inform_R[726][5];				r_cell_reg[749] = inform_R[758][5];				r_cell_reg[750] = inform_R[727][5];				r_cell_reg[751] = inform_R[759][5];				r_cell_reg[752] = inform_R[728][5];				r_cell_reg[753] = inform_R[760][5];				r_cell_reg[754] = inform_R[729][5];				r_cell_reg[755] = inform_R[761][5];				r_cell_reg[756] = inform_R[730][5];				r_cell_reg[757] = inform_R[762][5];				r_cell_reg[758] = inform_R[731][5];				r_cell_reg[759] = inform_R[763][5];				r_cell_reg[760] = inform_R[732][5];				r_cell_reg[761] = inform_R[764][5];				r_cell_reg[762] = inform_R[733][5];				r_cell_reg[763] = inform_R[765][5];				r_cell_reg[764] = inform_R[734][5];				r_cell_reg[765] = inform_R[766][5];				r_cell_reg[766] = inform_R[735][5];				r_cell_reg[767] = inform_R[767][5];				r_cell_reg[768] = inform_R[768][5];				r_cell_reg[769] = inform_R[800][5];				r_cell_reg[770] = inform_R[769][5];				r_cell_reg[771] = inform_R[801][5];				r_cell_reg[772] = inform_R[770][5];				r_cell_reg[773] = inform_R[802][5];				r_cell_reg[774] = inform_R[771][5];				r_cell_reg[775] = inform_R[803][5];				r_cell_reg[776] = inform_R[772][5];				r_cell_reg[777] = inform_R[804][5];				r_cell_reg[778] = inform_R[773][5];				r_cell_reg[779] = inform_R[805][5];				r_cell_reg[780] = inform_R[774][5];				r_cell_reg[781] = inform_R[806][5];				r_cell_reg[782] = inform_R[775][5];				r_cell_reg[783] = inform_R[807][5];				r_cell_reg[784] = inform_R[776][5];				r_cell_reg[785] = inform_R[808][5];				r_cell_reg[786] = inform_R[777][5];				r_cell_reg[787] = inform_R[809][5];				r_cell_reg[788] = inform_R[778][5];				r_cell_reg[789] = inform_R[810][5];				r_cell_reg[790] = inform_R[779][5];				r_cell_reg[791] = inform_R[811][5];				r_cell_reg[792] = inform_R[780][5];				r_cell_reg[793] = inform_R[812][5];				r_cell_reg[794] = inform_R[781][5];				r_cell_reg[795] = inform_R[813][5];				r_cell_reg[796] = inform_R[782][5];				r_cell_reg[797] = inform_R[814][5];				r_cell_reg[798] = inform_R[783][5];				r_cell_reg[799] = inform_R[815][5];				r_cell_reg[800] = inform_R[784][5];				r_cell_reg[801] = inform_R[816][5];				r_cell_reg[802] = inform_R[785][5];				r_cell_reg[803] = inform_R[817][5];				r_cell_reg[804] = inform_R[786][5];				r_cell_reg[805] = inform_R[818][5];				r_cell_reg[806] = inform_R[787][5];				r_cell_reg[807] = inform_R[819][5];				r_cell_reg[808] = inform_R[788][5];				r_cell_reg[809] = inform_R[820][5];				r_cell_reg[810] = inform_R[789][5];				r_cell_reg[811] = inform_R[821][5];				r_cell_reg[812] = inform_R[790][5];				r_cell_reg[813] = inform_R[822][5];				r_cell_reg[814] = inform_R[791][5];				r_cell_reg[815] = inform_R[823][5];				r_cell_reg[816] = inform_R[792][5];				r_cell_reg[817] = inform_R[824][5];				r_cell_reg[818] = inform_R[793][5];				r_cell_reg[819] = inform_R[825][5];				r_cell_reg[820] = inform_R[794][5];				r_cell_reg[821] = inform_R[826][5];				r_cell_reg[822] = inform_R[795][5];				r_cell_reg[823] = inform_R[827][5];				r_cell_reg[824] = inform_R[796][5];				r_cell_reg[825] = inform_R[828][5];				r_cell_reg[826] = inform_R[797][5];				r_cell_reg[827] = inform_R[829][5];				r_cell_reg[828] = inform_R[798][5];				r_cell_reg[829] = inform_R[830][5];				r_cell_reg[830] = inform_R[799][5];				r_cell_reg[831] = inform_R[831][5];				r_cell_reg[832] = inform_R[832][5];				r_cell_reg[833] = inform_R[864][5];				r_cell_reg[834] = inform_R[833][5];				r_cell_reg[835] = inform_R[865][5];				r_cell_reg[836] = inform_R[834][5];				r_cell_reg[837] = inform_R[866][5];				r_cell_reg[838] = inform_R[835][5];				r_cell_reg[839] = inform_R[867][5];				r_cell_reg[840] = inform_R[836][5];				r_cell_reg[841] = inform_R[868][5];				r_cell_reg[842] = inform_R[837][5];				r_cell_reg[843] = inform_R[869][5];				r_cell_reg[844] = inform_R[838][5];				r_cell_reg[845] = inform_R[870][5];				r_cell_reg[846] = inform_R[839][5];				r_cell_reg[847] = inform_R[871][5];				r_cell_reg[848] = inform_R[840][5];				r_cell_reg[849] = inform_R[872][5];				r_cell_reg[850] = inform_R[841][5];				r_cell_reg[851] = inform_R[873][5];				r_cell_reg[852] = inform_R[842][5];				r_cell_reg[853] = inform_R[874][5];				r_cell_reg[854] = inform_R[843][5];				r_cell_reg[855] = inform_R[875][5];				r_cell_reg[856] = inform_R[844][5];				r_cell_reg[857] = inform_R[876][5];				r_cell_reg[858] = inform_R[845][5];				r_cell_reg[859] = inform_R[877][5];				r_cell_reg[860] = inform_R[846][5];				r_cell_reg[861] = inform_R[878][5];				r_cell_reg[862] = inform_R[847][5];				r_cell_reg[863] = inform_R[879][5];				r_cell_reg[864] = inform_R[848][5];				r_cell_reg[865] = inform_R[880][5];				r_cell_reg[866] = inform_R[849][5];				r_cell_reg[867] = inform_R[881][5];				r_cell_reg[868] = inform_R[850][5];				r_cell_reg[869] = inform_R[882][5];				r_cell_reg[870] = inform_R[851][5];				r_cell_reg[871] = inform_R[883][5];				r_cell_reg[872] = inform_R[852][5];				r_cell_reg[873] = inform_R[884][5];				r_cell_reg[874] = inform_R[853][5];				r_cell_reg[875] = inform_R[885][5];				r_cell_reg[876] = inform_R[854][5];				r_cell_reg[877] = inform_R[886][5];				r_cell_reg[878] = inform_R[855][5];				r_cell_reg[879] = inform_R[887][5];				r_cell_reg[880] = inform_R[856][5];				r_cell_reg[881] = inform_R[888][5];				r_cell_reg[882] = inform_R[857][5];				r_cell_reg[883] = inform_R[889][5];				r_cell_reg[884] = inform_R[858][5];				r_cell_reg[885] = inform_R[890][5];				r_cell_reg[886] = inform_R[859][5];				r_cell_reg[887] = inform_R[891][5];				r_cell_reg[888] = inform_R[860][5];				r_cell_reg[889] = inform_R[892][5];				r_cell_reg[890] = inform_R[861][5];				r_cell_reg[891] = inform_R[893][5];				r_cell_reg[892] = inform_R[862][5];				r_cell_reg[893] = inform_R[894][5];				r_cell_reg[894] = inform_R[863][5];				r_cell_reg[895] = inform_R[895][5];				r_cell_reg[896] = inform_R[896][5];				r_cell_reg[897] = inform_R[928][5];				r_cell_reg[898] = inform_R[897][5];				r_cell_reg[899] = inform_R[929][5];				r_cell_reg[900] = inform_R[898][5];				r_cell_reg[901] = inform_R[930][5];				r_cell_reg[902] = inform_R[899][5];				r_cell_reg[903] = inform_R[931][5];				r_cell_reg[904] = inform_R[900][5];				r_cell_reg[905] = inform_R[932][5];				r_cell_reg[906] = inform_R[901][5];				r_cell_reg[907] = inform_R[933][5];				r_cell_reg[908] = inform_R[902][5];				r_cell_reg[909] = inform_R[934][5];				r_cell_reg[910] = inform_R[903][5];				r_cell_reg[911] = inform_R[935][5];				r_cell_reg[912] = inform_R[904][5];				r_cell_reg[913] = inform_R[936][5];				r_cell_reg[914] = inform_R[905][5];				r_cell_reg[915] = inform_R[937][5];				r_cell_reg[916] = inform_R[906][5];				r_cell_reg[917] = inform_R[938][5];				r_cell_reg[918] = inform_R[907][5];				r_cell_reg[919] = inform_R[939][5];				r_cell_reg[920] = inform_R[908][5];				r_cell_reg[921] = inform_R[940][5];				r_cell_reg[922] = inform_R[909][5];				r_cell_reg[923] = inform_R[941][5];				r_cell_reg[924] = inform_R[910][5];				r_cell_reg[925] = inform_R[942][5];				r_cell_reg[926] = inform_R[911][5];				r_cell_reg[927] = inform_R[943][5];				r_cell_reg[928] = inform_R[912][5];				r_cell_reg[929] = inform_R[944][5];				r_cell_reg[930] = inform_R[913][5];				r_cell_reg[931] = inform_R[945][5];				r_cell_reg[932] = inform_R[914][5];				r_cell_reg[933] = inform_R[946][5];				r_cell_reg[934] = inform_R[915][5];				r_cell_reg[935] = inform_R[947][5];				r_cell_reg[936] = inform_R[916][5];				r_cell_reg[937] = inform_R[948][5];				r_cell_reg[938] = inform_R[917][5];				r_cell_reg[939] = inform_R[949][5];				r_cell_reg[940] = inform_R[918][5];				r_cell_reg[941] = inform_R[950][5];				r_cell_reg[942] = inform_R[919][5];				r_cell_reg[943] = inform_R[951][5];				r_cell_reg[944] = inform_R[920][5];				r_cell_reg[945] = inform_R[952][5];				r_cell_reg[946] = inform_R[921][5];				r_cell_reg[947] = inform_R[953][5];				r_cell_reg[948] = inform_R[922][5];				r_cell_reg[949] = inform_R[954][5];				r_cell_reg[950] = inform_R[923][5];				r_cell_reg[951] = inform_R[955][5];				r_cell_reg[952] = inform_R[924][5];				r_cell_reg[953] = inform_R[956][5];				r_cell_reg[954] = inform_R[925][5];				r_cell_reg[955] = inform_R[957][5];				r_cell_reg[956] = inform_R[926][5];				r_cell_reg[957] = inform_R[958][5];				r_cell_reg[958] = inform_R[927][5];				r_cell_reg[959] = inform_R[959][5];				r_cell_reg[960] = inform_R[960][5];				r_cell_reg[961] = inform_R[992][5];				r_cell_reg[962] = inform_R[961][5];				r_cell_reg[963] = inform_R[993][5];				r_cell_reg[964] = inform_R[962][5];				r_cell_reg[965] = inform_R[994][5];				r_cell_reg[966] = inform_R[963][5];				r_cell_reg[967] = inform_R[995][5];				r_cell_reg[968] = inform_R[964][5];				r_cell_reg[969] = inform_R[996][5];				r_cell_reg[970] = inform_R[965][5];				r_cell_reg[971] = inform_R[997][5];				r_cell_reg[972] = inform_R[966][5];				r_cell_reg[973] = inform_R[998][5];				r_cell_reg[974] = inform_R[967][5];				r_cell_reg[975] = inform_R[999][5];				r_cell_reg[976] = inform_R[968][5];				r_cell_reg[977] = inform_R[1000][5];				r_cell_reg[978] = inform_R[969][5];				r_cell_reg[979] = inform_R[1001][5];				r_cell_reg[980] = inform_R[970][5];				r_cell_reg[981] = inform_R[1002][5];				r_cell_reg[982] = inform_R[971][5];				r_cell_reg[983] = inform_R[1003][5];				r_cell_reg[984] = inform_R[972][5];				r_cell_reg[985] = inform_R[1004][5];				r_cell_reg[986] = inform_R[973][5];				r_cell_reg[987] = inform_R[1005][5];				r_cell_reg[988] = inform_R[974][5];				r_cell_reg[989] = inform_R[1006][5];				r_cell_reg[990] = inform_R[975][5];				r_cell_reg[991] = inform_R[1007][5];				r_cell_reg[992] = inform_R[976][5];				r_cell_reg[993] = inform_R[1008][5];				r_cell_reg[994] = inform_R[977][5];				r_cell_reg[995] = inform_R[1009][5];				r_cell_reg[996] = inform_R[978][5];				r_cell_reg[997] = inform_R[1010][5];				r_cell_reg[998] = inform_R[979][5];				r_cell_reg[999] = inform_R[1011][5];				r_cell_reg[1000] = inform_R[980][5];				r_cell_reg[1001] = inform_R[1012][5];				r_cell_reg[1002] = inform_R[981][5];				r_cell_reg[1003] = inform_R[1013][5];				r_cell_reg[1004] = inform_R[982][5];				r_cell_reg[1005] = inform_R[1014][5];				r_cell_reg[1006] = inform_R[983][5];				r_cell_reg[1007] = inform_R[1015][5];				r_cell_reg[1008] = inform_R[984][5];				r_cell_reg[1009] = inform_R[1016][5];				r_cell_reg[1010] = inform_R[985][5];				r_cell_reg[1011] = inform_R[1017][5];				r_cell_reg[1012] = inform_R[986][5];				r_cell_reg[1013] = inform_R[1018][5];				r_cell_reg[1014] = inform_R[987][5];				r_cell_reg[1015] = inform_R[1019][5];				r_cell_reg[1016] = inform_R[988][5];				r_cell_reg[1017] = inform_R[1020][5];				r_cell_reg[1018] = inform_R[989][5];				r_cell_reg[1019] = inform_R[1021][5];				r_cell_reg[1020] = inform_R[990][5];				r_cell_reg[1021] = inform_R[1022][5];				r_cell_reg[1022] = inform_R[991][5];				r_cell_reg[1023] = inform_R[1023][5];				l_cell_reg[0] = inform_L[0][6];				l_cell_reg[1] = inform_L[32][6];				l_cell_reg[2] = inform_L[1][6];				l_cell_reg[3] = inform_L[33][6];				l_cell_reg[4] = inform_L[2][6];				l_cell_reg[5] = inform_L[34][6];				l_cell_reg[6] = inform_L[3][6];				l_cell_reg[7] = inform_L[35][6];				l_cell_reg[8] = inform_L[4][6];				l_cell_reg[9] = inform_L[36][6];				l_cell_reg[10] = inform_L[5][6];				l_cell_reg[11] = inform_L[37][6];				l_cell_reg[12] = inform_L[6][6];				l_cell_reg[13] = inform_L[38][6];				l_cell_reg[14] = inform_L[7][6];				l_cell_reg[15] = inform_L[39][6];				l_cell_reg[16] = inform_L[8][6];				l_cell_reg[17] = inform_L[40][6];				l_cell_reg[18] = inform_L[9][6];				l_cell_reg[19] = inform_L[41][6];				l_cell_reg[20] = inform_L[10][6];				l_cell_reg[21] = inform_L[42][6];				l_cell_reg[22] = inform_L[11][6];				l_cell_reg[23] = inform_L[43][6];				l_cell_reg[24] = inform_L[12][6];				l_cell_reg[25] = inform_L[44][6];				l_cell_reg[26] = inform_L[13][6];				l_cell_reg[27] = inform_L[45][6];				l_cell_reg[28] = inform_L[14][6];				l_cell_reg[29] = inform_L[46][6];				l_cell_reg[30] = inform_L[15][6];				l_cell_reg[31] = inform_L[47][6];				l_cell_reg[32] = inform_L[16][6];				l_cell_reg[33] = inform_L[48][6];				l_cell_reg[34] = inform_L[17][6];				l_cell_reg[35] = inform_L[49][6];				l_cell_reg[36] = inform_L[18][6];				l_cell_reg[37] = inform_L[50][6];				l_cell_reg[38] = inform_L[19][6];				l_cell_reg[39] = inform_L[51][6];				l_cell_reg[40] = inform_L[20][6];				l_cell_reg[41] = inform_L[52][6];				l_cell_reg[42] = inform_L[21][6];				l_cell_reg[43] = inform_L[53][6];				l_cell_reg[44] = inform_L[22][6];				l_cell_reg[45] = inform_L[54][6];				l_cell_reg[46] = inform_L[23][6];				l_cell_reg[47] = inform_L[55][6];				l_cell_reg[48] = inform_L[24][6];				l_cell_reg[49] = inform_L[56][6];				l_cell_reg[50] = inform_L[25][6];				l_cell_reg[51] = inform_L[57][6];				l_cell_reg[52] = inform_L[26][6];				l_cell_reg[53] = inform_L[58][6];				l_cell_reg[54] = inform_L[27][6];				l_cell_reg[55] = inform_L[59][6];				l_cell_reg[56] = inform_L[28][6];				l_cell_reg[57] = inform_L[60][6];				l_cell_reg[58] = inform_L[29][6];				l_cell_reg[59] = inform_L[61][6];				l_cell_reg[60] = inform_L[30][6];				l_cell_reg[61] = inform_L[62][6];				l_cell_reg[62] = inform_L[31][6];				l_cell_reg[63] = inform_L[63][6];				l_cell_reg[64] = inform_L[64][6];				l_cell_reg[65] = inform_L[96][6];				l_cell_reg[66] = inform_L[65][6];				l_cell_reg[67] = inform_L[97][6];				l_cell_reg[68] = inform_L[66][6];				l_cell_reg[69] = inform_L[98][6];				l_cell_reg[70] = inform_L[67][6];				l_cell_reg[71] = inform_L[99][6];				l_cell_reg[72] = inform_L[68][6];				l_cell_reg[73] = inform_L[100][6];				l_cell_reg[74] = inform_L[69][6];				l_cell_reg[75] = inform_L[101][6];				l_cell_reg[76] = inform_L[70][6];				l_cell_reg[77] = inform_L[102][6];				l_cell_reg[78] = inform_L[71][6];				l_cell_reg[79] = inform_L[103][6];				l_cell_reg[80] = inform_L[72][6];				l_cell_reg[81] = inform_L[104][6];				l_cell_reg[82] = inform_L[73][6];				l_cell_reg[83] = inform_L[105][6];				l_cell_reg[84] = inform_L[74][6];				l_cell_reg[85] = inform_L[106][6];				l_cell_reg[86] = inform_L[75][6];				l_cell_reg[87] = inform_L[107][6];				l_cell_reg[88] = inform_L[76][6];				l_cell_reg[89] = inform_L[108][6];				l_cell_reg[90] = inform_L[77][6];				l_cell_reg[91] = inform_L[109][6];				l_cell_reg[92] = inform_L[78][6];				l_cell_reg[93] = inform_L[110][6];				l_cell_reg[94] = inform_L[79][6];				l_cell_reg[95] = inform_L[111][6];				l_cell_reg[96] = inform_L[80][6];				l_cell_reg[97] = inform_L[112][6];				l_cell_reg[98] = inform_L[81][6];				l_cell_reg[99] = inform_L[113][6];				l_cell_reg[100] = inform_L[82][6];				l_cell_reg[101] = inform_L[114][6];				l_cell_reg[102] = inform_L[83][6];				l_cell_reg[103] = inform_L[115][6];				l_cell_reg[104] = inform_L[84][6];				l_cell_reg[105] = inform_L[116][6];				l_cell_reg[106] = inform_L[85][6];				l_cell_reg[107] = inform_L[117][6];				l_cell_reg[108] = inform_L[86][6];				l_cell_reg[109] = inform_L[118][6];				l_cell_reg[110] = inform_L[87][6];				l_cell_reg[111] = inform_L[119][6];				l_cell_reg[112] = inform_L[88][6];				l_cell_reg[113] = inform_L[120][6];				l_cell_reg[114] = inform_L[89][6];				l_cell_reg[115] = inform_L[121][6];				l_cell_reg[116] = inform_L[90][6];				l_cell_reg[117] = inform_L[122][6];				l_cell_reg[118] = inform_L[91][6];				l_cell_reg[119] = inform_L[123][6];				l_cell_reg[120] = inform_L[92][6];				l_cell_reg[121] = inform_L[124][6];				l_cell_reg[122] = inform_L[93][6];				l_cell_reg[123] = inform_L[125][6];				l_cell_reg[124] = inform_L[94][6];				l_cell_reg[125] = inform_L[126][6];				l_cell_reg[126] = inform_L[95][6];				l_cell_reg[127] = inform_L[127][6];				l_cell_reg[128] = inform_L[128][6];				l_cell_reg[129] = inform_L[160][6];				l_cell_reg[130] = inform_L[129][6];				l_cell_reg[131] = inform_L[161][6];				l_cell_reg[132] = inform_L[130][6];				l_cell_reg[133] = inform_L[162][6];				l_cell_reg[134] = inform_L[131][6];				l_cell_reg[135] = inform_L[163][6];				l_cell_reg[136] = inform_L[132][6];				l_cell_reg[137] = inform_L[164][6];				l_cell_reg[138] = inform_L[133][6];				l_cell_reg[139] = inform_L[165][6];				l_cell_reg[140] = inform_L[134][6];				l_cell_reg[141] = inform_L[166][6];				l_cell_reg[142] = inform_L[135][6];				l_cell_reg[143] = inform_L[167][6];				l_cell_reg[144] = inform_L[136][6];				l_cell_reg[145] = inform_L[168][6];				l_cell_reg[146] = inform_L[137][6];				l_cell_reg[147] = inform_L[169][6];				l_cell_reg[148] = inform_L[138][6];				l_cell_reg[149] = inform_L[170][6];				l_cell_reg[150] = inform_L[139][6];				l_cell_reg[151] = inform_L[171][6];				l_cell_reg[152] = inform_L[140][6];				l_cell_reg[153] = inform_L[172][6];				l_cell_reg[154] = inform_L[141][6];				l_cell_reg[155] = inform_L[173][6];				l_cell_reg[156] = inform_L[142][6];				l_cell_reg[157] = inform_L[174][6];				l_cell_reg[158] = inform_L[143][6];				l_cell_reg[159] = inform_L[175][6];				l_cell_reg[160] = inform_L[144][6];				l_cell_reg[161] = inform_L[176][6];				l_cell_reg[162] = inform_L[145][6];				l_cell_reg[163] = inform_L[177][6];				l_cell_reg[164] = inform_L[146][6];				l_cell_reg[165] = inform_L[178][6];				l_cell_reg[166] = inform_L[147][6];				l_cell_reg[167] = inform_L[179][6];				l_cell_reg[168] = inform_L[148][6];				l_cell_reg[169] = inform_L[180][6];				l_cell_reg[170] = inform_L[149][6];				l_cell_reg[171] = inform_L[181][6];				l_cell_reg[172] = inform_L[150][6];				l_cell_reg[173] = inform_L[182][6];				l_cell_reg[174] = inform_L[151][6];				l_cell_reg[175] = inform_L[183][6];				l_cell_reg[176] = inform_L[152][6];				l_cell_reg[177] = inform_L[184][6];				l_cell_reg[178] = inform_L[153][6];				l_cell_reg[179] = inform_L[185][6];				l_cell_reg[180] = inform_L[154][6];				l_cell_reg[181] = inform_L[186][6];				l_cell_reg[182] = inform_L[155][6];				l_cell_reg[183] = inform_L[187][6];				l_cell_reg[184] = inform_L[156][6];				l_cell_reg[185] = inform_L[188][6];				l_cell_reg[186] = inform_L[157][6];				l_cell_reg[187] = inform_L[189][6];				l_cell_reg[188] = inform_L[158][6];				l_cell_reg[189] = inform_L[190][6];				l_cell_reg[190] = inform_L[159][6];				l_cell_reg[191] = inform_L[191][6];				l_cell_reg[192] = inform_L[192][6];				l_cell_reg[193] = inform_L[224][6];				l_cell_reg[194] = inform_L[193][6];				l_cell_reg[195] = inform_L[225][6];				l_cell_reg[196] = inform_L[194][6];				l_cell_reg[197] = inform_L[226][6];				l_cell_reg[198] = inform_L[195][6];				l_cell_reg[199] = inform_L[227][6];				l_cell_reg[200] = inform_L[196][6];				l_cell_reg[201] = inform_L[228][6];				l_cell_reg[202] = inform_L[197][6];				l_cell_reg[203] = inform_L[229][6];				l_cell_reg[204] = inform_L[198][6];				l_cell_reg[205] = inform_L[230][6];				l_cell_reg[206] = inform_L[199][6];				l_cell_reg[207] = inform_L[231][6];				l_cell_reg[208] = inform_L[200][6];				l_cell_reg[209] = inform_L[232][6];				l_cell_reg[210] = inform_L[201][6];				l_cell_reg[211] = inform_L[233][6];				l_cell_reg[212] = inform_L[202][6];				l_cell_reg[213] = inform_L[234][6];				l_cell_reg[214] = inform_L[203][6];				l_cell_reg[215] = inform_L[235][6];				l_cell_reg[216] = inform_L[204][6];				l_cell_reg[217] = inform_L[236][6];				l_cell_reg[218] = inform_L[205][6];				l_cell_reg[219] = inform_L[237][6];				l_cell_reg[220] = inform_L[206][6];				l_cell_reg[221] = inform_L[238][6];				l_cell_reg[222] = inform_L[207][6];				l_cell_reg[223] = inform_L[239][6];				l_cell_reg[224] = inform_L[208][6];				l_cell_reg[225] = inform_L[240][6];				l_cell_reg[226] = inform_L[209][6];				l_cell_reg[227] = inform_L[241][6];				l_cell_reg[228] = inform_L[210][6];				l_cell_reg[229] = inform_L[242][6];				l_cell_reg[230] = inform_L[211][6];				l_cell_reg[231] = inform_L[243][6];				l_cell_reg[232] = inform_L[212][6];				l_cell_reg[233] = inform_L[244][6];				l_cell_reg[234] = inform_L[213][6];				l_cell_reg[235] = inform_L[245][6];				l_cell_reg[236] = inform_L[214][6];				l_cell_reg[237] = inform_L[246][6];				l_cell_reg[238] = inform_L[215][6];				l_cell_reg[239] = inform_L[247][6];				l_cell_reg[240] = inform_L[216][6];				l_cell_reg[241] = inform_L[248][6];				l_cell_reg[242] = inform_L[217][6];				l_cell_reg[243] = inform_L[249][6];				l_cell_reg[244] = inform_L[218][6];				l_cell_reg[245] = inform_L[250][6];				l_cell_reg[246] = inform_L[219][6];				l_cell_reg[247] = inform_L[251][6];				l_cell_reg[248] = inform_L[220][6];				l_cell_reg[249] = inform_L[252][6];				l_cell_reg[250] = inform_L[221][6];				l_cell_reg[251] = inform_L[253][6];				l_cell_reg[252] = inform_L[222][6];				l_cell_reg[253] = inform_L[254][6];				l_cell_reg[254] = inform_L[223][6];				l_cell_reg[255] = inform_L[255][6];				l_cell_reg[256] = inform_L[256][6];				l_cell_reg[257] = inform_L[288][6];				l_cell_reg[258] = inform_L[257][6];				l_cell_reg[259] = inform_L[289][6];				l_cell_reg[260] = inform_L[258][6];				l_cell_reg[261] = inform_L[290][6];				l_cell_reg[262] = inform_L[259][6];				l_cell_reg[263] = inform_L[291][6];				l_cell_reg[264] = inform_L[260][6];				l_cell_reg[265] = inform_L[292][6];				l_cell_reg[266] = inform_L[261][6];				l_cell_reg[267] = inform_L[293][6];				l_cell_reg[268] = inform_L[262][6];				l_cell_reg[269] = inform_L[294][6];				l_cell_reg[270] = inform_L[263][6];				l_cell_reg[271] = inform_L[295][6];				l_cell_reg[272] = inform_L[264][6];				l_cell_reg[273] = inform_L[296][6];				l_cell_reg[274] = inform_L[265][6];				l_cell_reg[275] = inform_L[297][6];				l_cell_reg[276] = inform_L[266][6];				l_cell_reg[277] = inform_L[298][6];				l_cell_reg[278] = inform_L[267][6];				l_cell_reg[279] = inform_L[299][6];				l_cell_reg[280] = inform_L[268][6];				l_cell_reg[281] = inform_L[300][6];				l_cell_reg[282] = inform_L[269][6];				l_cell_reg[283] = inform_L[301][6];				l_cell_reg[284] = inform_L[270][6];				l_cell_reg[285] = inform_L[302][6];				l_cell_reg[286] = inform_L[271][6];				l_cell_reg[287] = inform_L[303][6];				l_cell_reg[288] = inform_L[272][6];				l_cell_reg[289] = inform_L[304][6];				l_cell_reg[290] = inform_L[273][6];				l_cell_reg[291] = inform_L[305][6];				l_cell_reg[292] = inform_L[274][6];				l_cell_reg[293] = inform_L[306][6];				l_cell_reg[294] = inform_L[275][6];				l_cell_reg[295] = inform_L[307][6];				l_cell_reg[296] = inform_L[276][6];				l_cell_reg[297] = inform_L[308][6];				l_cell_reg[298] = inform_L[277][6];				l_cell_reg[299] = inform_L[309][6];				l_cell_reg[300] = inform_L[278][6];				l_cell_reg[301] = inform_L[310][6];				l_cell_reg[302] = inform_L[279][6];				l_cell_reg[303] = inform_L[311][6];				l_cell_reg[304] = inform_L[280][6];				l_cell_reg[305] = inform_L[312][6];				l_cell_reg[306] = inform_L[281][6];				l_cell_reg[307] = inform_L[313][6];				l_cell_reg[308] = inform_L[282][6];				l_cell_reg[309] = inform_L[314][6];				l_cell_reg[310] = inform_L[283][6];				l_cell_reg[311] = inform_L[315][6];				l_cell_reg[312] = inform_L[284][6];				l_cell_reg[313] = inform_L[316][6];				l_cell_reg[314] = inform_L[285][6];				l_cell_reg[315] = inform_L[317][6];				l_cell_reg[316] = inform_L[286][6];				l_cell_reg[317] = inform_L[318][6];				l_cell_reg[318] = inform_L[287][6];				l_cell_reg[319] = inform_L[319][6];				l_cell_reg[320] = inform_L[320][6];				l_cell_reg[321] = inform_L[352][6];				l_cell_reg[322] = inform_L[321][6];				l_cell_reg[323] = inform_L[353][6];				l_cell_reg[324] = inform_L[322][6];				l_cell_reg[325] = inform_L[354][6];				l_cell_reg[326] = inform_L[323][6];				l_cell_reg[327] = inform_L[355][6];				l_cell_reg[328] = inform_L[324][6];				l_cell_reg[329] = inform_L[356][6];				l_cell_reg[330] = inform_L[325][6];				l_cell_reg[331] = inform_L[357][6];				l_cell_reg[332] = inform_L[326][6];				l_cell_reg[333] = inform_L[358][6];				l_cell_reg[334] = inform_L[327][6];				l_cell_reg[335] = inform_L[359][6];				l_cell_reg[336] = inform_L[328][6];				l_cell_reg[337] = inform_L[360][6];				l_cell_reg[338] = inform_L[329][6];				l_cell_reg[339] = inform_L[361][6];				l_cell_reg[340] = inform_L[330][6];				l_cell_reg[341] = inform_L[362][6];				l_cell_reg[342] = inform_L[331][6];				l_cell_reg[343] = inform_L[363][6];				l_cell_reg[344] = inform_L[332][6];				l_cell_reg[345] = inform_L[364][6];				l_cell_reg[346] = inform_L[333][6];				l_cell_reg[347] = inform_L[365][6];				l_cell_reg[348] = inform_L[334][6];				l_cell_reg[349] = inform_L[366][6];				l_cell_reg[350] = inform_L[335][6];				l_cell_reg[351] = inform_L[367][6];				l_cell_reg[352] = inform_L[336][6];				l_cell_reg[353] = inform_L[368][6];				l_cell_reg[354] = inform_L[337][6];				l_cell_reg[355] = inform_L[369][6];				l_cell_reg[356] = inform_L[338][6];				l_cell_reg[357] = inform_L[370][6];				l_cell_reg[358] = inform_L[339][6];				l_cell_reg[359] = inform_L[371][6];				l_cell_reg[360] = inform_L[340][6];				l_cell_reg[361] = inform_L[372][6];				l_cell_reg[362] = inform_L[341][6];				l_cell_reg[363] = inform_L[373][6];				l_cell_reg[364] = inform_L[342][6];				l_cell_reg[365] = inform_L[374][6];				l_cell_reg[366] = inform_L[343][6];				l_cell_reg[367] = inform_L[375][6];				l_cell_reg[368] = inform_L[344][6];				l_cell_reg[369] = inform_L[376][6];				l_cell_reg[370] = inform_L[345][6];				l_cell_reg[371] = inform_L[377][6];				l_cell_reg[372] = inform_L[346][6];				l_cell_reg[373] = inform_L[378][6];				l_cell_reg[374] = inform_L[347][6];				l_cell_reg[375] = inform_L[379][6];				l_cell_reg[376] = inform_L[348][6];				l_cell_reg[377] = inform_L[380][6];				l_cell_reg[378] = inform_L[349][6];				l_cell_reg[379] = inform_L[381][6];				l_cell_reg[380] = inform_L[350][6];				l_cell_reg[381] = inform_L[382][6];				l_cell_reg[382] = inform_L[351][6];				l_cell_reg[383] = inform_L[383][6];				l_cell_reg[384] = inform_L[384][6];				l_cell_reg[385] = inform_L[416][6];				l_cell_reg[386] = inform_L[385][6];				l_cell_reg[387] = inform_L[417][6];				l_cell_reg[388] = inform_L[386][6];				l_cell_reg[389] = inform_L[418][6];				l_cell_reg[390] = inform_L[387][6];				l_cell_reg[391] = inform_L[419][6];				l_cell_reg[392] = inform_L[388][6];				l_cell_reg[393] = inform_L[420][6];				l_cell_reg[394] = inform_L[389][6];				l_cell_reg[395] = inform_L[421][6];				l_cell_reg[396] = inform_L[390][6];				l_cell_reg[397] = inform_L[422][6];				l_cell_reg[398] = inform_L[391][6];				l_cell_reg[399] = inform_L[423][6];				l_cell_reg[400] = inform_L[392][6];				l_cell_reg[401] = inform_L[424][6];				l_cell_reg[402] = inform_L[393][6];				l_cell_reg[403] = inform_L[425][6];				l_cell_reg[404] = inform_L[394][6];				l_cell_reg[405] = inform_L[426][6];				l_cell_reg[406] = inform_L[395][6];				l_cell_reg[407] = inform_L[427][6];				l_cell_reg[408] = inform_L[396][6];				l_cell_reg[409] = inform_L[428][6];				l_cell_reg[410] = inform_L[397][6];				l_cell_reg[411] = inform_L[429][6];				l_cell_reg[412] = inform_L[398][6];				l_cell_reg[413] = inform_L[430][6];				l_cell_reg[414] = inform_L[399][6];				l_cell_reg[415] = inform_L[431][6];				l_cell_reg[416] = inform_L[400][6];				l_cell_reg[417] = inform_L[432][6];				l_cell_reg[418] = inform_L[401][6];				l_cell_reg[419] = inform_L[433][6];				l_cell_reg[420] = inform_L[402][6];				l_cell_reg[421] = inform_L[434][6];				l_cell_reg[422] = inform_L[403][6];				l_cell_reg[423] = inform_L[435][6];				l_cell_reg[424] = inform_L[404][6];				l_cell_reg[425] = inform_L[436][6];				l_cell_reg[426] = inform_L[405][6];				l_cell_reg[427] = inform_L[437][6];				l_cell_reg[428] = inform_L[406][6];				l_cell_reg[429] = inform_L[438][6];				l_cell_reg[430] = inform_L[407][6];				l_cell_reg[431] = inform_L[439][6];				l_cell_reg[432] = inform_L[408][6];				l_cell_reg[433] = inform_L[440][6];				l_cell_reg[434] = inform_L[409][6];				l_cell_reg[435] = inform_L[441][6];				l_cell_reg[436] = inform_L[410][6];				l_cell_reg[437] = inform_L[442][6];				l_cell_reg[438] = inform_L[411][6];				l_cell_reg[439] = inform_L[443][6];				l_cell_reg[440] = inform_L[412][6];				l_cell_reg[441] = inform_L[444][6];				l_cell_reg[442] = inform_L[413][6];				l_cell_reg[443] = inform_L[445][6];				l_cell_reg[444] = inform_L[414][6];				l_cell_reg[445] = inform_L[446][6];				l_cell_reg[446] = inform_L[415][6];				l_cell_reg[447] = inform_L[447][6];				l_cell_reg[448] = inform_L[448][6];				l_cell_reg[449] = inform_L[480][6];				l_cell_reg[450] = inform_L[449][6];				l_cell_reg[451] = inform_L[481][6];				l_cell_reg[452] = inform_L[450][6];				l_cell_reg[453] = inform_L[482][6];				l_cell_reg[454] = inform_L[451][6];				l_cell_reg[455] = inform_L[483][6];				l_cell_reg[456] = inform_L[452][6];				l_cell_reg[457] = inform_L[484][6];				l_cell_reg[458] = inform_L[453][6];				l_cell_reg[459] = inform_L[485][6];				l_cell_reg[460] = inform_L[454][6];				l_cell_reg[461] = inform_L[486][6];				l_cell_reg[462] = inform_L[455][6];				l_cell_reg[463] = inform_L[487][6];				l_cell_reg[464] = inform_L[456][6];				l_cell_reg[465] = inform_L[488][6];				l_cell_reg[466] = inform_L[457][6];				l_cell_reg[467] = inform_L[489][6];				l_cell_reg[468] = inform_L[458][6];				l_cell_reg[469] = inform_L[490][6];				l_cell_reg[470] = inform_L[459][6];				l_cell_reg[471] = inform_L[491][6];				l_cell_reg[472] = inform_L[460][6];				l_cell_reg[473] = inform_L[492][6];				l_cell_reg[474] = inform_L[461][6];				l_cell_reg[475] = inform_L[493][6];				l_cell_reg[476] = inform_L[462][6];				l_cell_reg[477] = inform_L[494][6];				l_cell_reg[478] = inform_L[463][6];				l_cell_reg[479] = inform_L[495][6];				l_cell_reg[480] = inform_L[464][6];				l_cell_reg[481] = inform_L[496][6];				l_cell_reg[482] = inform_L[465][6];				l_cell_reg[483] = inform_L[497][6];				l_cell_reg[484] = inform_L[466][6];				l_cell_reg[485] = inform_L[498][6];				l_cell_reg[486] = inform_L[467][6];				l_cell_reg[487] = inform_L[499][6];				l_cell_reg[488] = inform_L[468][6];				l_cell_reg[489] = inform_L[500][6];				l_cell_reg[490] = inform_L[469][6];				l_cell_reg[491] = inform_L[501][6];				l_cell_reg[492] = inform_L[470][6];				l_cell_reg[493] = inform_L[502][6];				l_cell_reg[494] = inform_L[471][6];				l_cell_reg[495] = inform_L[503][6];				l_cell_reg[496] = inform_L[472][6];				l_cell_reg[497] = inform_L[504][6];				l_cell_reg[498] = inform_L[473][6];				l_cell_reg[499] = inform_L[505][6];				l_cell_reg[500] = inform_L[474][6];				l_cell_reg[501] = inform_L[506][6];				l_cell_reg[502] = inform_L[475][6];				l_cell_reg[503] = inform_L[507][6];				l_cell_reg[504] = inform_L[476][6];				l_cell_reg[505] = inform_L[508][6];				l_cell_reg[506] = inform_L[477][6];				l_cell_reg[507] = inform_L[509][6];				l_cell_reg[508] = inform_L[478][6];				l_cell_reg[509] = inform_L[510][6];				l_cell_reg[510] = inform_L[479][6];				l_cell_reg[511] = inform_L[511][6];				l_cell_reg[512] = inform_L[512][6];				l_cell_reg[513] = inform_L[544][6];				l_cell_reg[514] = inform_L[513][6];				l_cell_reg[515] = inform_L[545][6];				l_cell_reg[516] = inform_L[514][6];				l_cell_reg[517] = inform_L[546][6];				l_cell_reg[518] = inform_L[515][6];				l_cell_reg[519] = inform_L[547][6];				l_cell_reg[520] = inform_L[516][6];				l_cell_reg[521] = inform_L[548][6];				l_cell_reg[522] = inform_L[517][6];				l_cell_reg[523] = inform_L[549][6];				l_cell_reg[524] = inform_L[518][6];				l_cell_reg[525] = inform_L[550][6];				l_cell_reg[526] = inform_L[519][6];				l_cell_reg[527] = inform_L[551][6];				l_cell_reg[528] = inform_L[520][6];				l_cell_reg[529] = inform_L[552][6];				l_cell_reg[530] = inform_L[521][6];				l_cell_reg[531] = inform_L[553][6];				l_cell_reg[532] = inform_L[522][6];				l_cell_reg[533] = inform_L[554][6];				l_cell_reg[534] = inform_L[523][6];				l_cell_reg[535] = inform_L[555][6];				l_cell_reg[536] = inform_L[524][6];				l_cell_reg[537] = inform_L[556][6];				l_cell_reg[538] = inform_L[525][6];				l_cell_reg[539] = inform_L[557][6];				l_cell_reg[540] = inform_L[526][6];				l_cell_reg[541] = inform_L[558][6];				l_cell_reg[542] = inform_L[527][6];				l_cell_reg[543] = inform_L[559][6];				l_cell_reg[544] = inform_L[528][6];				l_cell_reg[545] = inform_L[560][6];				l_cell_reg[546] = inform_L[529][6];				l_cell_reg[547] = inform_L[561][6];				l_cell_reg[548] = inform_L[530][6];				l_cell_reg[549] = inform_L[562][6];				l_cell_reg[550] = inform_L[531][6];				l_cell_reg[551] = inform_L[563][6];				l_cell_reg[552] = inform_L[532][6];				l_cell_reg[553] = inform_L[564][6];				l_cell_reg[554] = inform_L[533][6];				l_cell_reg[555] = inform_L[565][6];				l_cell_reg[556] = inform_L[534][6];				l_cell_reg[557] = inform_L[566][6];				l_cell_reg[558] = inform_L[535][6];				l_cell_reg[559] = inform_L[567][6];				l_cell_reg[560] = inform_L[536][6];				l_cell_reg[561] = inform_L[568][6];				l_cell_reg[562] = inform_L[537][6];				l_cell_reg[563] = inform_L[569][6];				l_cell_reg[564] = inform_L[538][6];				l_cell_reg[565] = inform_L[570][6];				l_cell_reg[566] = inform_L[539][6];				l_cell_reg[567] = inform_L[571][6];				l_cell_reg[568] = inform_L[540][6];				l_cell_reg[569] = inform_L[572][6];				l_cell_reg[570] = inform_L[541][6];				l_cell_reg[571] = inform_L[573][6];				l_cell_reg[572] = inform_L[542][6];				l_cell_reg[573] = inform_L[574][6];				l_cell_reg[574] = inform_L[543][6];				l_cell_reg[575] = inform_L[575][6];				l_cell_reg[576] = inform_L[576][6];				l_cell_reg[577] = inform_L[608][6];				l_cell_reg[578] = inform_L[577][6];				l_cell_reg[579] = inform_L[609][6];				l_cell_reg[580] = inform_L[578][6];				l_cell_reg[581] = inform_L[610][6];				l_cell_reg[582] = inform_L[579][6];				l_cell_reg[583] = inform_L[611][6];				l_cell_reg[584] = inform_L[580][6];				l_cell_reg[585] = inform_L[612][6];				l_cell_reg[586] = inform_L[581][6];				l_cell_reg[587] = inform_L[613][6];				l_cell_reg[588] = inform_L[582][6];				l_cell_reg[589] = inform_L[614][6];				l_cell_reg[590] = inform_L[583][6];				l_cell_reg[591] = inform_L[615][6];				l_cell_reg[592] = inform_L[584][6];				l_cell_reg[593] = inform_L[616][6];				l_cell_reg[594] = inform_L[585][6];				l_cell_reg[595] = inform_L[617][6];				l_cell_reg[596] = inform_L[586][6];				l_cell_reg[597] = inform_L[618][6];				l_cell_reg[598] = inform_L[587][6];				l_cell_reg[599] = inform_L[619][6];				l_cell_reg[600] = inform_L[588][6];				l_cell_reg[601] = inform_L[620][6];				l_cell_reg[602] = inform_L[589][6];				l_cell_reg[603] = inform_L[621][6];				l_cell_reg[604] = inform_L[590][6];				l_cell_reg[605] = inform_L[622][6];				l_cell_reg[606] = inform_L[591][6];				l_cell_reg[607] = inform_L[623][6];				l_cell_reg[608] = inform_L[592][6];				l_cell_reg[609] = inform_L[624][6];				l_cell_reg[610] = inform_L[593][6];				l_cell_reg[611] = inform_L[625][6];				l_cell_reg[612] = inform_L[594][6];				l_cell_reg[613] = inform_L[626][6];				l_cell_reg[614] = inform_L[595][6];				l_cell_reg[615] = inform_L[627][6];				l_cell_reg[616] = inform_L[596][6];				l_cell_reg[617] = inform_L[628][6];				l_cell_reg[618] = inform_L[597][6];				l_cell_reg[619] = inform_L[629][6];				l_cell_reg[620] = inform_L[598][6];				l_cell_reg[621] = inform_L[630][6];				l_cell_reg[622] = inform_L[599][6];				l_cell_reg[623] = inform_L[631][6];				l_cell_reg[624] = inform_L[600][6];				l_cell_reg[625] = inform_L[632][6];				l_cell_reg[626] = inform_L[601][6];				l_cell_reg[627] = inform_L[633][6];				l_cell_reg[628] = inform_L[602][6];				l_cell_reg[629] = inform_L[634][6];				l_cell_reg[630] = inform_L[603][6];				l_cell_reg[631] = inform_L[635][6];				l_cell_reg[632] = inform_L[604][6];				l_cell_reg[633] = inform_L[636][6];				l_cell_reg[634] = inform_L[605][6];				l_cell_reg[635] = inform_L[637][6];				l_cell_reg[636] = inform_L[606][6];				l_cell_reg[637] = inform_L[638][6];				l_cell_reg[638] = inform_L[607][6];				l_cell_reg[639] = inform_L[639][6];				l_cell_reg[640] = inform_L[640][6];				l_cell_reg[641] = inform_L[672][6];				l_cell_reg[642] = inform_L[641][6];				l_cell_reg[643] = inform_L[673][6];				l_cell_reg[644] = inform_L[642][6];				l_cell_reg[645] = inform_L[674][6];				l_cell_reg[646] = inform_L[643][6];				l_cell_reg[647] = inform_L[675][6];				l_cell_reg[648] = inform_L[644][6];				l_cell_reg[649] = inform_L[676][6];				l_cell_reg[650] = inform_L[645][6];				l_cell_reg[651] = inform_L[677][6];				l_cell_reg[652] = inform_L[646][6];				l_cell_reg[653] = inform_L[678][6];				l_cell_reg[654] = inform_L[647][6];				l_cell_reg[655] = inform_L[679][6];				l_cell_reg[656] = inform_L[648][6];				l_cell_reg[657] = inform_L[680][6];				l_cell_reg[658] = inform_L[649][6];				l_cell_reg[659] = inform_L[681][6];				l_cell_reg[660] = inform_L[650][6];				l_cell_reg[661] = inform_L[682][6];				l_cell_reg[662] = inform_L[651][6];				l_cell_reg[663] = inform_L[683][6];				l_cell_reg[664] = inform_L[652][6];				l_cell_reg[665] = inform_L[684][6];				l_cell_reg[666] = inform_L[653][6];				l_cell_reg[667] = inform_L[685][6];				l_cell_reg[668] = inform_L[654][6];				l_cell_reg[669] = inform_L[686][6];				l_cell_reg[670] = inform_L[655][6];				l_cell_reg[671] = inform_L[687][6];				l_cell_reg[672] = inform_L[656][6];				l_cell_reg[673] = inform_L[688][6];				l_cell_reg[674] = inform_L[657][6];				l_cell_reg[675] = inform_L[689][6];				l_cell_reg[676] = inform_L[658][6];				l_cell_reg[677] = inform_L[690][6];				l_cell_reg[678] = inform_L[659][6];				l_cell_reg[679] = inform_L[691][6];				l_cell_reg[680] = inform_L[660][6];				l_cell_reg[681] = inform_L[692][6];				l_cell_reg[682] = inform_L[661][6];				l_cell_reg[683] = inform_L[693][6];				l_cell_reg[684] = inform_L[662][6];				l_cell_reg[685] = inform_L[694][6];				l_cell_reg[686] = inform_L[663][6];				l_cell_reg[687] = inform_L[695][6];				l_cell_reg[688] = inform_L[664][6];				l_cell_reg[689] = inform_L[696][6];				l_cell_reg[690] = inform_L[665][6];				l_cell_reg[691] = inform_L[697][6];				l_cell_reg[692] = inform_L[666][6];				l_cell_reg[693] = inform_L[698][6];				l_cell_reg[694] = inform_L[667][6];				l_cell_reg[695] = inform_L[699][6];				l_cell_reg[696] = inform_L[668][6];				l_cell_reg[697] = inform_L[700][6];				l_cell_reg[698] = inform_L[669][6];				l_cell_reg[699] = inform_L[701][6];				l_cell_reg[700] = inform_L[670][6];				l_cell_reg[701] = inform_L[702][6];				l_cell_reg[702] = inform_L[671][6];				l_cell_reg[703] = inform_L[703][6];				l_cell_reg[704] = inform_L[704][6];				l_cell_reg[705] = inform_L[736][6];				l_cell_reg[706] = inform_L[705][6];				l_cell_reg[707] = inform_L[737][6];				l_cell_reg[708] = inform_L[706][6];				l_cell_reg[709] = inform_L[738][6];				l_cell_reg[710] = inform_L[707][6];				l_cell_reg[711] = inform_L[739][6];				l_cell_reg[712] = inform_L[708][6];				l_cell_reg[713] = inform_L[740][6];				l_cell_reg[714] = inform_L[709][6];				l_cell_reg[715] = inform_L[741][6];				l_cell_reg[716] = inform_L[710][6];				l_cell_reg[717] = inform_L[742][6];				l_cell_reg[718] = inform_L[711][6];				l_cell_reg[719] = inform_L[743][6];				l_cell_reg[720] = inform_L[712][6];				l_cell_reg[721] = inform_L[744][6];				l_cell_reg[722] = inform_L[713][6];				l_cell_reg[723] = inform_L[745][6];				l_cell_reg[724] = inform_L[714][6];				l_cell_reg[725] = inform_L[746][6];				l_cell_reg[726] = inform_L[715][6];				l_cell_reg[727] = inform_L[747][6];				l_cell_reg[728] = inform_L[716][6];				l_cell_reg[729] = inform_L[748][6];				l_cell_reg[730] = inform_L[717][6];				l_cell_reg[731] = inform_L[749][6];				l_cell_reg[732] = inform_L[718][6];				l_cell_reg[733] = inform_L[750][6];				l_cell_reg[734] = inform_L[719][6];				l_cell_reg[735] = inform_L[751][6];				l_cell_reg[736] = inform_L[720][6];				l_cell_reg[737] = inform_L[752][6];				l_cell_reg[738] = inform_L[721][6];				l_cell_reg[739] = inform_L[753][6];				l_cell_reg[740] = inform_L[722][6];				l_cell_reg[741] = inform_L[754][6];				l_cell_reg[742] = inform_L[723][6];				l_cell_reg[743] = inform_L[755][6];				l_cell_reg[744] = inform_L[724][6];				l_cell_reg[745] = inform_L[756][6];				l_cell_reg[746] = inform_L[725][6];				l_cell_reg[747] = inform_L[757][6];				l_cell_reg[748] = inform_L[726][6];				l_cell_reg[749] = inform_L[758][6];				l_cell_reg[750] = inform_L[727][6];				l_cell_reg[751] = inform_L[759][6];				l_cell_reg[752] = inform_L[728][6];				l_cell_reg[753] = inform_L[760][6];				l_cell_reg[754] = inform_L[729][6];				l_cell_reg[755] = inform_L[761][6];				l_cell_reg[756] = inform_L[730][6];				l_cell_reg[757] = inform_L[762][6];				l_cell_reg[758] = inform_L[731][6];				l_cell_reg[759] = inform_L[763][6];				l_cell_reg[760] = inform_L[732][6];				l_cell_reg[761] = inform_L[764][6];				l_cell_reg[762] = inform_L[733][6];				l_cell_reg[763] = inform_L[765][6];				l_cell_reg[764] = inform_L[734][6];				l_cell_reg[765] = inform_L[766][6];				l_cell_reg[766] = inform_L[735][6];				l_cell_reg[767] = inform_L[767][6];				l_cell_reg[768] = inform_L[768][6];				l_cell_reg[769] = inform_L[800][6];				l_cell_reg[770] = inform_L[769][6];				l_cell_reg[771] = inform_L[801][6];				l_cell_reg[772] = inform_L[770][6];				l_cell_reg[773] = inform_L[802][6];				l_cell_reg[774] = inform_L[771][6];				l_cell_reg[775] = inform_L[803][6];				l_cell_reg[776] = inform_L[772][6];				l_cell_reg[777] = inform_L[804][6];				l_cell_reg[778] = inform_L[773][6];				l_cell_reg[779] = inform_L[805][6];				l_cell_reg[780] = inform_L[774][6];				l_cell_reg[781] = inform_L[806][6];				l_cell_reg[782] = inform_L[775][6];				l_cell_reg[783] = inform_L[807][6];				l_cell_reg[784] = inform_L[776][6];				l_cell_reg[785] = inform_L[808][6];				l_cell_reg[786] = inform_L[777][6];				l_cell_reg[787] = inform_L[809][6];				l_cell_reg[788] = inform_L[778][6];				l_cell_reg[789] = inform_L[810][6];				l_cell_reg[790] = inform_L[779][6];				l_cell_reg[791] = inform_L[811][6];				l_cell_reg[792] = inform_L[780][6];				l_cell_reg[793] = inform_L[812][6];				l_cell_reg[794] = inform_L[781][6];				l_cell_reg[795] = inform_L[813][6];				l_cell_reg[796] = inform_L[782][6];				l_cell_reg[797] = inform_L[814][6];				l_cell_reg[798] = inform_L[783][6];				l_cell_reg[799] = inform_L[815][6];				l_cell_reg[800] = inform_L[784][6];				l_cell_reg[801] = inform_L[816][6];				l_cell_reg[802] = inform_L[785][6];				l_cell_reg[803] = inform_L[817][6];				l_cell_reg[804] = inform_L[786][6];				l_cell_reg[805] = inform_L[818][6];				l_cell_reg[806] = inform_L[787][6];				l_cell_reg[807] = inform_L[819][6];				l_cell_reg[808] = inform_L[788][6];				l_cell_reg[809] = inform_L[820][6];				l_cell_reg[810] = inform_L[789][6];				l_cell_reg[811] = inform_L[821][6];				l_cell_reg[812] = inform_L[790][6];				l_cell_reg[813] = inform_L[822][6];				l_cell_reg[814] = inform_L[791][6];				l_cell_reg[815] = inform_L[823][6];				l_cell_reg[816] = inform_L[792][6];				l_cell_reg[817] = inform_L[824][6];				l_cell_reg[818] = inform_L[793][6];				l_cell_reg[819] = inform_L[825][6];				l_cell_reg[820] = inform_L[794][6];				l_cell_reg[821] = inform_L[826][6];				l_cell_reg[822] = inform_L[795][6];				l_cell_reg[823] = inform_L[827][6];				l_cell_reg[824] = inform_L[796][6];				l_cell_reg[825] = inform_L[828][6];				l_cell_reg[826] = inform_L[797][6];				l_cell_reg[827] = inform_L[829][6];				l_cell_reg[828] = inform_L[798][6];				l_cell_reg[829] = inform_L[830][6];				l_cell_reg[830] = inform_L[799][6];				l_cell_reg[831] = inform_L[831][6];				l_cell_reg[832] = inform_L[832][6];				l_cell_reg[833] = inform_L[864][6];				l_cell_reg[834] = inform_L[833][6];				l_cell_reg[835] = inform_L[865][6];				l_cell_reg[836] = inform_L[834][6];				l_cell_reg[837] = inform_L[866][6];				l_cell_reg[838] = inform_L[835][6];				l_cell_reg[839] = inform_L[867][6];				l_cell_reg[840] = inform_L[836][6];				l_cell_reg[841] = inform_L[868][6];				l_cell_reg[842] = inform_L[837][6];				l_cell_reg[843] = inform_L[869][6];				l_cell_reg[844] = inform_L[838][6];				l_cell_reg[845] = inform_L[870][6];				l_cell_reg[846] = inform_L[839][6];				l_cell_reg[847] = inform_L[871][6];				l_cell_reg[848] = inform_L[840][6];				l_cell_reg[849] = inform_L[872][6];				l_cell_reg[850] = inform_L[841][6];				l_cell_reg[851] = inform_L[873][6];				l_cell_reg[852] = inform_L[842][6];				l_cell_reg[853] = inform_L[874][6];				l_cell_reg[854] = inform_L[843][6];				l_cell_reg[855] = inform_L[875][6];				l_cell_reg[856] = inform_L[844][6];				l_cell_reg[857] = inform_L[876][6];				l_cell_reg[858] = inform_L[845][6];				l_cell_reg[859] = inform_L[877][6];				l_cell_reg[860] = inform_L[846][6];				l_cell_reg[861] = inform_L[878][6];				l_cell_reg[862] = inform_L[847][6];				l_cell_reg[863] = inform_L[879][6];				l_cell_reg[864] = inform_L[848][6];				l_cell_reg[865] = inform_L[880][6];				l_cell_reg[866] = inform_L[849][6];				l_cell_reg[867] = inform_L[881][6];				l_cell_reg[868] = inform_L[850][6];				l_cell_reg[869] = inform_L[882][6];				l_cell_reg[870] = inform_L[851][6];				l_cell_reg[871] = inform_L[883][6];				l_cell_reg[872] = inform_L[852][6];				l_cell_reg[873] = inform_L[884][6];				l_cell_reg[874] = inform_L[853][6];				l_cell_reg[875] = inform_L[885][6];				l_cell_reg[876] = inform_L[854][6];				l_cell_reg[877] = inform_L[886][6];				l_cell_reg[878] = inform_L[855][6];				l_cell_reg[879] = inform_L[887][6];				l_cell_reg[880] = inform_L[856][6];				l_cell_reg[881] = inform_L[888][6];				l_cell_reg[882] = inform_L[857][6];				l_cell_reg[883] = inform_L[889][6];				l_cell_reg[884] = inform_L[858][6];				l_cell_reg[885] = inform_L[890][6];				l_cell_reg[886] = inform_L[859][6];				l_cell_reg[887] = inform_L[891][6];				l_cell_reg[888] = inform_L[860][6];				l_cell_reg[889] = inform_L[892][6];				l_cell_reg[890] = inform_L[861][6];				l_cell_reg[891] = inform_L[893][6];				l_cell_reg[892] = inform_L[862][6];				l_cell_reg[893] = inform_L[894][6];				l_cell_reg[894] = inform_L[863][6];				l_cell_reg[895] = inform_L[895][6];				l_cell_reg[896] = inform_L[896][6];				l_cell_reg[897] = inform_L[928][6];				l_cell_reg[898] = inform_L[897][6];				l_cell_reg[899] = inform_L[929][6];				l_cell_reg[900] = inform_L[898][6];				l_cell_reg[901] = inform_L[930][6];				l_cell_reg[902] = inform_L[899][6];				l_cell_reg[903] = inform_L[931][6];				l_cell_reg[904] = inform_L[900][6];				l_cell_reg[905] = inform_L[932][6];				l_cell_reg[906] = inform_L[901][6];				l_cell_reg[907] = inform_L[933][6];				l_cell_reg[908] = inform_L[902][6];				l_cell_reg[909] = inform_L[934][6];				l_cell_reg[910] = inform_L[903][6];				l_cell_reg[911] = inform_L[935][6];				l_cell_reg[912] = inform_L[904][6];				l_cell_reg[913] = inform_L[936][6];				l_cell_reg[914] = inform_L[905][6];				l_cell_reg[915] = inform_L[937][6];				l_cell_reg[916] = inform_L[906][6];				l_cell_reg[917] = inform_L[938][6];				l_cell_reg[918] = inform_L[907][6];				l_cell_reg[919] = inform_L[939][6];				l_cell_reg[920] = inform_L[908][6];				l_cell_reg[921] = inform_L[940][6];				l_cell_reg[922] = inform_L[909][6];				l_cell_reg[923] = inform_L[941][6];				l_cell_reg[924] = inform_L[910][6];				l_cell_reg[925] = inform_L[942][6];				l_cell_reg[926] = inform_L[911][6];				l_cell_reg[927] = inform_L[943][6];				l_cell_reg[928] = inform_L[912][6];				l_cell_reg[929] = inform_L[944][6];				l_cell_reg[930] = inform_L[913][6];				l_cell_reg[931] = inform_L[945][6];				l_cell_reg[932] = inform_L[914][6];				l_cell_reg[933] = inform_L[946][6];				l_cell_reg[934] = inform_L[915][6];				l_cell_reg[935] = inform_L[947][6];				l_cell_reg[936] = inform_L[916][6];				l_cell_reg[937] = inform_L[948][6];				l_cell_reg[938] = inform_L[917][6];				l_cell_reg[939] = inform_L[949][6];				l_cell_reg[940] = inform_L[918][6];				l_cell_reg[941] = inform_L[950][6];				l_cell_reg[942] = inform_L[919][6];				l_cell_reg[943] = inform_L[951][6];				l_cell_reg[944] = inform_L[920][6];				l_cell_reg[945] = inform_L[952][6];				l_cell_reg[946] = inform_L[921][6];				l_cell_reg[947] = inform_L[953][6];				l_cell_reg[948] = inform_L[922][6];				l_cell_reg[949] = inform_L[954][6];				l_cell_reg[950] = inform_L[923][6];				l_cell_reg[951] = inform_L[955][6];				l_cell_reg[952] = inform_L[924][6];				l_cell_reg[953] = inform_L[956][6];				l_cell_reg[954] = inform_L[925][6];				l_cell_reg[955] = inform_L[957][6];				l_cell_reg[956] = inform_L[926][6];				l_cell_reg[957] = inform_L[958][6];				l_cell_reg[958] = inform_L[927][6];				l_cell_reg[959] = inform_L[959][6];				l_cell_reg[960] = inform_L[960][6];				l_cell_reg[961] = inform_L[992][6];				l_cell_reg[962] = inform_L[961][6];				l_cell_reg[963] = inform_L[993][6];				l_cell_reg[964] = inform_L[962][6];				l_cell_reg[965] = inform_L[994][6];				l_cell_reg[966] = inform_L[963][6];				l_cell_reg[967] = inform_L[995][6];				l_cell_reg[968] = inform_L[964][6];				l_cell_reg[969] = inform_L[996][6];				l_cell_reg[970] = inform_L[965][6];				l_cell_reg[971] = inform_L[997][6];				l_cell_reg[972] = inform_L[966][6];				l_cell_reg[973] = inform_L[998][6];				l_cell_reg[974] = inform_L[967][6];				l_cell_reg[975] = inform_L[999][6];				l_cell_reg[976] = inform_L[968][6];				l_cell_reg[977] = inform_L[1000][6];				l_cell_reg[978] = inform_L[969][6];				l_cell_reg[979] = inform_L[1001][6];				l_cell_reg[980] = inform_L[970][6];				l_cell_reg[981] = inform_L[1002][6];				l_cell_reg[982] = inform_L[971][6];				l_cell_reg[983] = inform_L[1003][6];				l_cell_reg[984] = inform_L[972][6];				l_cell_reg[985] = inform_L[1004][6];				l_cell_reg[986] = inform_L[973][6];				l_cell_reg[987] = inform_L[1005][6];				l_cell_reg[988] = inform_L[974][6];				l_cell_reg[989] = inform_L[1006][6];				l_cell_reg[990] = inform_L[975][6];				l_cell_reg[991] = inform_L[1007][6];				l_cell_reg[992] = inform_L[976][6];				l_cell_reg[993] = inform_L[1008][6];				l_cell_reg[994] = inform_L[977][6];				l_cell_reg[995] = inform_L[1009][6];				l_cell_reg[996] = inform_L[978][6];				l_cell_reg[997] = inform_L[1010][6];				l_cell_reg[998] = inform_L[979][6];				l_cell_reg[999] = inform_L[1011][6];				l_cell_reg[1000] = inform_L[980][6];				l_cell_reg[1001] = inform_L[1012][6];				l_cell_reg[1002] = inform_L[981][6];				l_cell_reg[1003] = inform_L[1013][6];				l_cell_reg[1004] = inform_L[982][6];				l_cell_reg[1005] = inform_L[1014][6];				l_cell_reg[1006] = inform_L[983][6];				l_cell_reg[1007] = inform_L[1015][6];				l_cell_reg[1008] = inform_L[984][6];				l_cell_reg[1009] = inform_L[1016][6];				l_cell_reg[1010] = inform_L[985][6];				l_cell_reg[1011] = inform_L[1017][6];				l_cell_reg[1012] = inform_L[986][6];				l_cell_reg[1013] = inform_L[1018][6];				l_cell_reg[1014] = inform_L[987][6];				l_cell_reg[1015] = inform_L[1019][6];				l_cell_reg[1016] = inform_L[988][6];				l_cell_reg[1017] = inform_L[1020][6];				l_cell_reg[1018] = inform_L[989][6];				l_cell_reg[1019] = inform_L[1021][6];				l_cell_reg[1020] = inform_L[990][6];				l_cell_reg[1021] = inform_L[1022][6];				l_cell_reg[1022] = inform_L[991][6];				l_cell_reg[1023] = inform_L[1023][6];			end
			7:			begin				r_cell_reg[0] = inform_R[0][6];				r_cell_reg[1] = inform_R[64][6];				r_cell_reg[2] = inform_R[1][6];				r_cell_reg[3] = inform_R[65][6];				r_cell_reg[4] = inform_R[2][6];				r_cell_reg[5] = inform_R[66][6];				r_cell_reg[6] = inform_R[3][6];				r_cell_reg[7] = inform_R[67][6];				r_cell_reg[8] = inform_R[4][6];				r_cell_reg[9] = inform_R[68][6];				r_cell_reg[10] = inform_R[5][6];				r_cell_reg[11] = inform_R[69][6];				r_cell_reg[12] = inform_R[6][6];				r_cell_reg[13] = inform_R[70][6];				r_cell_reg[14] = inform_R[7][6];				r_cell_reg[15] = inform_R[71][6];				r_cell_reg[16] = inform_R[8][6];				r_cell_reg[17] = inform_R[72][6];				r_cell_reg[18] = inform_R[9][6];				r_cell_reg[19] = inform_R[73][6];				r_cell_reg[20] = inform_R[10][6];				r_cell_reg[21] = inform_R[74][6];				r_cell_reg[22] = inform_R[11][6];				r_cell_reg[23] = inform_R[75][6];				r_cell_reg[24] = inform_R[12][6];				r_cell_reg[25] = inform_R[76][6];				r_cell_reg[26] = inform_R[13][6];				r_cell_reg[27] = inform_R[77][6];				r_cell_reg[28] = inform_R[14][6];				r_cell_reg[29] = inform_R[78][6];				r_cell_reg[30] = inform_R[15][6];				r_cell_reg[31] = inform_R[79][6];				r_cell_reg[32] = inform_R[16][6];				r_cell_reg[33] = inform_R[80][6];				r_cell_reg[34] = inform_R[17][6];				r_cell_reg[35] = inform_R[81][6];				r_cell_reg[36] = inform_R[18][6];				r_cell_reg[37] = inform_R[82][6];				r_cell_reg[38] = inform_R[19][6];				r_cell_reg[39] = inform_R[83][6];				r_cell_reg[40] = inform_R[20][6];				r_cell_reg[41] = inform_R[84][6];				r_cell_reg[42] = inform_R[21][6];				r_cell_reg[43] = inform_R[85][6];				r_cell_reg[44] = inform_R[22][6];				r_cell_reg[45] = inform_R[86][6];				r_cell_reg[46] = inform_R[23][6];				r_cell_reg[47] = inform_R[87][6];				r_cell_reg[48] = inform_R[24][6];				r_cell_reg[49] = inform_R[88][6];				r_cell_reg[50] = inform_R[25][6];				r_cell_reg[51] = inform_R[89][6];				r_cell_reg[52] = inform_R[26][6];				r_cell_reg[53] = inform_R[90][6];				r_cell_reg[54] = inform_R[27][6];				r_cell_reg[55] = inform_R[91][6];				r_cell_reg[56] = inform_R[28][6];				r_cell_reg[57] = inform_R[92][6];				r_cell_reg[58] = inform_R[29][6];				r_cell_reg[59] = inform_R[93][6];				r_cell_reg[60] = inform_R[30][6];				r_cell_reg[61] = inform_R[94][6];				r_cell_reg[62] = inform_R[31][6];				r_cell_reg[63] = inform_R[95][6];				r_cell_reg[64] = inform_R[32][6];				r_cell_reg[65] = inform_R[96][6];				r_cell_reg[66] = inform_R[33][6];				r_cell_reg[67] = inform_R[97][6];				r_cell_reg[68] = inform_R[34][6];				r_cell_reg[69] = inform_R[98][6];				r_cell_reg[70] = inform_R[35][6];				r_cell_reg[71] = inform_R[99][6];				r_cell_reg[72] = inform_R[36][6];				r_cell_reg[73] = inform_R[100][6];				r_cell_reg[74] = inform_R[37][6];				r_cell_reg[75] = inform_R[101][6];				r_cell_reg[76] = inform_R[38][6];				r_cell_reg[77] = inform_R[102][6];				r_cell_reg[78] = inform_R[39][6];				r_cell_reg[79] = inform_R[103][6];				r_cell_reg[80] = inform_R[40][6];				r_cell_reg[81] = inform_R[104][6];				r_cell_reg[82] = inform_R[41][6];				r_cell_reg[83] = inform_R[105][6];				r_cell_reg[84] = inform_R[42][6];				r_cell_reg[85] = inform_R[106][6];				r_cell_reg[86] = inform_R[43][6];				r_cell_reg[87] = inform_R[107][6];				r_cell_reg[88] = inform_R[44][6];				r_cell_reg[89] = inform_R[108][6];				r_cell_reg[90] = inform_R[45][6];				r_cell_reg[91] = inform_R[109][6];				r_cell_reg[92] = inform_R[46][6];				r_cell_reg[93] = inform_R[110][6];				r_cell_reg[94] = inform_R[47][6];				r_cell_reg[95] = inform_R[111][6];				r_cell_reg[96] = inform_R[48][6];				r_cell_reg[97] = inform_R[112][6];				r_cell_reg[98] = inform_R[49][6];				r_cell_reg[99] = inform_R[113][6];				r_cell_reg[100] = inform_R[50][6];				r_cell_reg[101] = inform_R[114][6];				r_cell_reg[102] = inform_R[51][6];				r_cell_reg[103] = inform_R[115][6];				r_cell_reg[104] = inform_R[52][6];				r_cell_reg[105] = inform_R[116][6];				r_cell_reg[106] = inform_R[53][6];				r_cell_reg[107] = inform_R[117][6];				r_cell_reg[108] = inform_R[54][6];				r_cell_reg[109] = inform_R[118][6];				r_cell_reg[110] = inform_R[55][6];				r_cell_reg[111] = inform_R[119][6];				r_cell_reg[112] = inform_R[56][6];				r_cell_reg[113] = inform_R[120][6];				r_cell_reg[114] = inform_R[57][6];				r_cell_reg[115] = inform_R[121][6];				r_cell_reg[116] = inform_R[58][6];				r_cell_reg[117] = inform_R[122][6];				r_cell_reg[118] = inform_R[59][6];				r_cell_reg[119] = inform_R[123][6];				r_cell_reg[120] = inform_R[60][6];				r_cell_reg[121] = inform_R[124][6];				r_cell_reg[122] = inform_R[61][6];				r_cell_reg[123] = inform_R[125][6];				r_cell_reg[124] = inform_R[62][6];				r_cell_reg[125] = inform_R[126][6];				r_cell_reg[126] = inform_R[63][6];				r_cell_reg[127] = inform_R[127][6];				r_cell_reg[128] = inform_R[128][6];				r_cell_reg[129] = inform_R[192][6];				r_cell_reg[130] = inform_R[129][6];				r_cell_reg[131] = inform_R[193][6];				r_cell_reg[132] = inform_R[130][6];				r_cell_reg[133] = inform_R[194][6];				r_cell_reg[134] = inform_R[131][6];				r_cell_reg[135] = inform_R[195][6];				r_cell_reg[136] = inform_R[132][6];				r_cell_reg[137] = inform_R[196][6];				r_cell_reg[138] = inform_R[133][6];				r_cell_reg[139] = inform_R[197][6];				r_cell_reg[140] = inform_R[134][6];				r_cell_reg[141] = inform_R[198][6];				r_cell_reg[142] = inform_R[135][6];				r_cell_reg[143] = inform_R[199][6];				r_cell_reg[144] = inform_R[136][6];				r_cell_reg[145] = inform_R[200][6];				r_cell_reg[146] = inform_R[137][6];				r_cell_reg[147] = inform_R[201][6];				r_cell_reg[148] = inform_R[138][6];				r_cell_reg[149] = inform_R[202][6];				r_cell_reg[150] = inform_R[139][6];				r_cell_reg[151] = inform_R[203][6];				r_cell_reg[152] = inform_R[140][6];				r_cell_reg[153] = inform_R[204][6];				r_cell_reg[154] = inform_R[141][6];				r_cell_reg[155] = inform_R[205][6];				r_cell_reg[156] = inform_R[142][6];				r_cell_reg[157] = inform_R[206][6];				r_cell_reg[158] = inform_R[143][6];				r_cell_reg[159] = inform_R[207][6];				r_cell_reg[160] = inform_R[144][6];				r_cell_reg[161] = inform_R[208][6];				r_cell_reg[162] = inform_R[145][6];				r_cell_reg[163] = inform_R[209][6];				r_cell_reg[164] = inform_R[146][6];				r_cell_reg[165] = inform_R[210][6];				r_cell_reg[166] = inform_R[147][6];				r_cell_reg[167] = inform_R[211][6];				r_cell_reg[168] = inform_R[148][6];				r_cell_reg[169] = inform_R[212][6];				r_cell_reg[170] = inform_R[149][6];				r_cell_reg[171] = inform_R[213][6];				r_cell_reg[172] = inform_R[150][6];				r_cell_reg[173] = inform_R[214][6];				r_cell_reg[174] = inform_R[151][6];				r_cell_reg[175] = inform_R[215][6];				r_cell_reg[176] = inform_R[152][6];				r_cell_reg[177] = inform_R[216][6];				r_cell_reg[178] = inform_R[153][6];				r_cell_reg[179] = inform_R[217][6];				r_cell_reg[180] = inform_R[154][6];				r_cell_reg[181] = inform_R[218][6];				r_cell_reg[182] = inform_R[155][6];				r_cell_reg[183] = inform_R[219][6];				r_cell_reg[184] = inform_R[156][6];				r_cell_reg[185] = inform_R[220][6];				r_cell_reg[186] = inform_R[157][6];				r_cell_reg[187] = inform_R[221][6];				r_cell_reg[188] = inform_R[158][6];				r_cell_reg[189] = inform_R[222][6];				r_cell_reg[190] = inform_R[159][6];				r_cell_reg[191] = inform_R[223][6];				r_cell_reg[192] = inform_R[160][6];				r_cell_reg[193] = inform_R[224][6];				r_cell_reg[194] = inform_R[161][6];				r_cell_reg[195] = inform_R[225][6];				r_cell_reg[196] = inform_R[162][6];				r_cell_reg[197] = inform_R[226][6];				r_cell_reg[198] = inform_R[163][6];				r_cell_reg[199] = inform_R[227][6];				r_cell_reg[200] = inform_R[164][6];				r_cell_reg[201] = inform_R[228][6];				r_cell_reg[202] = inform_R[165][6];				r_cell_reg[203] = inform_R[229][6];				r_cell_reg[204] = inform_R[166][6];				r_cell_reg[205] = inform_R[230][6];				r_cell_reg[206] = inform_R[167][6];				r_cell_reg[207] = inform_R[231][6];				r_cell_reg[208] = inform_R[168][6];				r_cell_reg[209] = inform_R[232][6];				r_cell_reg[210] = inform_R[169][6];				r_cell_reg[211] = inform_R[233][6];				r_cell_reg[212] = inform_R[170][6];				r_cell_reg[213] = inform_R[234][6];				r_cell_reg[214] = inform_R[171][6];				r_cell_reg[215] = inform_R[235][6];				r_cell_reg[216] = inform_R[172][6];				r_cell_reg[217] = inform_R[236][6];				r_cell_reg[218] = inform_R[173][6];				r_cell_reg[219] = inform_R[237][6];				r_cell_reg[220] = inform_R[174][6];				r_cell_reg[221] = inform_R[238][6];				r_cell_reg[222] = inform_R[175][6];				r_cell_reg[223] = inform_R[239][6];				r_cell_reg[224] = inform_R[176][6];				r_cell_reg[225] = inform_R[240][6];				r_cell_reg[226] = inform_R[177][6];				r_cell_reg[227] = inform_R[241][6];				r_cell_reg[228] = inform_R[178][6];				r_cell_reg[229] = inform_R[242][6];				r_cell_reg[230] = inform_R[179][6];				r_cell_reg[231] = inform_R[243][6];				r_cell_reg[232] = inform_R[180][6];				r_cell_reg[233] = inform_R[244][6];				r_cell_reg[234] = inform_R[181][6];				r_cell_reg[235] = inform_R[245][6];				r_cell_reg[236] = inform_R[182][6];				r_cell_reg[237] = inform_R[246][6];				r_cell_reg[238] = inform_R[183][6];				r_cell_reg[239] = inform_R[247][6];				r_cell_reg[240] = inform_R[184][6];				r_cell_reg[241] = inform_R[248][6];				r_cell_reg[242] = inform_R[185][6];				r_cell_reg[243] = inform_R[249][6];				r_cell_reg[244] = inform_R[186][6];				r_cell_reg[245] = inform_R[250][6];				r_cell_reg[246] = inform_R[187][6];				r_cell_reg[247] = inform_R[251][6];				r_cell_reg[248] = inform_R[188][6];				r_cell_reg[249] = inform_R[252][6];				r_cell_reg[250] = inform_R[189][6];				r_cell_reg[251] = inform_R[253][6];				r_cell_reg[252] = inform_R[190][6];				r_cell_reg[253] = inform_R[254][6];				r_cell_reg[254] = inform_R[191][6];				r_cell_reg[255] = inform_R[255][6];				r_cell_reg[256] = inform_R[256][6];				r_cell_reg[257] = inform_R[320][6];				r_cell_reg[258] = inform_R[257][6];				r_cell_reg[259] = inform_R[321][6];				r_cell_reg[260] = inform_R[258][6];				r_cell_reg[261] = inform_R[322][6];				r_cell_reg[262] = inform_R[259][6];				r_cell_reg[263] = inform_R[323][6];				r_cell_reg[264] = inform_R[260][6];				r_cell_reg[265] = inform_R[324][6];				r_cell_reg[266] = inform_R[261][6];				r_cell_reg[267] = inform_R[325][6];				r_cell_reg[268] = inform_R[262][6];				r_cell_reg[269] = inform_R[326][6];				r_cell_reg[270] = inform_R[263][6];				r_cell_reg[271] = inform_R[327][6];				r_cell_reg[272] = inform_R[264][6];				r_cell_reg[273] = inform_R[328][6];				r_cell_reg[274] = inform_R[265][6];				r_cell_reg[275] = inform_R[329][6];				r_cell_reg[276] = inform_R[266][6];				r_cell_reg[277] = inform_R[330][6];				r_cell_reg[278] = inform_R[267][6];				r_cell_reg[279] = inform_R[331][6];				r_cell_reg[280] = inform_R[268][6];				r_cell_reg[281] = inform_R[332][6];				r_cell_reg[282] = inform_R[269][6];				r_cell_reg[283] = inform_R[333][6];				r_cell_reg[284] = inform_R[270][6];				r_cell_reg[285] = inform_R[334][6];				r_cell_reg[286] = inform_R[271][6];				r_cell_reg[287] = inform_R[335][6];				r_cell_reg[288] = inform_R[272][6];				r_cell_reg[289] = inform_R[336][6];				r_cell_reg[290] = inform_R[273][6];				r_cell_reg[291] = inform_R[337][6];				r_cell_reg[292] = inform_R[274][6];				r_cell_reg[293] = inform_R[338][6];				r_cell_reg[294] = inform_R[275][6];				r_cell_reg[295] = inform_R[339][6];				r_cell_reg[296] = inform_R[276][6];				r_cell_reg[297] = inform_R[340][6];				r_cell_reg[298] = inform_R[277][6];				r_cell_reg[299] = inform_R[341][6];				r_cell_reg[300] = inform_R[278][6];				r_cell_reg[301] = inform_R[342][6];				r_cell_reg[302] = inform_R[279][6];				r_cell_reg[303] = inform_R[343][6];				r_cell_reg[304] = inform_R[280][6];				r_cell_reg[305] = inform_R[344][6];				r_cell_reg[306] = inform_R[281][6];				r_cell_reg[307] = inform_R[345][6];				r_cell_reg[308] = inform_R[282][6];				r_cell_reg[309] = inform_R[346][6];				r_cell_reg[310] = inform_R[283][6];				r_cell_reg[311] = inform_R[347][6];				r_cell_reg[312] = inform_R[284][6];				r_cell_reg[313] = inform_R[348][6];				r_cell_reg[314] = inform_R[285][6];				r_cell_reg[315] = inform_R[349][6];				r_cell_reg[316] = inform_R[286][6];				r_cell_reg[317] = inform_R[350][6];				r_cell_reg[318] = inform_R[287][6];				r_cell_reg[319] = inform_R[351][6];				r_cell_reg[320] = inform_R[288][6];				r_cell_reg[321] = inform_R[352][6];				r_cell_reg[322] = inform_R[289][6];				r_cell_reg[323] = inform_R[353][6];				r_cell_reg[324] = inform_R[290][6];				r_cell_reg[325] = inform_R[354][6];				r_cell_reg[326] = inform_R[291][6];				r_cell_reg[327] = inform_R[355][6];				r_cell_reg[328] = inform_R[292][6];				r_cell_reg[329] = inform_R[356][6];				r_cell_reg[330] = inform_R[293][6];				r_cell_reg[331] = inform_R[357][6];				r_cell_reg[332] = inform_R[294][6];				r_cell_reg[333] = inform_R[358][6];				r_cell_reg[334] = inform_R[295][6];				r_cell_reg[335] = inform_R[359][6];				r_cell_reg[336] = inform_R[296][6];				r_cell_reg[337] = inform_R[360][6];				r_cell_reg[338] = inform_R[297][6];				r_cell_reg[339] = inform_R[361][6];				r_cell_reg[340] = inform_R[298][6];				r_cell_reg[341] = inform_R[362][6];				r_cell_reg[342] = inform_R[299][6];				r_cell_reg[343] = inform_R[363][6];				r_cell_reg[344] = inform_R[300][6];				r_cell_reg[345] = inform_R[364][6];				r_cell_reg[346] = inform_R[301][6];				r_cell_reg[347] = inform_R[365][6];				r_cell_reg[348] = inform_R[302][6];				r_cell_reg[349] = inform_R[366][6];				r_cell_reg[350] = inform_R[303][6];				r_cell_reg[351] = inform_R[367][6];				r_cell_reg[352] = inform_R[304][6];				r_cell_reg[353] = inform_R[368][6];				r_cell_reg[354] = inform_R[305][6];				r_cell_reg[355] = inform_R[369][6];				r_cell_reg[356] = inform_R[306][6];				r_cell_reg[357] = inform_R[370][6];				r_cell_reg[358] = inform_R[307][6];				r_cell_reg[359] = inform_R[371][6];				r_cell_reg[360] = inform_R[308][6];				r_cell_reg[361] = inform_R[372][6];				r_cell_reg[362] = inform_R[309][6];				r_cell_reg[363] = inform_R[373][6];				r_cell_reg[364] = inform_R[310][6];				r_cell_reg[365] = inform_R[374][6];				r_cell_reg[366] = inform_R[311][6];				r_cell_reg[367] = inform_R[375][6];				r_cell_reg[368] = inform_R[312][6];				r_cell_reg[369] = inform_R[376][6];				r_cell_reg[370] = inform_R[313][6];				r_cell_reg[371] = inform_R[377][6];				r_cell_reg[372] = inform_R[314][6];				r_cell_reg[373] = inform_R[378][6];				r_cell_reg[374] = inform_R[315][6];				r_cell_reg[375] = inform_R[379][6];				r_cell_reg[376] = inform_R[316][6];				r_cell_reg[377] = inform_R[380][6];				r_cell_reg[378] = inform_R[317][6];				r_cell_reg[379] = inform_R[381][6];				r_cell_reg[380] = inform_R[318][6];				r_cell_reg[381] = inform_R[382][6];				r_cell_reg[382] = inform_R[319][6];				r_cell_reg[383] = inform_R[383][6];				r_cell_reg[384] = inform_R[384][6];				r_cell_reg[385] = inform_R[448][6];				r_cell_reg[386] = inform_R[385][6];				r_cell_reg[387] = inform_R[449][6];				r_cell_reg[388] = inform_R[386][6];				r_cell_reg[389] = inform_R[450][6];				r_cell_reg[390] = inform_R[387][6];				r_cell_reg[391] = inform_R[451][6];				r_cell_reg[392] = inform_R[388][6];				r_cell_reg[393] = inform_R[452][6];				r_cell_reg[394] = inform_R[389][6];				r_cell_reg[395] = inform_R[453][6];				r_cell_reg[396] = inform_R[390][6];				r_cell_reg[397] = inform_R[454][6];				r_cell_reg[398] = inform_R[391][6];				r_cell_reg[399] = inform_R[455][6];				r_cell_reg[400] = inform_R[392][6];				r_cell_reg[401] = inform_R[456][6];				r_cell_reg[402] = inform_R[393][6];				r_cell_reg[403] = inform_R[457][6];				r_cell_reg[404] = inform_R[394][6];				r_cell_reg[405] = inform_R[458][6];				r_cell_reg[406] = inform_R[395][6];				r_cell_reg[407] = inform_R[459][6];				r_cell_reg[408] = inform_R[396][6];				r_cell_reg[409] = inform_R[460][6];				r_cell_reg[410] = inform_R[397][6];				r_cell_reg[411] = inform_R[461][6];				r_cell_reg[412] = inform_R[398][6];				r_cell_reg[413] = inform_R[462][6];				r_cell_reg[414] = inform_R[399][6];				r_cell_reg[415] = inform_R[463][6];				r_cell_reg[416] = inform_R[400][6];				r_cell_reg[417] = inform_R[464][6];				r_cell_reg[418] = inform_R[401][6];				r_cell_reg[419] = inform_R[465][6];				r_cell_reg[420] = inform_R[402][6];				r_cell_reg[421] = inform_R[466][6];				r_cell_reg[422] = inform_R[403][6];				r_cell_reg[423] = inform_R[467][6];				r_cell_reg[424] = inform_R[404][6];				r_cell_reg[425] = inform_R[468][6];				r_cell_reg[426] = inform_R[405][6];				r_cell_reg[427] = inform_R[469][6];				r_cell_reg[428] = inform_R[406][6];				r_cell_reg[429] = inform_R[470][6];				r_cell_reg[430] = inform_R[407][6];				r_cell_reg[431] = inform_R[471][6];				r_cell_reg[432] = inform_R[408][6];				r_cell_reg[433] = inform_R[472][6];				r_cell_reg[434] = inform_R[409][6];				r_cell_reg[435] = inform_R[473][6];				r_cell_reg[436] = inform_R[410][6];				r_cell_reg[437] = inform_R[474][6];				r_cell_reg[438] = inform_R[411][6];				r_cell_reg[439] = inform_R[475][6];				r_cell_reg[440] = inform_R[412][6];				r_cell_reg[441] = inform_R[476][6];				r_cell_reg[442] = inform_R[413][6];				r_cell_reg[443] = inform_R[477][6];				r_cell_reg[444] = inform_R[414][6];				r_cell_reg[445] = inform_R[478][6];				r_cell_reg[446] = inform_R[415][6];				r_cell_reg[447] = inform_R[479][6];				r_cell_reg[448] = inform_R[416][6];				r_cell_reg[449] = inform_R[480][6];				r_cell_reg[450] = inform_R[417][6];				r_cell_reg[451] = inform_R[481][6];				r_cell_reg[452] = inform_R[418][6];				r_cell_reg[453] = inform_R[482][6];				r_cell_reg[454] = inform_R[419][6];				r_cell_reg[455] = inform_R[483][6];				r_cell_reg[456] = inform_R[420][6];				r_cell_reg[457] = inform_R[484][6];				r_cell_reg[458] = inform_R[421][6];				r_cell_reg[459] = inform_R[485][6];				r_cell_reg[460] = inform_R[422][6];				r_cell_reg[461] = inform_R[486][6];				r_cell_reg[462] = inform_R[423][6];				r_cell_reg[463] = inform_R[487][6];				r_cell_reg[464] = inform_R[424][6];				r_cell_reg[465] = inform_R[488][6];				r_cell_reg[466] = inform_R[425][6];				r_cell_reg[467] = inform_R[489][6];				r_cell_reg[468] = inform_R[426][6];				r_cell_reg[469] = inform_R[490][6];				r_cell_reg[470] = inform_R[427][6];				r_cell_reg[471] = inform_R[491][6];				r_cell_reg[472] = inform_R[428][6];				r_cell_reg[473] = inform_R[492][6];				r_cell_reg[474] = inform_R[429][6];				r_cell_reg[475] = inform_R[493][6];				r_cell_reg[476] = inform_R[430][6];				r_cell_reg[477] = inform_R[494][6];				r_cell_reg[478] = inform_R[431][6];				r_cell_reg[479] = inform_R[495][6];				r_cell_reg[480] = inform_R[432][6];				r_cell_reg[481] = inform_R[496][6];				r_cell_reg[482] = inform_R[433][6];				r_cell_reg[483] = inform_R[497][6];				r_cell_reg[484] = inform_R[434][6];				r_cell_reg[485] = inform_R[498][6];				r_cell_reg[486] = inform_R[435][6];				r_cell_reg[487] = inform_R[499][6];				r_cell_reg[488] = inform_R[436][6];				r_cell_reg[489] = inform_R[500][6];				r_cell_reg[490] = inform_R[437][6];				r_cell_reg[491] = inform_R[501][6];				r_cell_reg[492] = inform_R[438][6];				r_cell_reg[493] = inform_R[502][6];				r_cell_reg[494] = inform_R[439][6];				r_cell_reg[495] = inform_R[503][6];				r_cell_reg[496] = inform_R[440][6];				r_cell_reg[497] = inform_R[504][6];				r_cell_reg[498] = inform_R[441][6];				r_cell_reg[499] = inform_R[505][6];				r_cell_reg[500] = inform_R[442][6];				r_cell_reg[501] = inform_R[506][6];				r_cell_reg[502] = inform_R[443][6];				r_cell_reg[503] = inform_R[507][6];				r_cell_reg[504] = inform_R[444][6];				r_cell_reg[505] = inform_R[508][6];				r_cell_reg[506] = inform_R[445][6];				r_cell_reg[507] = inform_R[509][6];				r_cell_reg[508] = inform_R[446][6];				r_cell_reg[509] = inform_R[510][6];				r_cell_reg[510] = inform_R[447][6];				r_cell_reg[511] = inform_R[511][6];				r_cell_reg[512] = inform_R[512][6];				r_cell_reg[513] = inform_R[576][6];				r_cell_reg[514] = inform_R[513][6];				r_cell_reg[515] = inform_R[577][6];				r_cell_reg[516] = inform_R[514][6];				r_cell_reg[517] = inform_R[578][6];				r_cell_reg[518] = inform_R[515][6];				r_cell_reg[519] = inform_R[579][6];				r_cell_reg[520] = inform_R[516][6];				r_cell_reg[521] = inform_R[580][6];				r_cell_reg[522] = inform_R[517][6];				r_cell_reg[523] = inform_R[581][6];				r_cell_reg[524] = inform_R[518][6];				r_cell_reg[525] = inform_R[582][6];				r_cell_reg[526] = inform_R[519][6];				r_cell_reg[527] = inform_R[583][6];				r_cell_reg[528] = inform_R[520][6];				r_cell_reg[529] = inform_R[584][6];				r_cell_reg[530] = inform_R[521][6];				r_cell_reg[531] = inform_R[585][6];				r_cell_reg[532] = inform_R[522][6];				r_cell_reg[533] = inform_R[586][6];				r_cell_reg[534] = inform_R[523][6];				r_cell_reg[535] = inform_R[587][6];				r_cell_reg[536] = inform_R[524][6];				r_cell_reg[537] = inform_R[588][6];				r_cell_reg[538] = inform_R[525][6];				r_cell_reg[539] = inform_R[589][6];				r_cell_reg[540] = inform_R[526][6];				r_cell_reg[541] = inform_R[590][6];				r_cell_reg[542] = inform_R[527][6];				r_cell_reg[543] = inform_R[591][6];				r_cell_reg[544] = inform_R[528][6];				r_cell_reg[545] = inform_R[592][6];				r_cell_reg[546] = inform_R[529][6];				r_cell_reg[547] = inform_R[593][6];				r_cell_reg[548] = inform_R[530][6];				r_cell_reg[549] = inform_R[594][6];				r_cell_reg[550] = inform_R[531][6];				r_cell_reg[551] = inform_R[595][6];				r_cell_reg[552] = inform_R[532][6];				r_cell_reg[553] = inform_R[596][6];				r_cell_reg[554] = inform_R[533][6];				r_cell_reg[555] = inform_R[597][6];				r_cell_reg[556] = inform_R[534][6];				r_cell_reg[557] = inform_R[598][6];				r_cell_reg[558] = inform_R[535][6];				r_cell_reg[559] = inform_R[599][6];				r_cell_reg[560] = inform_R[536][6];				r_cell_reg[561] = inform_R[600][6];				r_cell_reg[562] = inform_R[537][6];				r_cell_reg[563] = inform_R[601][6];				r_cell_reg[564] = inform_R[538][6];				r_cell_reg[565] = inform_R[602][6];				r_cell_reg[566] = inform_R[539][6];				r_cell_reg[567] = inform_R[603][6];				r_cell_reg[568] = inform_R[540][6];				r_cell_reg[569] = inform_R[604][6];				r_cell_reg[570] = inform_R[541][6];				r_cell_reg[571] = inform_R[605][6];				r_cell_reg[572] = inform_R[542][6];				r_cell_reg[573] = inform_R[606][6];				r_cell_reg[574] = inform_R[543][6];				r_cell_reg[575] = inform_R[607][6];				r_cell_reg[576] = inform_R[544][6];				r_cell_reg[577] = inform_R[608][6];				r_cell_reg[578] = inform_R[545][6];				r_cell_reg[579] = inform_R[609][6];				r_cell_reg[580] = inform_R[546][6];				r_cell_reg[581] = inform_R[610][6];				r_cell_reg[582] = inform_R[547][6];				r_cell_reg[583] = inform_R[611][6];				r_cell_reg[584] = inform_R[548][6];				r_cell_reg[585] = inform_R[612][6];				r_cell_reg[586] = inform_R[549][6];				r_cell_reg[587] = inform_R[613][6];				r_cell_reg[588] = inform_R[550][6];				r_cell_reg[589] = inform_R[614][6];				r_cell_reg[590] = inform_R[551][6];				r_cell_reg[591] = inform_R[615][6];				r_cell_reg[592] = inform_R[552][6];				r_cell_reg[593] = inform_R[616][6];				r_cell_reg[594] = inform_R[553][6];				r_cell_reg[595] = inform_R[617][6];				r_cell_reg[596] = inform_R[554][6];				r_cell_reg[597] = inform_R[618][6];				r_cell_reg[598] = inform_R[555][6];				r_cell_reg[599] = inform_R[619][6];				r_cell_reg[600] = inform_R[556][6];				r_cell_reg[601] = inform_R[620][6];				r_cell_reg[602] = inform_R[557][6];				r_cell_reg[603] = inform_R[621][6];				r_cell_reg[604] = inform_R[558][6];				r_cell_reg[605] = inform_R[622][6];				r_cell_reg[606] = inform_R[559][6];				r_cell_reg[607] = inform_R[623][6];				r_cell_reg[608] = inform_R[560][6];				r_cell_reg[609] = inform_R[624][6];				r_cell_reg[610] = inform_R[561][6];				r_cell_reg[611] = inform_R[625][6];				r_cell_reg[612] = inform_R[562][6];				r_cell_reg[613] = inform_R[626][6];				r_cell_reg[614] = inform_R[563][6];				r_cell_reg[615] = inform_R[627][6];				r_cell_reg[616] = inform_R[564][6];				r_cell_reg[617] = inform_R[628][6];				r_cell_reg[618] = inform_R[565][6];				r_cell_reg[619] = inform_R[629][6];				r_cell_reg[620] = inform_R[566][6];				r_cell_reg[621] = inform_R[630][6];				r_cell_reg[622] = inform_R[567][6];				r_cell_reg[623] = inform_R[631][6];				r_cell_reg[624] = inform_R[568][6];				r_cell_reg[625] = inform_R[632][6];				r_cell_reg[626] = inform_R[569][6];				r_cell_reg[627] = inform_R[633][6];				r_cell_reg[628] = inform_R[570][6];				r_cell_reg[629] = inform_R[634][6];				r_cell_reg[630] = inform_R[571][6];				r_cell_reg[631] = inform_R[635][6];				r_cell_reg[632] = inform_R[572][6];				r_cell_reg[633] = inform_R[636][6];				r_cell_reg[634] = inform_R[573][6];				r_cell_reg[635] = inform_R[637][6];				r_cell_reg[636] = inform_R[574][6];				r_cell_reg[637] = inform_R[638][6];				r_cell_reg[638] = inform_R[575][6];				r_cell_reg[639] = inform_R[639][6];				r_cell_reg[640] = inform_R[640][6];				r_cell_reg[641] = inform_R[704][6];				r_cell_reg[642] = inform_R[641][6];				r_cell_reg[643] = inform_R[705][6];				r_cell_reg[644] = inform_R[642][6];				r_cell_reg[645] = inform_R[706][6];				r_cell_reg[646] = inform_R[643][6];				r_cell_reg[647] = inform_R[707][6];				r_cell_reg[648] = inform_R[644][6];				r_cell_reg[649] = inform_R[708][6];				r_cell_reg[650] = inform_R[645][6];				r_cell_reg[651] = inform_R[709][6];				r_cell_reg[652] = inform_R[646][6];				r_cell_reg[653] = inform_R[710][6];				r_cell_reg[654] = inform_R[647][6];				r_cell_reg[655] = inform_R[711][6];				r_cell_reg[656] = inform_R[648][6];				r_cell_reg[657] = inform_R[712][6];				r_cell_reg[658] = inform_R[649][6];				r_cell_reg[659] = inform_R[713][6];				r_cell_reg[660] = inform_R[650][6];				r_cell_reg[661] = inform_R[714][6];				r_cell_reg[662] = inform_R[651][6];				r_cell_reg[663] = inform_R[715][6];				r_cell_reg[664] = inform_R[652][6];				r_cell_reg[665] = inform_R[716][6];				r_cell_reg[666] = inform_R[653][6];				r_cell_reg[667] = inform_R[717][6];				r_cell_reg[668] = inform_R[654][6];				r_cell_reg[669] = inform_R[718][6];				r_cell_reg[670] = inform_R[655][6];				r_cell_reg[671] = inform_R[719][6];				r_cell_reg[672] = inform_R[656][6];				r_cell_reg[673] = inform_R[720][6];				r_cell_reg[674] = inform_R[657][6];				r_cell_reg[675] = inform_R[721][6];				r_cell_reg[676] = inform_R[658][6];				r_cell_reg[677] = inform_R[722][6];				r_cell_reg[678] = inform_R[659][6];				r_cell_reg[679] = inform_R[723][6];				r_cell_reg[680] = inform_R[660][6];				r_cell_reg[681] = inform_R[724][6];				r_cell_reg[682] = inform_R[661][6];				r_cell_reg[683] = inform_R[725][6];				r_cell_reg[684] = inform_R[662][6];				r_cell_reg[685] = inform_R[726][6];				r_cell_reg[686] = inform_R[663][6];				r_cell_reg[687] = inform_R[727][6];				r_cell_reg[688] = inform_R[664][6];				r_cell_reg[689] = inform_R[728][6];				r_cell_reg[690] = inform_R[665][6];				r_cell_reg[691] = inform_R[729][6];				r_cell_reg[692] = inform_R[666][6];				r_cell_reg[693] = inform_R[730][6];				r_cell_reg[694] = inform_R[667][6];				r_cell_reg[695] = inform_R[731][6];				r_cell_reg[696] = inform_R[668][6];				r_cell_reg[697] = inform_R[732][6];				r_cell_reg[698] = inform_R[669][6];				r_cell_reg[699] = inform_R[733][6];				r_cell_reg[700] = inform_R[670][6];				r_cell_reg[701] = inform_R[734][6];				r_cell_reg[702] = inform_R[671][6];				r_cell_reg[703] = inform_R[735][6];				r_cell_reg[704] = inform_R[672][6];				r_cell_reg[705] = inform_R[736][6];				r_cell_reg[706] = inform_R[673][6];				r_cell_reg[707] = inform_R[737][6];				r_cell_reg[708] = inform_R[674][6];				r_cell_reg[709] = inform_R[738][6];				r_cell_reg[710] = inform_R[675][6];				r_cell_reg[711] = inform_R[739][6];				r_cell_reg[712] = inform_R[676][6];				r_cell_reg[713] = inform_R[740][6];				r_cell_reg[714] = inform_R[677][6];				r_cell_reg[715] = inform_R[741][6];				r_cell_reg[716] = inform_R[678][6];				r_cell_reg[717] = inform_R[742][6];				r_cell_reg[718] = inform_R[679][6];				r_cell_reg[719] = inform_R[743][6];				r_cell_reg[720] = inform_R[680][6];				r_cell_reg[721] = inform_R[744][6];				r_cell_reg[722] = inform_R[681][6];				r_cell_reg[723] = inform_R[745][6];				r_cell_reg[724] = inform_R[682][6];				r_cell_reg[725] = inform_R[746][6];				r_cell_reg[726] = inform_R[683][6];				r_cell_reg[727] = inform_R[747][6];				r_cell_reg[728] = inform_R[684][6];				r_cell_reg[729] = inform_R[748][6];				r_cell_reg[730] = inform_R[685][6];				r_cell_reg[731] = inform_R[749][6];				r_cell_reg[732] = inform_R[686][6];				r_cell_reg[733] = inform_R[750][6];				r_cell_reg[734] = inform_R[687][6];				r_cell_reg[735] = inform_R[751][6];				r_cell_reg[736] = inform_R[688][6];				r_cell_reg[737] = inform_R[752][6];				r_cell_reg[738] = inform_R[689][6];				r_cell_reg[739] = inform_R[753][6];				r_cell_reg[740] = inform_R[690][6];				r_cell_reg[741] = inform_R[754][6];				r_cell_reg[742] = inform_R[691][6];				r_cell_reg[743] = inform_R[755][6];				r_cell_reg[744] = inform_R[692][6];				r_cell_reg[745] = inform_R[756][6];				r_cell_reg[746] = inform_R[693][6];				r_cell_reg[747] = inform_R[757][6];				r_cell_reg[748] = inform_R[694][6];				r_cell_reg[749] = inform_R[758][6];				r_cell_reg[750] = inform_R[695][6];				r_cell_reg[751] = inform_R[759][6];				r_cell_reg[752] = inform_R[696][6];				r_cell_reg[753] = inform_R[760][6];				r_cell_reg[754] = inform_R[697][6];				r_cell_reg[755] = inform_R[761][6];				r_cell_reg[756] = inform_R[698][6];				r_cell_reg[757] = inform_R[762][6];				r_cell_reg[758] = inform_R[699][6];				r_cell_reg[759] = inform_R[763][6];				r_cell_reg[760] = inform_R[700][6];				r_cell_reg[761] = inform_R[764][6];				r_cell_reg[762] = inform_R[701][6];				r_cell_reg[763] = inform_R[765][6];				r_cell_reg[764] = inform_R[702][6];				r_cell_reg[765] = inform_R[766][6];				r_cell_reg[766] = inform_R[703][6];				r_cell_reg[767] = inform_R[767][6];				r_cell_reg[768] = inform_R[768][6];				r_cell_reg[769] = inform_R[832][6];				r_cell_reg[770] = inform_R[769][6];				r_cell_reg[771] = inform_R[833][6];				r_cell_reg[772] = inform_R[770][6];				r_cell_reg[773] = inform_R[834][6];				r_cell_reg[774] = inform_R[771][6];				r_cell_reg[775] = inform_R[835][6];				r_cell_reg[776] = inform_R[772][6];				r_cell_reg[777] = inform_R[836][6];				r_cell_reg[778] = inform_R[773][6];				r_cell_reg[779] = inform_R[837][6];				r_cell_reg[780] = inform_R[774][6];				r_cell_reg[781] = inform_R[838][6];				r_cell_reg[782] = inform_R[775][6];				r_cell_reg[783] = inform_R[839][6];				r_cell_reg[784] = inform_R[776][6];				r_cell_reg[785] = inform_R[840][6];				r_cell_reg[786] = inform_R[777][6];				r_cell_reg[787] = inform_R[841][6];				r_cell_reg[788] = inform_R[778][6];				r_cell_reg[789] = inform_R[842][6];				r_cell_reg[790] = inform_R[779][6];				r_cell_reg[791] = inform_R[843][6];				r_cell_reg[792] = inform_R[780][6];				r_cell_reg[793] = inform_R[844][6];				r_cell_reg[794] = inform_R[781][6];				r_cell_reg[795] = inform_R[845][6];				r_cell_reg[796] = inform_R[782][6];				r_cell_reg[797] = inform_R[846][6];				r_cell_reg[798] = inform_R[783][6];				r_cell_reg[799] = inform_R[847][6];				r_cell_reg[800] = inform_R[784][6];				r_cell_reg[801] = inform_R[848][6];				r_cell_reg[802] = inform_R[785][6];				r_cell_reg[803] = inform_R[849][6];				r_cell_reg[804] = inform_R[786][6];				r_cell_reg[805] = inform_R[850][6];				r_cell_reg[806] = inform_R[787][6];				r_cell_reg[807] = inform_R[851][6];				r_cell_reg[808] = inform_R[788][6];				r_cell_reg[809] = inform_R[852][6];				r_cell_reg[810] = inform_R[789][6];				r_cell_reg[811] = inform_R[853][6];				r_cell_reg[812] = inform_R[790][6];				r_cell_reg[813] = inform_R[854][6];				r_cell_reg[814] = inform_R[791][6];				r_cell_reg[815] = inform_R[855][6];				r_cell_reg[816] = inform_R[792][6];				r_cell_reg[817] = inform_R[856][6];				r_cell_reg[818] = inform_R[793][6];				r_cell_reg[819] = inform_R[857][6];				r_cell_reg[820] = inform_R[794][6];				r_cell_reg[821] = inform_R[858][6];				r_cell_reg[822] = inform_R[795][6];				r_cell_reg[823] = inform_R[859][6];				r_cell_reg[824] = inform_R[796][6];				r_cell_reg[825] = inform_R[860][6];				r_cell_reg[826] = inform_R[797][6];				r_cell_reg[827] = inform_R[861][6];				r_cell_reg[828] = inform_R[798][6];				r_cell_reg[829] = inform_R[862][6];				r_cell_reg[830] = inform_R[799][6];				r_cell_reg[831] = inform_R[863][6];				r_cell_reg[832] = inform_R[800][6];				r_cell_reg[833] = inform_R[864][6];				r_cell_reg[834] = inform_R[801][6];				r_cell_reg[835] = inform_R[865][6];				r_cell_reg[836] = inform_R[802][6];				r_cell_reg[837] = inform_R[866][6];				r_cell_reg[838] = inform_R[803][6];				r_cell_reg[839] = inform_R[867][6];				r_cell_reg[840] = inform_R[804][6];				r_cell_reg[841] = inform_R[868][6];				r_cell_reg[842] = inform_R[805][6];				r_cell_reg[843] = inform_R[869][6];				r_cell_reg[844] = inform_R[806][6];				r_cell_reg[845] = inform_R[870][6];				r_cell_reg[846] = inform_R[807][6];				r_cell_reg[847] = inform_R[871][6];				r_cell_reg[848] = inform_R[808][6];				r_cell_reg[849] = inform_R[872][6];				r_cell_reg[850] = inform_R[809][6];				r_cell_reg[851] = inform_R[873][6];				r_cell_reg[852] = inform_R[810][6];				r_cell_reg[853] = inform_R[874][6];				r_cell_reg[854] = inform_R[811][6];				r_cell_reg[855] = inform_R[875][6];				r_cell_reg[856] = inform_R[812][6];				r_cell_reg[857] = inform_R[876][6];				r_cell_reg[858] = inform_R[813][6];				r_cell_reg[859] = inform_R[877][6];				r_cell_reg[860] = inform_R[814][6];				r_cell_reg[861] = inform_R[878][6];				r_cell_reg[862] = inform_R[815][6];				r_cell_reg[863] = inform_R[879][6];				r_cell_reg[864] = inform_R[816][6];				r_cell_reg[865] = inform_R[880][6];				r_cell_reg[866] = inform_R[817][6];				r_cell_reg[867] = inform_R[881][6];				r_cell_reg[868] = inform_R[818][6];				r_cell_reg[869] = inform_R[882][6];				r_cell_reg[870] = inform_R[819][6];				r_cell_reg[871] = inform_R[883][6];				r_cell_reg[872] = inform_R[820][6];				r_cell_reg[873] = inform_R[884][6];				r_cell_reg[874] = inform_R[821][6];				r_cell_reg[875] = inform_R[885][6];				r_cell_reg[876] = inform_R[822][6];				r_cell_reg[877] = inform_R[886][6];				r_cell_reg[878] = inform_R[823][6];				r_cell_reg[879] = inform_R[887][6];				r_cell_reg[880] = inform_R[824][6];				r_cell_reg[881] = inform_R[888][6];				r_cell_reg[882] = inform_R[825][6];				r_cell_reg[883] = inform_R[889][6];				r_cell_reg[884] = inform_R[826][6];				r_cell_reg[885] = inform_R[890][6];				r_cell_reg[886] = inform_R[827][6];				r_cell_reg[887] = inform_R[891][6];				r_cell_reg[888] = inform_R[828][6];				r_cell_reg[889] = inform_R[892][6];				r_cell_reg[890] = inform_R[829][6];				r_cell_reg[891] = inform_R[893][6];				r_cell_reg[892] = inform_R[830][6];				r_cell_reg[893] = inform_R[894][6];				r_cell_reg[894] = inform_R[831][6];				r_cell_reg[895] = inform_R[895][6];				r_cell_reg[896] = inform_R[896][6];				r_cell_reg[897] = inform_R[960][6];				r_cell_reg[898] = inform_R[897][6];				r_cell_reg[899] = inform_R[961][6];				r_cell_reg[900] = inform_R[898][6];				r_cell_reg[901] = inform_R[962][6];				r_cell_reg[902] = inform_R[899][6];				r_cell_reg[903] = inform_R[963][6];				r_cell_reg[904] = inform_R[900][6];				r_cell_reg[905] = inform_R[964][6];				r_cell_reg[906] = inform_R[901][6];				r_cell_reg[907] = inform_R[965][6];				r_cell_reg[908] = inform_R[902][6];				r_cell_reg[909] = inform_R[966][6];				r_cell_reg[910] = inform_R[903][6];				r_cell_reg[911] = inform_R[967][6];				r_cell_reg[912] = inform_R[904][6];				r_cell_reg[913] = inform_R[968][6];				r_cell_reg[914] = inform_R[905][6];				r_cell_reg[915] = inform_R[969][6];				r_cell_reg[916] = inform_R[906][6];				r_cell_reg[917] = inform_R[970][6];				r_cell_reg[918] = inform_R[907][6];				r_cell_reg[919] = inform_R[971][6];				r_cell_reg[920] = inform_R[908][6];				r_cell_reg[921] = inform_R[972][6];				r_cell_reg[922] = inform_R[909][6];				r_cell_reg[923] = inform_R[973][6];				r_cell_reg[924] = inform_R[910][6];				r_cell_reg[925] = inform_R[974][6];				r_cell_reg[926] = inform_R[911][6];				r_cell_reg[927] = inform_R[975][6];				r_cell_reg[928] = inform_R[912][6];				r_cell_reg[929] = inform_R[976][6];				r_cell_reg[930] = inform_R[913][6];				r_cell_reg[931] = inform_R[977][6];				r_cell_reg[932] = inform_R[914][6];				r_cell_reg[933] = inform_R[978][6];				r_cell_reg[934] = inform_R[915][6];				r_cell_reg[935] = inform_R[979][6];				r_cell_reg[936] = inform_R[916][6];				r_cell_reg[937] = inform_R[980][6];				r_cell_reg[938] = inform_R[917][6];				r_cell_reg[939] = inform_R[981][6];				r_cell_reg[940] = inform_R[918][6];				r_cell_reg[941] = inform_R[982][6];				r_cell_reg[942] = inform_R[919][6];				r_cell_reg[943] = inform_R[983][6];				r_cell_reg[944] = inform_R[920][6];				r_cell_reg[945] = inform_R[984][6];				r_cell_reg[946] = inform_R[921][6];				r_cell_reg[947] = inform_R[985][6];				r_cell_reg[948] = inform_R[922][6];				r_cell_reg[949] = inform_R[986][6];				r_cell_reg[950] = inform_R[923][6];				r_cell_reg[951] = inform_R[987][6];				r_cell_reg[952] = inform_R[924][6];				r_cell_reg[953] = inform_R[988][6];				r_cell_reg[954] = inform_R[925][6];				r_cell_reg[955] = inform_R[989][6];				r_cell_reg[956] = inform_R[926][6];				r_cell_reg[957] = inform_R[990][6];				r_cell_reg[958] = inform_R[927][6];				r_cell_reg[959] = inform_R[991][6];				r_cell_reg[960] = inform_R[928][6];				r_cell_reg[961] = inform_R[992][6];				r_cell_reg[962] = inform_R[929][6];				r_cell_reg[963] = inform_R[993][6];				r_cell_reg[964] = inform_R[930][6];				r_cell_reg[965] = inform_R[994][6];				r_cell_reg[966] = inform_R[931][6];				r_cell_reg[967] = inform_R[995][6];				r_cell_reg[968] = inform_R[932][6];				r_cell_reg[969] = inform_R[996][6];				r_cell_reg[970] = inform_R[933][6];				r_cell_reg[971] = inform_R[997][6];				r_cell_reg[972] = inform_R[934][6];				r_cell_reg[973] = inform_R[998][6];				r_cell_reg[974] = inform_R[935][6];				r_cell_reg[975] = inform_R[999][6];				r_cell_reg[976] = inform_R[936][6];				r_cell_reg[977] = inform_R[1000][6];				r_cell_reg[978] = inform_R[937][6];				r_cell_reg[979] = inform_R[1001][6];				r_cell_reg[980] = inform_R[938][6];				r_cell_reg[981] = inform_R[1002][6];				r_cell_reg[982] = inform_R[939][6];				r_cell_reg[983] = inform_R[1003][6];				r_cell_reg[984] = inform_R[940][6];				r_cell_reg[985] = inform_R[1004][6];				r_cell_reg[986] = inform_R[941][6];				r_cell_reg[987] = inform_R[1005][6];				r_cell_reg[988] = inform_R[942][6];				r_cell_reg[989] = inform_R[1006][6];				r_cell_reg[990] = inform_R[943][6];				r_cell_reg[991] = inform_R[1007][6];				r_cell_reg[992] = inform_R[944][6];				r_cell_reg[993] = inform_R[1008][6];				r_cell_reg[994] = inform_R[945][6];				r_cell_reg[995] = inform_R[1009][6];				r_cell_reg[996] = inform_R[946][6];				r_cell_reg[997] = inform_R[1010][6];				r_cell_reg[998] = inform_R[947][6];				r_cell_reg[999] = inform_R[1011][6];				r_cell_reg[1000] = inform_R[948][6];				r_cell_reg[1001] = inform_R[1012][6];				r_cell_reg[1002] = inform_R[949][6];				r_cell_reg[1003] = inform_R[1013][6];				r_cell_reg[1004] = inform_R[950][6];				r_cell_reg[1005] = inform_R[1014][6];				r_cell_reg[1006] = inform_R[951][6];				r_cell_reg[1007] = inform_R[1015][6];				r_cell_reg[1008] = inform_R[952][6];				r_cell_reg[1009] = inform_R[1016][6];				r_cell_reg[1010] = inform_R[953][6];				r_cell_reg[1011] = inform_R[1017][6];				r_cell_reg[1012] = inform_R[954][6];				r_cell_reg[1013] = inform_R[1018][6];				r_cell_reg[1014] = inform_R[955][6];				r_cell_reg[1015] = inform_R[1019][6];				r_cell_reg[1016] = inform_R[956][6];				r_cell_reg[1017] = inform_R[1020][6];				r_cell_reg[1018] = inform_R[957][6];				r_cell_reg[1019] = inform_R[1021][6];				r_cell_reg[1020] = inform_R[958][6];				r_cell_reg[1021] = inform_R[1022][6];				r_cell_reg[1022] = inform_R[959][6];				r_cell_reg[1023] = inform_R[1023][6];				l_cell_reg[0] = inform_L[0][7];				l_cell_reg[1] = inform_L[64][7];				l_cell_reg[2] = inform_L[1][7];				l_cell_reg[3] = inform_L[65][7];				l_cell_reg[4] = inform_L[2][7];				l_cell_reg[5] = inform_L[66][7];				l_cell_reg[6] = inform_L[3][7];				l_cell_reg[7] = inform_L[67][7];				l_cell_reg[8] = inform_L[4][7];				l_cell_reg[9] = inform_L[68][7];				l_cell_reg[10] = inform_L[5][7];				l_cell_reg[11] = inform_L[69][7];				l_cell_reg[12] = inform_L[6][7];				l_cell_reg[13] = inform_L[70][7];				l_cell_reg[14] = inform_L[7][7];				l_cell_reg[15] = inform_L[71][7];				l_cell_reg[16] = inform_L[8][7];				l_cell_reg[17] = inform_L[72][7];				l_cell_reg[18] = inform_L[9][7];				l_cell_reg[19] = inform_L[73][7];				l_cell_reg[20] = inform_L[10][7];				l_cell_reg[21] = inform_L[74][7];				l_cell_reg[22] = inform_L[11][7];				l_cell_reg[23] = inform_L[75][7];				l_cell_reg[24] = inform_L[12][7];				l_cell_reg[25] = inform_L[76][7];				l_cell_reg[26] = inform_L[13][7];				l_cell_reg[27] = inform_L[77][7];				l_cell_reg[28] = inform_L[14][7];				l_cell_reg[29] = inform_L[78][7];				l_cell_reg[30] = inform_L[15][7];				l_cell_reg[31] = inform_L[79][7];				l_cell_reg[32] = inform_L[16][7];				l_cell_reg[33] = inform_L[80][7];				l_cell_reg[34] = inform_L[17][7];				l_cell_reg[35] = inform_L[81][7];				l_cell_reg[36] = inform_L[18][7];				l_cell_reg[37] = inform_L[82][7];				l_cell_reg[38] = inform_L[19][7];				l_cell_reg[39] = inform_L[83][7];				l_cell_reg[40] = inform_L[20][7];				l_cell_reg[41] = inform_L[84][7];				l_cell_reg[42] = inform_L[21][7];				l_cell_reg[43] = inform_L[85][7];				l_cell_reg[44] = inform_L[22][7];				l_cell_reg[45] = inform_L[86][7];				l_cell_reg[46] = inform_L[23][7];				l_cell_reg[47] = inform_L[87][7];				l_cell_reg[48] = inform_L[24][7];				l_cell_reg[49] = inform_L[88][7];				l_cell_reg[50] = inform_L[25][7];				l_cell_reg[51] = inform_L[89][7];				l_cell_reg[52] = inform_L[26][7];				l_cell_reg[53] = inform_L[90][7];				l_cell_reg[54] = inform_L[27][7];				l_cell_reg[55] = inform_L[91][7];				l_cell_reg[56] = inform_L[28][7];				l_cell_reg[57] = inform_L[92][7];				l_cell_reg[58] = inform_L[29][7];				l_cell_reg[59] = inform_L[93][7];				l_cell_reg[60] = inform_L[30][7];				l_cell_reg[61] = inform_L[94][7];				l_cell_reg[62] = inform_L[31][7];				l_cell_reg[63] = inform_L[95][7];				l_cell_reg[64] = inform_L[32][7];				l_cell_reg[65] = inform_L[96][7];				l_cell_reg[66] = inform_L[33][7];				l_cell_reg[67] = inform_L[97][7];				l_cell_reg[68] = inform_L[34][7];				l_cell_reg[69] = inform_L[98][7];				l_cell_reg[70] = inform_L[35][7];				l_cell_reg[71] = inform_L[99][7];				l_cell_reg[72] = inform_L[36][7];				l_cell_reg[73] = inform_L[100][7];				l_cell_reg[74] = inform_L[37][7];				l_cell_reg[75] = inform_L[101][7];				l_cell_reg[76] = inform_L[38][7];				l_cell_reg[77] = inform_L[102][7];				l_cell_reg[78] = inform_L[39][7];				l_cell_reg[79] = inform_L[103][7];				l_cell_reg[80] = inform_L[40][7];				l_cell_reg[81] = inform_L[104][7];				l_cell_reg[82] = inform_L[41][7];				l_cell_reg[83] = inform_L[105][7];				l_cell_reg[84] = inform_L[42][7];				l_cell_reg[85] = inform_L[106][7];				l_cell_reg[86] = inform_L[43][7];				l_cell_reg[87] = inform_L[107][7];				l_cell_reg[88] = inform_L[44][7];				l_cell_reg[89] = inform_L[108][7];				l_cell_reg[90] = inform_L[45][7];				l_cell_reg[91] = inform_L[109][7];				l_cell_reg[92] = inform_L[46][7];				l_cell_reg[93] = inform_L[110][7];				l_cell_reg[94] = inform_L[47][7];				l_cell_reg[95] = inform_L[111][7];				l_cell_reg[96] = inform_L[48][7];				l_cell_reg[97] = inform_L[112][7];				l_cell_reg[98] = inform_L[49][7];				l_cell_reg[99] = inform_L[113][7];				l_cell_reg[100] = inform_L[50][7];				l_cell_reg[101] = inform_L[114][7];				l_cell_reg[102] = inform_L[51][7];				l_cell_reg[103] = inform_L[115][7];				l_cell_reg[104] = inform_L[52][7];				l_cell_reg[105] = inform_L[116][7];				l_cell_reg[106] = inform_L[53][7];				l_cell_reg[107] = inform_L[117][7];				l_cell_reg[108] = inform_L[54][7];				l_cell_reg[109] = inform_L[118][7];				l_cell_reg[110] = inform_L[55][7];				l_cell_reg[111] = inform_L[119][7];				l_cell_reg[112] = inform_L[56][7];				l_cell_reg[113] = inform_L[120][7];				l_cell_reg[114] = inform_L[57][7];				l_cell_reg[115] = inform_L[121][7];				l_cell_reg[116] = inform_L[58][7];				l_cell_reg[117] = inform_L[122][7];				l_cell_reg[118] = inform_L[59][7];				l_cell_reg[119] = inform_L[123][7];				l_cell_reg[120] = inform_L[60][7];				l_cell_reg[121] = inform_L[124][7];				l_cell_reg[122] = inform_L[61][7];				l_cell_reg[123] = inform_L[125][7];				l_cell_reg[124] = inform_L[62][7];				l_cell_reg[125] = inform_L[126][7];				l_cell_reg[126] = inform_L[63][7];				l_cell_reg[127] = inform_L[127][7];				l_cell_reg[128] = inform_L[128][7];				l_cell_reg[129] = inform_L[192][7];				l_cell_reg[130] = inform_L[129][7];				l_cell_reg[131] = inform_L[193][7];				l_cell_reg[132] = inform_L[130][7];				l_cell_reg[133] = inform_L[194][7];				l_cell_reg[134] = inform_L[131][7];				l_cell_reg[135] = inform_L[195][7];				l_cell_reg[136] = inform_L[132][7];				l_cell_reg[137] = inform_L[196][7];				l_cell_reg[138] = inform_L[133][7];				l_cell_reg[139] = inform_L[197][7];				l_cell_reg[140] = inform_L[134][7];				l_cell_reg[141] = inform_L[198][7];				l_cell_reg[142] = inform_L[135][7];				l_cell_reg[143] = inform_L[199][7];				l_cell_reg[144] = inform_L[136][7];				l_cell_reg[145] = inform_L[200][7];				l_cell_reg[146] = inform_L[137][7];				l_cell_reg[147] = inform_L[201][7];				l_cell_reg[148] = inform_L[138][7];				l_cell_reg[149] = inform_L[202][7];				l_cell_reg[150] = inform_L[139][7];				l_cell_reg[151] = inform_L[203][7];				l_cell_reg[152] = inform_L[140][7];				l_cell_reg[153] = inform_L[204][7];				l_cell_reg[154] = inform_L[141][7];				l_cell_reg[155] = inform_L[205][7];				l_cell_reg[156] = inform_L[142][7];				l_cell_reg[157] = inform_L[206][7];				l_cell_reg[158] = inform_L[143][7];				l_cell_reg[159] = inform_L[207][7];				l_cell_reg[160] = inform_L[144][7];				l_cell_reg[161] = inform_L[208][7];				l_cell_reg[162] = inform_L[145][7];				l_cell_reg[163] = inform_L[209][7];				l_cell_reg[164] = inform_L[146][7];				l_cell_reg[165] = inform_L[210][7];				l_cell_reg[166] = inform_L[147][7];				l_cell_reg[167] = inform_L[211][7];				l_cell_reg[168] = inform_L[148][7];				l_cell_reg[169] = inform_L[212][7];				l_cell_reg[170] = inform_L[149][7];				l_cell_reg[171] = inform_L[213][7];				l_cell_reg[172] = inform_L[150][7];				l_cell_reg[173] = inform_L[214][7];				l_cell_reg[174] = inform_L[151][7];				l_cell_reg[175] = inform_L[215][7];				l_cell_reg[176] = inform_L[152][7];				l_cell_reg[177] = inform_L[216][7];				l_cell_reg[178] = inform_L[153][7];				l_cell_reg[179] = inform_L[217][7];				l_cell_reg[180] = inform_L[154][7];				l_cell_reg[181] = inform_L[218][7];				l_cell_reg[182] = inform_L[155][7];				l_cell_reg[183] = inform_L[219][7];				l_cell_reg[184] = inform_L[156][7];				l_cell_reg[185] = inform_L[220][7];				l_cell_reg[186] = inform_L[157][7];				l_cell_reg[187] = inform_L[221][7];				l_cell_reg[188] = inform_L[158][7];				l_cell_reg[189] = inform_L[222][7];				l_cell_reg[190] = inform_L[159][7];				l_cell_reg[191] = inform_L[223][7];				l_cell_reg[192] = inform_L[160][7];				l_cell_reg[193] = inform_L[224][7];				l_cell_reg[194] = inform_L[161][7];				l_cell_reg[195] = inform_L[225][7];				l_cell_reg[196] = inform_L[162][7];				l_cell_reg[197] = inform_L[226][7];				l_cell_reg[198] = inform_L[163][7];				l_cell_reg[199] = inform_L[227][7];				l_cell_reg[200] = inform_L[164][7];				l_cell_reg[201] = inform_L[228][7];				l_cell_reg[202] = inform_L[165][7];				l_cell_reg[203] = inform_L[229][7];				l_cell_reg[204] = inform_L[166][7];				l_cell_reg[205] = inform_L[230][7];				l_cell_reg[206] = inform_L[167][7];				l_cell_reg[207] = inform_L[231][7];				l_cell_reg[208] = inform_L[168][7];				l_cell_reg[209] = inform_L[232][7];				l_cell_reg[210] = inform_L[169][7];				l_cell_reg[211] = inform_L[233][7];				l_cell_reg[212] = inform_L[170][7];				l_cell_reg[213] = inform_L[234][7];				l_cell_reg[214] = inform_L[171][7];				l_cell_reg[215] = inform_L[235][7];				l_cell_reg[216] = inform_L[172][7];				l_cell_reg[217] = inform_L[236][7];				l_cell_reg[218] = inform_L[173][7];				l_cell_reg[219] = inform_L[237][7];				l_cell_reg[220] = inform_L[174][7];				l_cell_reg[221] = inform_L[238][7];				l_cell_reg[222] = inform_L[175][7];				l_cell_reg[223] = inform_L[239][7];				l_cell_reg[224] = inform_L[176][7];				l_cell_reg[225] = inform_L[240][7];				l_cell_reg[226] = inform_L[177][7];				l_cell_reg[227] = inform_L[241][7];				l_cell_reg[228] = inform_L[178][7];				l_cell_reg[229] = inform_L[242][7];				l_cell_reg[230] = inform_L[179][7];				l_cell_reg[231] = inform_L[243][7];				l_cell_reg[232] = inform_L[180][7];				l_cell_reg[233] = inform_L[244][7];				l_cell_reg[234] = inform_L[181][7];				l_cell_reg[235] = inform_L[245][7];				l_cell_reg[236] = inform_L[182][7];				l_cell_reg[237] = inform_L[246][7];				l_cell_reg[238] = inform_L[183][7];				l_cell_reg[239] = inform_L[247][7];				l_cell_reg[240] = inform_L[184][7];				l_cell_reg[241] = inform_L[248][7];				l_cell_reg[242] = inform_L[185][7];				l_cell_reg[243] = inform_L[249][7];				l_cell_reg[244] = inform_L[186][7];				l_cell_reg[245] = inform_L[250][7];				l_cell_reg[246] = inform_L[187][7];				l_cell_reg[247] = inform_L[251][7];				l_cell_reg[248] = inform_L[188][7];				l_cell_reg[249] = inform_L[252][7];				l_cell_reg[250] = inform_L[189][7];				l_cell_reg[251] = inform_L[253][7];				l_cell_reg[252] = inform_L[190][7];				l_cell_reg[253] = inform_L[254][7];				l_cell_reg[254] = inform_L[191][7];				l_cell_reg[255] = inform_L[255][7];				l_cell_reg[256] = inform_L[256][7];				l_cell_reg[257] = inform_L[320][7];				l_cell_reg[258] = inform_L[257][7];				l_cell_reg[259] = inform_L[321][7];				l_cell_reg[260] = inform_L[258][7];				l_cell_reg[261] = inform_L[322][7];				l_cell_reg[262] = inform_L[259][7];				l_cell_reg[263] = inform_L[323][7];				l_cell_reg[264] = inform_L[260][7];				l_cell_reg[265] = inform_L[324][7];				l_cell_reg[266] = inform_L[261][7];				l_cell_reg[267] = inform_L[325][7];				l_cell_reg[268] = inform_L[262][7];				l_cell_reg[269] = inform_L[326][7];				l_cell_reg[270] = inform_L[263][7];				l_cell_reg[271] = inform_L[327][7];				l_cell_reg[272] = inform_L[264][7];				l_cell_reg[273] = inform_L[328][7];				l_cell_reg[274] = inform_L[265][7];				l_cell_reg[275] = inform_L[329][7];				l_cell_reg[276] = inform_L[266][7];				l_cell_reg[277] = inform_L[330][7];				l_cell_reg[278] = inform_L[267][7];				l_cell_reg[279] = inform_L[331][7];				l_cell_reg[280] = inform_L[268][7];				l_cell_reg[281] = inform_L[332][7];				l_cell_reg[282] = inform_L[269][7];				l_cell_reg[283] = inform_L[333][7];				l_cell_reg[284] = inform_L[270][7];				l_cell_reg[285] = inform_L[334][7];				l_cell_reg[286] = inform_L[271][7];				l_cell_reg[287] = inform_L[335][7];				l_cell_reg[288] = inform_L[272][7];				l_cell_reg[289] = inform_L[336][7];				l_cell_reg[290] = inform_L[273][7];				l_cell_reg[291] = inform_L[337][7];				l_cell_reg[292] = inform_L[274][7];				l_cell_reg[293] = inform_L[338][7];				l_cell_reg[294] = inform_L[275][7];				l_cell_reg[295] = inform_L[339][7];				l_cell_reg[296] = inform_L[276][7];				l_cell_reg[297] = inform_L[340][7];				l_cell_reg[298] = inform_L[277][7];				l_cell_reg[299] = inform_L[341][7];				l_cell_reg[300] = inform_L[278][7];				l_cell_reg[301] = inform_L[342][7];				l_cell_reg[302] = inform_L[279][7];				l_cell_reg[303] = inform_L[343][7];				l_cell_reg[304] = inform_L[280][7];				l_cell_reg[305] = inform_L[344][7];				l_cell_reg[306] = inform_L[281][7];				l_cell_reg[307] = inform_L[345][7];				l_cell_reg[308] = inform_L[282][7];				l_cell_reg[309] = inform_L[346][7];				l_cell_reg[310] = inform_L[283][7];				l_cell_reg[311] = inform_L[347][7];				l_cell_reg[312] = inform_L[284][7];				l_cell_reg[313] = inform_L[348][7];				l_cell_reg[314] = inform_L[285][7];				l_cell_reg[315] = inform_L[349][7];				l_cell_reg[316] = inform_L[286][7];				l_cell_reg[317] = inform_L[350][7];				l_cell_reg[318] = inform_L[287][7];				l_cell_reg[319] = inform_L[351][7];				l_cell_reg[320] = inform_L[288][7];				l_cell_reg[321] = inform_L[352][7];				l_cell_reg[322] = inform_L[289][7];				l_cell_reg[323] = inform_L[353][7];				l_cell_reg[324] = inform_L[290][7];				l_cell_reg[325] = inform_L[354][7];				l_cell_reg[326] = inform_L[291][7];				l_cell_reg[327] = inform_L[355][7];				l_cell_reg[328] = inform_L[292][7];				l_cell_reg[329] = inform_L[356][7];				l_cell_reg[330] = inform_L[293][7];				l_cell_reg[331] = inform_L[357][7];				l_cell_reg[332] = inform_L[294][7];				l_cell_reg[333] = inform_L[358][7];				l_cell_reg[334] = inform_L[295][7];				l_cell_reg[335] = inform_L[359][7];				l_cell_reg[336] = inform_L[296][7];				l_cell_reg[337] = inform_L[360][7];				l_cell_reg[338] = inform_L[297][7];				l_cell_reg[339] = inform_L[361][7];				l_cell_reg[340] = inform_L[298][7];				l_cell_reg[341] = inform_L[362][7];				l_cell_reg[342] = inform_L[299][7];				l_cell_reg[343] = inform_L[363][7];				l_cell_reg[344] = inform_L[300][7];				l_cell_reg[345] = inform_L[364][7];				l_cell_reg[346] = inform_L[301][7];				l_cell_reg[347] = inform_L[365][7];				l_cell_reg[348] = inform_L[302][7];				l_cell_reg[349] = inform_L[366][7];				l_cell_reg[350] = inform_L[303][7];				l_cell_reg[351] = inform_L[367][7];				l_cell_reg[352] = inform_L[304][7];				l_cell_reg[353] = inform_L[368][7];				l_cell_reg[354] = inform_L[305][7];				l_cell_reg[355] = inform_L[369][7];				l_cell_reg[356] = inform_L[306][7];				l_cell_reg[357] = inform_L[370][7];				l_cell_reg[358] = inform_L[307][7];				l_cell_reg[359] = inform_L[371][7];				l_cell_reg[360] = inform_L[308][7];				l_cell_reg[361] = inform_L[372][7];				l_cell_reg[362] = inform_L[309][7];				l_cell_reg[363] = inform_L[373][7];				l_cell_reg[364] = inform_L[310][7];				l_cell_reg[365] = inform_L[374][7];				l_cell_reg[366] = inform_L[311][7];				l_cell_reg[367] = inform_L[375][7];				l_cell_reg[368] = inform_L[312][7];				l_cell_reg[369] = inform_L[376][7];				l_cell_reg[370] = inform_L[313][7];				l_cell_reg[371] = inform_L[377][7];				l_cell_reg[372] = inform_L[314][7];				l_cell_reg[373] = inform_L[378][7];				l_cell_reg[374] = inform_L[315][7];				l_cell_reg[375] = inform_L[379][7];				l_cell_reg[376] = inform_L[316][7];				l_cell_reg[377] = inform_L[380][7];				l_cell_reg[378] = inform_L[317][7];				l_cell_reg[379] = inform_L[381][7];				l_cell_reg[380] = inform_L[318][7];				l_cell_reg[381] = inform_L[382][7];				l_cell_reg[382] = inform_L[319][7];				l_cell_reg[383] = inform_L[383][7];				l_cell_reg[384] = inform_L[384][7];				l_cell_reg[385] = inform_L[448][7];				l_cell_reg[386] = inform_L[385][7];				l_cell_reg[387] = inform_L[449][7];				l_cell_reg[388] = inform_L[386][7];				l_cell_reg[389] = inform_L[450][7];				l_cell_reg[390] = inform_L[387][7];				l_cell_reg[391] = inform_L[451][7];				l_cell_reg[392] = inform_L[388][7];				l_cell_reg[393] = inform_L[452][7];				l_cell_reg[394] = inform_L[389][7];				l_cell_reg[395] = inform_L[453][7];				l_cell_reg[396] = inform_L[390][7];				l_cell_reg[397] = inform_L[454][7];				l_cell_reg[398] = inform_L[391][7];				l_cell_reg[399] = inform_L[455][7];				l_cell_reg[400] = inform_L[392][7];				l_cell_reg[401] = inform_L[456][7];				l_cell_reg[402] = inform_L[393][7];				l_cell_reg[403] = inform_L[457][7];				l_cell_reg[404] = inform_L[394][7];				l_cell_reg[405] = inform_L[458][7];				l_cell_reg[406] = inform_L[395][7];				l_cell_reg[407] = inform_L[459][7];				l_cell_reg[408] = inform_L[396][7];				l_cell_reg[409] = inform_L[460][7];				l_cell_reg[410] = inform_L[397][7];				l_cell_reg[411] = inform_L[461][7];				l_cell_reg[412] = inform_L[398][7];				l_cell_reg[413] = inform_L[462][7];				l_cell_reg[414] = inform_L[399][7];				l_cell_reg[415] = inform_L[463][7];				l_cell_reg[416] = inform_L[400][7];				l_cell_reg[417] = inform_L[464][7];				l_cell_reg[418] = inform_L[401][7];				l_cell_reg[419] = inform_L[465][7];				l_cell_reg[420] = inform_L[402][7];				l_cell_reg[421] = inform_L[466][7];				l_cell_reg[422] = inform_L[403][7];				l_cell_reg[423] = inform_L[467][7];				l_cell_reg[424] = inform_L[404][7];				l_cell_reg[425] = inform_L[468][7];				l_cell_reg[426] = inform_L[405][7];				l_cell_reg[427] = inform_L[469][7];				l_cell_reg[428] = inform_L[406][7];				l_cell_reg[429] = inform_L[470][7];				l_cell_reg[430] = inform_L[407][7];				l_cell_reg[431] = inform_L[471][7];				l_cell_reg[432] = inform_L[408][7];				l_cell_reg[433] = inform_L[472][7];				l_cell_reg[434] = inform_L[409][7];				l_cell_reg[435] = inform_L[473][7];				l_cell_reg[436] = inform_L[410][7];				l_cell_reg[437] = inform_L[474][7];				l_cell_reg[438] = inform_L[411][7];				l_cell_reg[439] = inform_L[475][7];				l_cell_reg[440] = inform_L[412][7];				l_cell_reg[441] = inform_L[476][7];				l_cell_reg[442] = inform_L[413][7];				l_cell_reg[443] = inform_L[477][7];				l_cell_reg[444] = inform_L[414][7];				l_cell_reg[445] = inform_L[478][7];				l_cell_reg[446] = inform_L[415][7];				l_cell_reg[447] = inform_L[479][7];				l_cell_reg[448] = inform_L[416][7];				l_cell_reg[449] = inform_L[480][7];				l_cell_reg[450] = inform_L[417][7];				l_cell_reg[451] = inform_L[481][7];				l_cell_reg[452] = inform_L[418][7];				l_cell_reg[453] = inform_L[482][7];				l_cell_reg[454] = inform_L[419][7];				l_cell_reg[455] = inform_L[483][7];				l_cell_reg[456] = inform_L[420][7];				l_cell_reg[457] = inform_L[484][7];				l_cell_reg[458] = inform_L[421][7];				l_cell_reg[459] = inform_L[485][7];				l_cell_reg[460] = inform_L[422][7];				l_cell_reg[461] = inform_L[486][7];				l_cell_reg[462] = inform_L[423][7];				l_cell_reg[463] = inform_L[487][7];				l_cell_reg[464] = inform_L[424][7];				l_cell_reg[465] = inform_L[488][7];				l_cell_reg[466] = inform_L[425][7];				l_cell_reg[467] = inform_L[489][7];				l_cell_reg[468] = inform_L[426][7];				l_cell_reg[469] = inform_L[490][7];				l_cell_reg[470] = inform_L[427][7];				l_cell_reg[471] = inform_L[491][7];				l_cell_reg[472] = inform_L[428][7];				l_cell_reg[473] = inform_L[492][7];				l_cell_reg[474] = inform_L[429][7];				l_cell_reg[475] = inform_L[493][7];				l_cell_reg[476] = inform_L[430][7];				l_cell_reg[477] = inform_L[494][7];				l_cell_reg[478] = inform_L[431][7];				l_cell_reg[479] = inform_L[495][7];				l_cell_reg[480] = inform_L[432][7];				l_cell_reg[481] = inform_L[496][7];				l_cell_reg[482] = inform_L[433][7];				l_cell_reg[483] = inform_L[497][7];				l_cell_reg[484] = inform_L[434][7];				l_cell_reg[485] = inform_L[498][7];				l_cell_reg[486] = inform_L[435][7];				l_cell_reg[487] = inform_L[499][7];				l_cell_reg[488] = inform_L[436][7];				l_cell_reg[489] = inform_L[500][7];				l_cell_reg[490] = inform_L[437][7];				l_cell_reg[491] = inform_L[501][7];				l_cell_reg[492] = inform_L[438][7];				l_cell_reg[493] = inform_L[502][7];				l_cell_reg[494] = inform_L[439][7];				l_cell_reg[495] = inform_L[503][7];				l_cell_reg[496] = inform_L[440][7];				l_cell_reg[497] = inform_L[504][7];				l_cell_reg[498] = inform_L[441][7];				l_cell_reg[499] = inform_L[505][7];				l_cell_reg[500] = inform_L[442][7];				l_cell_reg[501] = inform_L[506][7];				l_cell_reg[502] = inform_L[443][7];				l_cell_reg[503] = inform_L[507][7];				l_cell_reg[504] = inform_L[444][7];				l_cell_reg[505] = inform_L[508][7];				l_cell_reg[506] = inform_L[445][7];				l_cell_reg[507] = inform_L[509][7];				l_cell_reg[508] = inform_L[446][7];				l_cell_reg[509] = inform_L[510][7];				l_cell_reg[510] = inform_L[447][7];				l_cell_reg[511] = inform_L[511][7];				l_cell_reg[512] = inform_L[512][7];				l_cell_reg[513] = inform_L[576][7];				l_cell_reg[514] = inform_L[513][7];				l_cell_reg[515] = inform_L[577][7];				l_cell_reg[516] = inform_L[514][7];				l_cell_reg[517] = inform_L[578][7];				l_cell_reg[518] = inform_L[515][7];				l_cell_reg[519] = inform_L[579][7];				l_cell_reg[520] = inform_L[516][7];				l_cell_reg[521] = inform_L[580][7];				l_cell_reg[522] = inform_L[517][7];				l_cell_reg[523] = inform_L[581][7];				l_cell_reg[524] = inform_L[518][7];				l_cell_reg[525] = inform_L[582][7];				l_cell_reg[526] = inform_L[519][7];				l_cell_reg[527] = inform_L[583][7];				l_cell_reg[528] = inform_L[520][7];				l_cell_reg[529] = inform_L[584][7];				l_cell_reg[530] = inform_L[521][7];				l_cell_reg[531] = inform_L[585][7];				l_cell_reg[532] = inform_L[522][7];				l_cell_reg[533] = inform_L[586][7];				l_cell_reg[534] = inform_L[523][7];				l_cell_reg[535] = inform_L[587][7];				l_cell_reg[536] = inform_L[524][7];				l_cell_reg[537] = inform_L[588][7];				l_cell_reg[538] = inform_L[525][7];				l_cell_reg[539] = inform_L[589][7];				l_cell_reg[540] = inform_L[526][7];				l_cell_reg[541] = inform_L[590][7];				l_cell_reg[542] = inform_L[527][7];				l_cell_reg[543] = inform_L[591][7];				l_cell_reg[544] = inform_L[528][7];				l_cell_reg[545] = inform_L[592][7];				l_cell_reg[546] = inform_L[529][7];				l_cell_reg[547] = inform_L[593][7];				l_cell_reg[548] = inform_L[530][7];				l_cell_reg[549] = inform_L[594][7];				l_cell_reg[550] = inform_L[531][7];				l_cell_reg[551] = inform_L[595][7];				l_cell_reg[552] = inform_L[532][7];				l_cell_reg[553] = inform_L[596][7];				l_cell_reg[554] = inform_L[533][7];				l_cell_reg[555] = inform_L[597][7];				l_cell_reg[556] = inform_L[534][7];				l_cell_reg[557] = inform_L[598][7];				l_cell_reg[558] = inform_L[535][7];				l_cell_reg[559] = inform_L[599][7];				l_cell_reg[560] = inform_L[536][7];				l_cell_reg[561] = inform_L[600][7];				l_cell_reg[562] = inform_L[537][7];				l_cell_reg[563] = inform_L[601][7];				l_cell_reg[564] = inform_L[538][7];				l_cell_reg[565] = inform_L[602][7];				l_cell_reg[566] = inform_L[539][7];				l_cell_reg[567] = inform_L[603][7];				l_cell_reg[568] = inform_L[540][7];				l_cell_reg[569] = inform_L[604][7];				l_cell_reg[570] = inform_L[541][7];				l_cell_reg[571] = inform_L[605][7];				l_cell_reg[572] = inform_L[542][7];				l_cell_reg[573] = inform_L[606][7];				l_cell_reg[574] = inform_L[543][7];				l_cell_reg[575] = inform_L[607][7];				l_cell_reg[576] = inform_L[544][7];				l_cell_reg[577] = inform_L[608][7];				l_cell_reg[578] = inform_L[545][7];				l_cell_reg[579] = inform_L[609][7];				l_cell_reg[580] = inform_L[546][7];				l_cell_reg[581] = inform_L[610][7];				l_cell_reg[582] = inform_L[547][7];				l_cell_reg[583] = inform_L[611][7];				l_cell_reg[584] = inform_L[548][7];				l_cell_reg[585] = inform_L[612][7];				l_cell_reg[586] = inform_L[549][7];				l_cell_reg[587] = inform_L[613][7];				l_cell_reg[588] = inform_L[550][7];				l_cell_reg[589] = inform_L[614][7];				l_cell_reg[590] = inform_L[551][7];				l_cell_reg[591] = inform_L[615][7];				l_cell_reg[592] = inform_L[552][7];				l_cell_reg[593] = inform_L[616][7];				l_cell_reg[594] = inform_L[553][7];				l_cell_reg[595] = inform_L[617][7];				l_cell_reg[596] = inform_L[554][7];				l_cell_reg[597] = inform_L[618][7];				l_cell_reg[598] = inform_L[555][7];				l_cell_reg[599] = inform_L[619][7];				l_cell_reg[600] = inform_L[556][7];				l_cell_reg[601] = inform_L[620][7];				l_cell_reg[602] = inform_L[557][7];				l_cell_reg[603] = inform_L[621][7];				l_cell_reg[604] = inform_L[558][7];				l_cell_reg[605] = inform_L[622][7];				l_cell_reg[606] = inform_L[559][7];				l_cell_reg[607] = inform_L[623][7];				l_cell_reg[608] = inform_L[560][7];				l_cell_reg[609] = inform_L[624][7];				l_cell_reg[610] = inform_L[561][7];				l_cell_reg[611] = inform_L[625][7];				l_cell_reg[612] = inform_L[562][7];				l_cell_reg[613] = inform_L[626][7];				l_cell_reg[614] = inform_L[563][7];				l_cell_reg[615] = inform_L[627][7];				l_cell_reg[616] = inform_L[564][7];				l_cell_reg[617] = inform_L[628][7];				l_cell_reg[618] = inform_L[565][7];				l_cell_reg[619] = inform_L[629][7];				l_cell_reg[620] = inform_L[566][7];				l_cell_reg[621] = inform_L[630][7];				l_cell_reg[622] = inform_L[567][7];				l_cell_reg[623] = inform_L[631][7];				l_cell_reg[624] = inform_L[568][7];				l_cell_reg[625] = inform_L[632][7];				l_cell_reg[626] = inform_L[569][7];				l_cell_reg[627] = inform_L[633][7];				l_cell_reg[628] = inform_L[570][7];				l_cell_reg[629] = inform_L[634][7];				l_cell_reg[630] = inform_L[571][7];				l_cell_reg[631] = inform_L[635][7];				l_cell_reg[632] = inform_L[572][7];				l_cell_reg[633] = inform_L[636][7];				l_cell_reg[634] = inform_L[573][7];				l_cell_reg[635] = inform_L[637][7];				l_cell_reg[636] = inform_L[574][7];				l_cell_reg[637] = inform_L[638][7];				l_cell_reg[638] = inform_L[575][7];				l_cell_reg[639] = inform_L[639][7];				l_cell_reg[640] = inform_L[640][7];				l_cell_reg[641] = inform_L[704][7];				l_cell_reg[642] = inform_L[641][7];				l_cell_reg[643] = inform_L[705][7];				l_cell_reg[644] = inform_L[642][7];				l_cell_reg[645] = inform_L[706][7];				l_cell_reg[646] = inform_L[643][7];				l_cell_reg[647] = inform_L[707][7];				l_cell_reg[648] = inform_L[644][7];				l_cell_reg[649] = inform_L[708][7];				l_cell_reg[650] = inform_L[645][7];				l_cell_reg[651] = inform_L[709][7];				l_cell_reg[652] = inform_L[646][7];				l_cell_reg[653] = inform_L[710][7];				l_cell_reg[654] = inform_L[647][7];				l_cell_reg[655] = inform_L[711][7];				l_cell_reg[656] = inform_L[648][7];				l_cell_reg[657] = inform_L[712][7];				l_cell_reg[658] = inform_L[649][7];				l_cell_reg[659] = inform_L[713][7];				l_cell_reg[660] = inform_L[650][7];				l_cell_reg[661] = inform_L[714][7];				l_cell_reg[662] = inform_L[651][7];				l_cell_reg[663] = inform_L[715][7];				l_cell_reg[664] = inform_L[652][7];				l_cell_reg[665] = inform_L[716][7];				l_cell_reg[666] = inform_L[653][7];				l_cell_reg[667] = inform_L[717][7];				l_cell_reg[668] = inform_L[654][7];				l_cell_reg[669] = inform_L[718][7];				l_cell_reg[670] = inform_L[655][7];				l_cell_reg[671] = inform_L[719][7];				l_cell_reg[672] = inform_L[656][7];				l_cell_reg[673] = inform_L[720][7];				l_cell_reg[674] = inform_L[657][7];				l_cell_reg[675] = inform_L[721][7];				l_cell_reg[676] = inform_L[658][7];				l_cell_reg[677] = inform_L[722][7];				l_cell_reg[678] = inform_L[659][7];				l_cell_reg[679] = inform_L[723][7];				l_cell_reg[680] = inform_L[660][7];				l_cell_reg[681] = inform_L[724][7];				l_cell_reg[682] = inform_L[661][7];				l_cell_reg[683] = inform_L[725][7];				l_cell_reg[684] = inform_L[662][7];				l_cell_reg[685] = inform_L[726][7];				l_cell_reg[686] = inform_L[663][7];				l_cell_reg[687] = inform_L[727][7];				l_cell_reg[688] = inform_L[664][7];				l_cell_reg[689] = inform_L[728][7];				l_cell_reg[690] = inform_L[665][7];				l_cell_reg[691] = inform_L[729][7];				l_cell_reg[692] = inform_L[666][7];				l_cell_reg[693] = inform_L[730][7];				l_cell_reg[694] = inform_L[667][7];				l_cell_reg[695] = inform_L[731][7];				l_cell_reg[696] = inform_L[668][7];				l_cell_reg[697] = inform_L[732][7];				l_cell_reg[698] = inform_L[669][7];				l_cell_reg[699] = inform_L[733][7];				l_cell_reg[700] = inform_L[670][7];				l_cell_reg[701] = inform_L[734][7];				l_cell_reg[702] = inform_L[671][7];				l_cell_reg[703] = inform_L[735][7];				l_cell_reg[704] = inform_L[672][7];				l_cell_reg[705] = inform_L[736][7];				l_cell_reg[706] = inform_L[673][7];				l_cell_reg[707] = inform_L[737][7];				l_cell_reg[708] = inform_L[674][7];				l_cell_reg[709] = inform_L[738][7];				l_cell_reg[710] = inform_L[675][7];				l_cell_reg[711] = inform_L[739][7];				l_cell_reg[712] = inform_L[676][7];				l_cell_reg[713] = inform_L[740][7];				l_cell_reg[714] = inform_L[677][7];				l_cell_reg[715] = inform_L[741][7];				l_cell_reg[716] = inform_L[678][7];				l_cell_reg[717] = inform_L[742][7];				l_cell_reg[718] = inform_L[679][7];				l_cell_reg[719] = inform_L[743][7];				l_cell_reg[720] = inform_L[680][7];				l_cell_reg[721] = inform_L[744][7];				l_cell_reg[722] = inform_L[681][7];				l_cell_reg[723] = inform_L[745][7];				l_cell_reg[724] = inform_L[682][7];				l_cell_reg[725] = inform_L[746][7];				l_cell_reg[726] = inform_L[683][7];				l_cell_reg[727] = inform_L[747][7];				l_cell_reg[728] = inform_L[684][7];				l_cell_reg[729] = inform_L[748][7];				l_cell_reg[730] = inform_L[685][7];				l_cell_reg[731] = inform_L[749][7];				l_cell_reg[732] = inform_L[686][7];				l_cell_reg[733] = inform_L[750][7];				l_cell_reg[734] = inform_L[687][7];				l_cell_reg[735] = inform_L[751][7];				l_cell_reg[736] = inform_L[688][7];				l_cell_reg[737] = inform_L[752][7];				l_cell_reg[738] = inform_L[689][7];				l_cell_reg[739] = inform_L[753][7];				l_cell_reg[740] = inform_L[690][7];				l_cell_reg[741] = inform_L[754][7];				l_cell_reg[742] = inform_L[691][7];				l_cell_reg[743] = inform_L[755][7];				l_cell_reg[744] = inform_L[692][7];				l_cell_reg[745] = inform_L[756][7];				l_cell_reg[746] = inform_L[693][7];				l_cell_reg[747] = inform_L[757][7];				l_cell_reg[748] = inform_L[694][7];				l_cell_reg[749] = inform_L[758][7];				l_cell_reg[750] = inform_L[695][7];				l_cell_reg[751] = inform_L[759][7];				l_cell_reg[752] = inform_L[696][7];				l_cell_reg[753] = inform_L[760][7];				l_cell_reg[754] = inform_L[697][7];				l_cell_reg[755] = inform_L[761][7];				l_cell_reg[756] = inform_L[698][7];				l_cell_reg[757] = inform_L[762][7];				l_cell_reg[758] = inform_L[699][7];				l_cell_reg[759] = inform_L[763][7];				l_cell_reg[760] = inform_L[700][7];				l_cell_reg[761] = inform_L[764][7];				l_cell_reg[762] = inform_L[701][7];				l_cell_reg[763] = inform_L[765][7];				l_cell_reg[764] = inform_L[702][7];				l_cell_reg[765] = inform_L[766][7];				l_cell_reg[766] = inform_L[703][7];				l_cell_reg[767] = inform_L[767][7];				l_cell_reg[768] = inform_L[768][7];				l_cell_reg[769] = inform_L[832][7];				l_cell_reg[770] = inform_L[769][7];				l_cell_reg[771] = inform_L[833][7];				l_cell_reg[772] = inform_L[770][7];				l_cell_reg[773] = inform_L[834][7];				l_cell_reg[774] = inform_L[771][7];				l_cell_reg[775] = inform_L[835][7];				l_cell_reg[776] = inform_L[772][7];				l_cell_reg[777] = inform_L[836][7];				l_cell_reg[778] = inform_L[773][7];				l_cell_reg[779] = inform_L[837][7];				l_cell_reg[780] = inform_L[774][7];				l_cell_reg[781] = inform_L[838][7];				l_cell_reg[782] = inform_L[775][7];				l_cell_reg[783] = inform_L[839][7];				l_cell_reg[784] = inform_L[776][7];				l_cell_reg[785] = inform_L[840][7];				l_cell_reg[786] = inform_L[777][7];				l_cell_reg[787] = inform_L[841][7];				l_cell_reg[788] = inform_L[778][7];				l_cell_reg[789] = inform_L[842][7];				l_cell_reg[790] = inform_L[779][7];				l_cell_reg[791] = inform_L[843][7];				l_cell_reg[792] = inform_L[780][7];				l_cell_reg[793] = inform_L[844][7];				l_cell_reg[794] = inform_L[781][7];				l_cell_reg[795] = inform_L[845][7];				l_cell_reg[796] = inform_L[782][7];				l_cell_reg[797] = inform_L[846][7];				l_cell_reg[798] = inform_L[783][7];				l_cell_reg[799] = inform_L[847][7];				l_cell_reg[800] = inform_L[784][7];				l_cell_reg[801] = inform_L[848][7];				l_cell_reg[802] = inform_L[785][7];				l_cell_reg[803] = inform_L[849][7];				l_cell_reg[804] = inform_L[786][7];				l_cell_reg[805] = inform_L[850][7];				l_cell_reg[806] = inform_L[787][7];				l_cell_reg[807] = inform_L[851][7];				l_cell_reg[808] = inform_L[788][7];				l_cell_reg[809] = inform_L[852][7];				l_cell_reg[810] = inform_L[789][7];				l_cell_reg[811] = inform_L[853][7];				l_cell_reg[812] = inform_L[790][7];				l_cell_reg[813] = inform_L[854][7];				l_cell_reg[814] = inform_L[791][7];				l_cell_reg[815] = inform_L[855][7];				l_cell_reg[816] = inform_L[792][7];				l_cell_reg[817] = inform_L[856][7];				l_cell_reg[818] = inform_L[793][7];				l_cell_reg[819] = inform_L[857][7];				l_cell_reg[820] = inform_L[794][7];				l_cell_reg[821] = inform_L[858][7];				l_cell_reg[822] = inform_L[795][7];				l_cell_reg[823] = inform_L[859][7];				l_cell_reg[824] = inform_L[796][7];				l_cell_reg[825] = inform_L[860][7];				l_cell_reg[826] = inform_L[797][7];				l_cell_reg[827] = inform_L[861][7];				l_cell_reg[828] = inform_L[798][7];				l_cell_reg[829] = inform_L[862][7];				l_cell_reg[830] = inform_L[799][7];				l_cell_reg[831] = inform_L[863][7];				l_cell_reg[832] = inform_L[800][7];				l_cell_reg[833] = inform_L[864][7];				l_cell_reg[834] = inform_L[801][7];				l_cell_reg[835] = inform_L[865][7];				l_cell_reg[836] = inform_L[802][7];				l_cell_reg[837] = inform_L[866][7];				l_cell_reg[838] = inform_L[803][7];				l_cell_reg[839] = inform_L[867][7];				l_cell_reg[840] = inform_L[804][7];				l_cell_reg[841] = inform_L[868][7];				l_cell_reg[842] = inform_L[805][7];				l_cell_reg[843] = inform_L[869][7];				l_cell_reg[844] = inform_L[806][7];				l_cell_reg[845] = inform_L[870][7];				l_cell_reg[846] = inform_L[807][7];				l_cell_reg[847] = inform_L[871][7];				l_cell_reg[848] = inform_L[808][7];				l_cell_reg[849] = inform_L[872][7];				l_cell_reg[850] = inform_L[809][7];				l_cell_reg[851] = inform_L[873][7];				l_cell_reg[852] = inform_L[810][7];				l_cell_reg[853] = inform_L[874][7];				l_cell_reg[854] = inform_L[811][7];				l_cell_reg[855] = inform_L[875][7];				l_cell_reg[856] = inform_L[812][7];				l_cell_reg[857] = inform_L[876][7];				l_cell_reg[858] = inform_L[813][7];				l_cell_reg[859] = inform_L[877][7];				l_cell_reg[860] = inform_L[814][7];				l_cell_reg[861] = inform_L[878][7];				l_cell_reg[862] = inform_L[815][7];				l_cell_reg[863] = inform_L[879][7];				l_cell_reg[864] = inform_L[816][7];				l_cell_reg[865] = inform_L[880][7];				l_cell_reg[866] = inform_L[817][7];				l_cell_reg[867] = inform_L[881][7];				l_cell_reg[868] = inform_L[818][7];				l_cell_reg[869] = inform_L[882][7];				l_cell_reg[870] = inform_L[819][7];				l_cell_reg[871] = inform_L[883][7];				l_cell_reg[872] = inform_L[820][7];				l_cell_reg[873] = inform_L[884][7];				l_cell_reg[874] = inform_L[821][7];				l_cell_reg[875] = inform_L[885][7];				l_cell_reg[876] = inform_L[822][7];				l_cell_reg[877] = inform_L[886][7];				l_cell_reg[878] = inform_L[823][7];				l_cell_reg[879] = inform_L[887][7];				l_cell_reg[880] = inform_L[824][7];				l_cell_reg[881] = inform_L[888][7];				l_cell_reg[882] = inform_L[825][7];				l_cell_reg[883] = inform_L[889][7];				l_cell_reg[884] = inform_L[826][7];				l_cell_reg[885] = inform_L[890][7];				l_cell_reg[886] = inform_L[827][7];				l_cell_reg[887] = inform_L[891][7];				l_cell_reg[888] = inform_L[828][7];				l_cell_reg[889] = inform_L[892][7];				l_cell_reg[890] = inform_L[829][7];				l_cell_reg[891] = inform_L[893][7];				l_cell_reg[892] = inform_L[830][7];				l_cell_reg[893] = inform_L[894][7];				l_cell_reg[894] = inform_L[831][7];				l_cell_reg[895] = inform_L[895][7];				l_cell_reg[896] = inform_L[896][7];				l_cell_reg[897] = inform_L[960][7];				l_cell_reg[898] = inform_L[897][7];				l_cell_reg[899] = inform_L[961][7];				l_cell_reg[900] = inform_L[898][7];				l_cell_reg[901] = inform_L[962][7];				l_cell_reg[902] = inform_L[899][7];				l_cell_reg[903] = inform_L[963][7];				l_cell_reg[904] = inform_L[900][7];				l_cell_reg[905] = inform_L[964][7];				l_cell_reg[906] = inform_L[901][7];				l_cell_reg[907] = inform_L[965][7];				l_cell_reg[908] = inform_L[902][7];				l_cell_reg[909] = inform_L[966][7];				l_cell_reg[910] = inform_L[903][7];				l_cell_reg[911] = inform_L[967][7];				l_cell_reg[912] = inform_L[904][7];				l_cell_reg[913] = inform_L[968][7];				l_cell_reg[914] = inform_L[905][7];				l_cell_reg[915] = inform_L[969][7];				l_cell_reg[916] = inform_L[906][7];				l_cell_reg[917] = inform_L[970][7];				l_cell_reg[918] = inform_L[907][7];				l_cell_reg[919] = inform_L[971][7];				l_cell_reg[920] = inform_L[908][7];				l_cell_reg[921] = inform_L[972][7];				l_cell_reg[922] = inform_L[909][7];				l_cell_reg[923] = inform_L[973][7];				l_cell_reg[924] = inform_L[910][7];				l_cell_reg[925] = inform_L[974][7];				l_cell_reg[926] = inform_L[911][7];				l_cell_reg[927] = inform_L[975][7];				l_cell_reg[928] = inform_L[912][7];				l_cell_reg[929] = inform_L[976][7];				l_cell_reg[930] = inform_L[913][7];				l_cell_reg[931] = inform_L[977][7];				l_cell_reg[932] = inform_L[914][7];				l_cell_reg[933] = inform_L[978][7];				l_cell_reg[934] = inform_L[915][7];				l_cell_reg[935] = inform_L[979][7];				l_cell_reg[936] = inform_L[916][7];				l_cell_reg[937] = inform_L[980][7];				l_cell_reg[938] = inform_L[917][7];				l_cell_reg[939] = inform_L[981][7];				l_cell_reg[940] = inform_L[918][7];				l_cell_reg[941] = inform_L[982][7];				l_cell_reg[942] = inform_L[919][7];				l_cell_reg[943] = inform_L[983][7];				l_cell_reg[944] = inform_L[920][7];				l_cell_reg[945] = inform_L[984][7];				l_cell_reg[946] = inform_L[921][7];				l_cell_reg[947] = inform_L[985][7];				l_cell_reg[948] = inform_L[922][7];				l_cell_reg[949] = inform_L[986][7];				l_cell_reg[950] = inform_L[923][7];				l_cell_reg[951] = inform_L[987][7];				l_cell_reg[952] = inform_L[924][7];				l_cell_reg[953] = inform_L[988][7];				l_cell_reg[954] = inform_L[925][7];				l_cell_reg[955] = inform_L[989][7];				l_cell_reg[956] = inform_L[926][7];				l_cell_reg[957] = inform_L[990][7];				l_cell_reg[958] = inform_L[927][7];				l_cell_reg[959] = inform_L[991][7];				l_cell_reg[960] = inform_L[928][7];				l_cell_reg[961] = inform_L[992][7];				l_cell_reg[962] = inform_L[929][7];				l_cell_reg[963] = inform_L[993][7];				l_cell_reg[964] = inform_L[930][7];				l_cell_reg[965] = inform_L[994][7];				l_cell_reg[966] = inform_L[931][7];				l_cell_reg[967] = inform_L[995][7];				l_cell_reg[968] = inform_L[932][7];				l_cell_reg[969] = inform_L[996][7];				l_cell_reg[970] = inform_L[933][7];				l_cell_reg[971] = inform_L[997][7];				l_cell_reg[972] = inform_L[934][7];				l_cell_reg[973] = inform_L[998][7];				l_cell_reg[974] = inform_L[935][7];				l_cell_reg[975] = inform_L[999][7];				l_cell_reg[976] = inform_L[936][7];				l_cell_reg[977] = inform_L[1000][7];				l_cell_reg[978] = inform_L[937][7];				l_cell_reg[979] = inform_L[1001][7];				l_cell_reg[980] = inform_L[938][7];				l_cell_reg[981] = inform_L[1002][7];				l_cell_reg[982] = inform_L[939][7];				l_cell_reg[983] = inform_L[1003][7];				l_cell_reg[984] = inform_L[940][7];				l_cell_reg[985] = inform_L[1004][7];				l_cell_reg[986] = inform_L[941][7];				l_cell_reg[987] = inform_L[1005][7];				l_cell_reg[988] = inform_L[942][7];				l_cell_reg[989] = inform_L[1006][7];				l_cell_reg[990] = inform_L[943][7];				l_cell_reg[991] = inform_L[1007][7];				l_cell_reg[992] = inform_L[944][7];				l_cell_reg[993] = inform_L[1008][7];				l_cell_reg[994] = inform_L[945][7];				l_cell_reg[995] = inform_L[1009][7];				l_cell_reg[996] = inform_L[946][7];				l_cell_reg[997] = inform_L[1010][7];				l_cell_reg[998] = inform_L[947][7];				l_cell_reg[999] = inform_L[1011][7];				l_cell_reg[1000] = inform_L[948][7];				l_cell_reg[1001] = inform_L[1012][7];				l_cell_reg[1002] = inform_L[949][7];				l_cell_reg[1003] = inform_L[1013][7];				l_cell_reg[1004] = inform_L[950][7];				l_cell_reg[1005] = inform_L[1014][7];				l_cell_reg[1006] = inform_L[951][7];				l_cell_reg[1007] = inform_L[1015][7];				l_cell_reg[1008] = inform_L[952][7];				l_cell_reg[1009] = inform_L[1016][7];				l_cell_reg[1010] = inform_L[953][7];				l_cell_reg[1011] = inform_L[1017][7];				l_cell_reg[1012] = inform_L[954][7];				l_cell_reg[1013] = inform_L[1018][7];				l_cell_reg[1014] = inform_L[955][7];				l_cell_reg[1015] = inform_L[1019][7];				l_cell_reg[1016] = inform_L[956][7];				l_cell_reg[1017] = inform_L[1020][7];				l_cell_reg[1018] = inform_L[957][7];				l_cell_reg[1019] = inform_L[1021][7];				l_cell_reg[1020] = inform_L[958][7];				l_cell_reg[1021] = inform_L[1022][7];				l_cell_reg[1022] = inform_L[959][7];				l_cell_reg[1023] = inform_L[1023][7];			end
			8:			begin				r_cell_reg[0] = inform_R[0][7];				r_cell_reg[1] = inform_R[128][7];				r_cell_reg[2] = inform_R[1][7];				r_cell_reg[3] = inform_R[129][7];				r_cell_reg[4] = inform_R[2][7];				r_cell_reg[5] = inform_R[130][7];				r_cell_reg[6] = inform_R[3][7];				r_cell_reg[7] = inform_R[131][7];				r_cell_reg[8] = inform_R[4][7];				r_cell_reg[9] = inform_R[132][7];				r_cell_reg[10] = inform_R[5][7];				r_cell_reg[11] = inform_R[133][7];				r_cell_reg[12] = inform_R[6][7];				r_cell_reg[13] = inform_R[134][7];				r_cell_reg[14] = inform_R[7][7];				r_cell_reg[15] = inform_R[135][7];				r_cell_reg[16] = inform_R[8][7];				r_cell_reg[17] = inform_R[136][7];				r_cell_reg[18] = inform_R[9][7];				r_cell_reg[19] = inform_R[137][7];				r_cell_reg[20] = inform_R[10][7];				r_cell_reg[21] = inform_R[138][7];				r_cell_reg[22] = inform_R[11][7];				r_cell_reg[23] = inform_R[139][7];				r_cell_reg[24] = inform_R[12][7];				r_cell_reg[25] = inform_R[140][7];				r_cell_reg[26] = inform_R[13][7];				r_cell_reg[27] = inform_R[141][7];				r_cell_reg[28] = inform_R[14][7];				r_cell_reg[29] = inform_R[142][7];				r_cell_reg[30] = inform_R[15][7];				r_cell_reg[31] = inform_R[143][7];				r_cell_reg[32] = inform_R[16][7];				r_cell_reg[33] = inform_R[144][7];				r_cell_reg[34] = inform_R[17][7];				r_cell_reg[35] = inform_R[145][7];				r_cell_reg[36] = inform_R[18][7];				r_cell_reg[37] = inform_R[146][7];				r_cell_reg[38] = inform_R[19][7];				r_cell_reg[39] = inform_R[147][7];				r_cell_reg[40] = inform_R[20][7];				r_cell_reg[41] = inform_R[148][7];				r_cell_reg[42] = inform_R[21][7];				r_cell_reg[43] = inform_R[149][7];				r_cell_reg[44] = inform_R[22][7];				r_cell_reg[45] = inform_R[150][7];				r_cell_reg[46] = inform_R[23][7];				r_cell_reg[47] = inform_R[151][7];				r_cell_reg[48] = inform_R[24][7];				r_cell_reg[49] = inform_R[152][7];				r_cell_reg[50] = inform_R[25][7];				r_cell_reg[51] = inform_R[153][7];				r_cell_reg[52] = inform_R[26][7];				r_cell_reg[53] = inform_R[154][7];				r_cell_reg[54] = inform_R[27][7];				r_cell_reg[55] = inform_R[155][7];				r_cell_reg[56] = inform_R[28][7];				r_cell_reg[57] = inform_R[156][7];				r_cell_reg[58] = inform_R[29][7];				r_cell_reg[59] = inform_R[157][7];				r_cell_reg[60] = inform_R[30][7];				r_cell_reg[61] = inform_R[158][7];				r_cell_reg[62] = inform_R[31][7];				r_cell_reg[63] = inform_R[159][7];				r_cell_reg[64] = inform_R[32][7];				r_cell_reg[65] = inform_R[160][7];				r_cell_reg[66] = inform_R[33][7];				r_cell_reg[67] = inform_R[161][7];				r_cell_reg[68] = inform_R[34][7];				r_cell_reg[69] = inform_R[162][7];				r_cell_reg[70] = inform_R[35][7];				r_cell_reg[71] = inform_R[163][7];				r_cell_reg[72] = inform_R[36][7];				r_cell_reg[73] = inform_R[164][7];				r_cell_reg[74] = inform_R[37][7];				r_cell_reg[75] = inform_R[165][7];				r_cell_reg[76] = inform_R[38][7];				r_cell_reg[77] = inform_R[166][7];				r_cell_reg[78] = inform_R[39][7];				r_cell_reg[79] = inform_R[167][7];				r_cell_reg[80] = inform_R[40][7];				r_cell_reg[81] = inform_R[168][7];				r_cell_reg[82] = inform_R[41][7];				r_cell_reg[83] = inform_R[169][7];				r_cell_reg[84] = inform_R[42][7];				r_cell_reg[85] = inform_R[170][7];				r_cell_reg[86] = inform_R[43][7];				r_cell_reg[87] = inform_R[171][7];				r_cell_reg[88] = inform_R[44][7];				r_cell_reg[89] = inform_R[172][7];				r_cell_reg[90] = inform_R[45][7];				r_cell_reg[91] = inform_R[173][7];				r_cell_reg[92] = inform_R[46][7];				r_cell_reg[93] = inform_R[174][7];				r_cell_reg[94] = inform_R[47][7];				r_cell_reg[95] = inform_R[175][7];				r_cell_reg[96] = inform_R[48][7];				r_cell_reg[97] = inform_R[176][7];				r_cell_reg[98] = inform_R[49][7];				r_cell_reg[99] = inform_R[177][7];				r_cell_reg[100] = inform_R[50][7];				r_cell_reg[101] = inform_R[178][7];				r_cell_reg[102] = inform_R[51][7];				r_cell_reg[103] = inform_R[179][7];				r_cell_reg[104] = inform_R[52][7];				r_cell_reg[105] = inform_R[180][7];				r_cell_reg[106] = inform_R[53][7];				r_cell_reg[107] = inform_R[181][7];				r_cell_reg[108] = inform_R[54][7];				r_cell_reg[109] = inform_R[182][7];				r_cell_reg[110] = inform_R[55][7];				r_cell_reg[111] = inform_R[183][7];				r_cell_reg[112] = inform_R[56][7];				r_cell_reg[113] = inform_R[184][7];				r_cell_reg[114] = inform_R[57][7];				r_cell_reg[115] = inform_R[185][7];				r_cell_reg[116] = inform_R[58][7];				r_cell_reg[117] = inform_R[186][7];				r_cell_reg[118] = inform_R[59][7];				r_cell_reg[119] = inform_R[187][7];				r_cell_reg[120] = inform_R[60][7];				r_cell_reg[121] = inform_R[188][7];				r_cell_reg[122] = inform_R[61][7];				r_cell_reg[123] = inform_R[189][7];				r_cell_reg[124] = inform_R[62][7];				r_cell_reg[125] = inform_R[190][7];				r_cell_reg[126] = inform_R[63][7];				r_cell_reg[127] = inform_R[191][7];				r_cell_reg[128] = inform_R[64][7];				r_cell_reg[129] = inform_R[192][7];				r_cell_reg[130] = inform_R[65][7];				r_cell_reg[131] = inform_R[193][7];				r_cell_reg[132] = inform_R[66][7];				r_cell_reg[133] = inform_R[194][7];				r_cell_reg[134] = inform_R[67][7];				r_cell_reg[135] = inform_R[195][7];				r_cell_reg[136] = inform_R[68][7];				r_cell_reg[137] = inform_R[196][7];				r_cell_reg[138] = inform_R[69][7];				r_cell_reg[139] = inform_R[197][7];				r_cell_reg[140] = inform_R[70][7];				r_cell_reg[141] = inform_R[198][7];				r_cell_reg[142] = inform_R[71][7];				r_cell_reg[143] = inform_R[199][7];				r_cell_reg[144] = inform_R[72][7];				r_cell_reg[145] = inform_R[200][7];				r_cell_reg[146] = inform_R[73][7];				r_cell_reg[147] = inform_R[201][7];				r_cell_reg[148] = inform_R[74][7];				r_cell_reg[149] = inform_R[202][7];				r_cell_reg[150] = inform_R[75][7];				r_cell_reg[151] = inform_R[203][7];				r_cell_reg[152] = inform_R[76][7];				r_cell_reg[153] = inform_R[204][7];				r_cell_reg[154] = inform_R[77][7];				r_cell_reg[155] = inform_R[205][7];				r_cell_reg[156] = inform_R[78][7];				r_cell_reg[157] = inform_R[206][7];				r_cell_reg[158] = inform_R[79][7];				r_cell_reg[159] = inform_R[207][7];				r_cell_reg[160] = inform_R[80][7];				r_cell_reg[161] = inform_R[208][7];				r_cell_reg[162] = inform_R[81][7];				r_cell_reg[163] = inform_R[209][7];				r_cell_reg[164] = inform_R[82][7];				r_cell_reg[165] = inform_R[210][7];				r_cell_reg[166] = inform_R[83][7];				r_cell_reg[167] = inform_R[211][7];				r_cell_reg[168] = inform_R[84][7];				r_cell_reg[169] = inform_R[212][7];				r_cell_reg[170] = inform_R[85][7];				r_cell_reg[171] = inform_R[213][7];				r_cell_reg[172] = inform_R[86][7];				r_cell_reg[173] = inform_R[214][7];				r_cell_reg[174] = inform_R[87][7];				r_cell_reg[175] = inform_R[215][7];				r_cell_reg[176] = inform_R[88][7];				r_cell_reg[177] = inform_R[216][7];				r_cell_reg[178] = inform_R[89][7];				r_cell_reg[179] = inform_R[217][7];				r_cell_reg[180] = inform_R[90][7];				r_cell_reg[181] = inform_R[218][7];				r_cell_reg[182] = inform_R[91][7];				r_cell_reg[183] = inform_R[219][7];				r_cell_reg[184] = inform_R[92][7];				r_cell_reg[185] = inform_R[220][7];				r_cell_reg[186] = inform_R[93][7];				r_cell_reg[187] = inform_R[221][7];				r_cell_reg[188] = inform_R[94][7];				r_cell_reg[189] = inform_R[222][7];				r_cell_reg[190] = inform_R[95][7];				r_cell_reg[191] = inform_R[223][7];				r_cell_reg[192] = inform_R[96][7];				r_cell_reg[193] = inform_R[224][7];				r_cell_reg[194] = inform_R[97][7];				r_cell_reg[195] = inform_R[225][7];				r_cell_reg[196] = inform_R[98][7];				r_cell_reg[197] = inform_R[226][7];				r_cell_reg[198] = inform_R[99][7];				r_cell_reg[199] = inform_R[227][7];				r_cell_reg[200] = inform_R[100][7];				r_cell_reg[201] = inform_R[228][7];				r_cell_reg[202] = inform_R[101][7];				r_cell_reg[203] = inform_R[229][7];				r_cell_reg[204] = inform_R[102][7];				r_cell_reg[205] = inform_R[230][7];				r_cell_reg[206] = inform_R[103][7];				r_cell_reg[207] = inform_R[231][7];				r_cell_reg[208] = inform_R[104][7];				r_cell_reg[209] = inform_R[232][7];				r_cell_reg[210] = inform_R[105][7];				r_cell_reg[211] = inform_R[233][7];				r_cell_reg[212] = inform_R[106][7];				r_cell_reg[213] = inform_R[234][7];				r_cell_reg[214] = inform_R[107][7];				r_cell_reg[215] = inform_R[235][7];				r_cell_reg[216] = inform_R[108][7];				r_cell_reg[217] = inform_R[236][7];				r_cell_reg[218] = inform_R[109][7];				r_cell_reg[219] = inform_R[237][7];				r_cell_reg[220] = inform_R[110][7];				r_cell_reg[221] = inform_R[238][7];				r_cell_reg[222] = inform_R[111][7];				r_cell_reg[223] = inform_R[239][7];				r_cell_reg[224] = inform_R[112][7];				r_cell_reg[225] = inform_R[240][7];				r_cell_reg[226] = inform_R[113][7];				r_cell_reg[227] = inform_R[241][7];				r_cell_reg[228] = inform_R[114][7];				r_cell_reg[229] = inform_R[242][7];				r_cell_reg[230] = inform_R[115][7];				r_cell_reg[231] = inform_R[243][7];				r_cell_reg[232] = inform_R[116][7];				r_cell_reg[233] = inform_R[244][7];				r_cell_reg[234] = inform_R[117][7];				r_cell_reg[235] = inform_R[245][7];				r_cell_reg[236] = inform_R[118][7];				r_cell_reg[237] = inform_R[246][7];				r_cell_reg[238] = inform_R[119][7];				r_cell_reg[239] = inform_R[247][7];				r_cell_reg[240] = inform_R[120][7];				r_cell_reg[241] = inform_R[248][7];				r_cell_reg[242] = inform_R[121][7];				r_cell_reg[243] = inform_R[249][7];				r_cell_reg[244] = inform_R[122][7];				r_cell_reg[245] = inform_R[250][7];				r_cell_reg[246] = inform_R[123][7];				r_cell_reg[247] = inform_R[251][7];				r_cell_reg[248] = inform_R[124][7];				r_cell_reg[249] = inform_R[252][7];				r_cell_reg[250] = inform_R[125][7];				r_cell_reg[251] = inform_R[253][7];				r_cell_reg[252] = inform_R[126][7];				r_cell_reg[253] = inform_R[254][7];				r_cell_reg[254] = inform_R[127][7];				r_cell_reg[255] = inform_R[255][7];				r_cell_reg[256] = inform_R[256][7];				r_cell_reg[257] = inform_R[384][7];				r_cell_reg[258] = inform_R[257][7];				r_cell_reg[259] = inform_R[385][7];				r_cell_reg[260] = inform_R[258][7];				r_cell_reg[261] = inform_R[386][7];				r_cell_reg[262] = inform_R[259][7];				r_cell_reg[263] = inform_R[387][7];				r_cell_reg[264] = inform_R[260][7];				r_cell_reg[265] = inform_R[388][7];				r_cell_reg[266] = inform_R[261][7];				r_cell_reg[267] = inform_R[389][7];				r_cell_reg[268] = inform_R[262][7];				r_cell_reg[269] = inform_R[390][7];				r_cell_reg[270] = inform_R[263][7];				r_cell_reg[271] = inform_R[391][7];				r_cell_reg[272] = inform_R[264][7];				r_cell_reg[273] = inform_R[392][7];				r_cell_reg[274] = inform_R[265][7];				r_cell_reg[275] = inform_R[393][7];				r_cell_reg[276] = inform_R[266][7];				r_cell_reg[277] = inform_R[394][7];				r_cell_reg[278] = inform_R[267][7];				r_cell_reg[279] = inform_R[395][7];				r_cell_reg[280] = inform_R[268][7];				r_cell_reg[281] = inform_R[396][7];				r_cell_reg[282] = inform_R[269][7];				r_cell_reg[283] = inform_R[397][7];				r_cell_reg[284] = inform_R[270][7];				r_cell_reg[285] = inform_R[398][7];				r_cell_reg[286] = inform_R[271][7];				r_cell_reg[287] = inform_R[399][7];				r_cell_reg[288] = inform_R[272][7];				r_cell_reg[289] = inform_R[400][7];				r_cell_reg[290] = inform_R[273][7];				r_cell_reg[291] = inform_R[401][7];				r_cell_reg[292] = inform_R[274][7];				r_cell_reg[293] = inform_R[402][7];				r_cell_reg[294] = inform_R[275][7];				r_cell_reg[295] = inform_R[403][7];				r_cell_reg[296] = inform_R[276][7];				r_cell_reg[297] = inform_R[404][7];				r_cell_reg[298] = inform_R[277][7];				r_cell_reg[299] = inform_R[405][7];				r_cell_reg[300] = inform_R[278][7];				r_cell_reg[301] = inform_R[406][7];				r_cell_reg[302] = inform_R[279][7];				r_cell_reg[303] = inform_R[407][7];				r_cell_reg[304] = inform_R[280][7];				r_cell_reg[305] = inform_R[408][7];				r_cell_reg[306] = inform_R[281][7];				r_cell_reg[307] = inform_R[409][7];				r_cell_reg[308] = inform_R[282][7];				r_cell_reg[309] = inform_R[410][7];				r_cell_reg[310] = inform_R[283][7];				r_cell_reg[311] = inform_R[411][7];				r_cell_reg[312] = inform_R[284][7];				r_cell_reg[313] = inform_R[412][7];				r_cell_reg[314] = inform_R[285][7];				r_cell_reg[315] = inform_R[413][7];				r_cell_reg[316] = inform_R[286][7];				r_cell_reg[317] = inform_R[414][7];				r_cell_reg[318] = inform_R[287][7];				r_cell_reg[319] = inform_R[415][7];				r_cell_reg[320] = inform_R[288][7];				r_cell_reg[321] = inform_R[416][7];				r_cell_reg[322] = inform_R[289][7];				r_cell_reg[323] = inform_R[417][7];				r_cell_reg[324] = inform_R[290][7];				r_cell_reg[325] = inform_R[418][7];				r_cell_reg[326] = inform_R[291][7];				r_cell_reg[327] = inform_R[419][7];				r_cell_reg[328] = inform_R[292][7];				r_cell_reg[329] = inform_R[420][7];				r_cell_reg[330] = inform_R[293][7];				r_cell_reg[331] = inform_R[421][7];				r_cell_reg[332] = inform_R[294][7];				r_cell_reg[333] = inform_R[422][7];				r_cell_reg[334] = inform_R[295][7];				r_cell_reg[335] = inform_R[423][7];				r_cell_reg[336] = inform_R[296][7];				r_cell_reg[337] = inform_R[424][7];				r_cell_reg[338] = inform_R[297][7];				r_cell_reg[339] = inform_R[425][7];				r_cell_reg[340] = inform_R[298][7];				r_cell_reg[341] = inform_R[426][7];				r_cell_reg[342] = inform_R[299][7];				r_cell_reg[343] = inform_R[427][7];				r_cell_reg[344] = inform_R[300][7];				r_cell_reg[345] = inform_R[428][7];				r_cell_reg[346] = inform_R[301][7];				r_cell_reg[347] = inform_R[429][7];				r_cell_reg[348] = inform_R[302][7];				r_cell_reg[349] = inform_R[430][7];				r_cell_reg[350] = inform_R[303][7];				r_cell_reg[351] = inform_R[431][7];				r_cell_reg[352] = inform_R[304][7];				r_cell_reg[353] = inform_R[432][7];				r_cell_reg[354] = inform_R[305][7];				r_cell_reg[355] = inform_R[433][7];				r_cell_reg[356] = inform_R[306][7];				r_cell_reg[357] = inform_R[434][7];				r_cell_reg[358] = inform_R[307][7];				r_cell_reg[359] = inform_R[435][7];				r_cell_reg[360] = inform_R[308][7];				r_cell_reg[361] = inform_R[436][7];				r_cell_reg[362] = inform_R[309][7];				r_cell_reg[363] = inform_R[437][7];				r_cell_reg[364] = inform_R[310][7];				r_cell_reg[365] = inform_R[438][7];				r_cell_reg[366] = inform_R[311][7];				r_cell_reg[367] = inform_R[439][7];				r_cell_reg[368] = inform_R[312][7];				r_cell_reg[369] = inform_R[440][7];				r_cell_reg[370] = inform_R[313][7];				r_cell_reg[371] = inform_R[441][7];				r_cell_reg[372] = inform_R[314][7];				r_cell_reg[373] = inform_R[442][7];				r_cell_reg[374] = inform_R[315][7];				r_cell_reg[375] = inform_R[443][7];				r_cell_reg[376] = inform_R[316][7];				r_cell_reg[377] = inform_R[444][7];				r_cell_reg[378] = inform_R[317][7];				r_cell_reg[379] = inform_R[445][7];				r_cell_reg[380] = inform_R[318][7];				r_cell_reg[381] = inform_R[446][7];				r_cell_reg[382] = inform_R[319][7];				r_cell_reg[383] = inform_R[447][7];				r_cell_reg[384] = inform_R[320][7];				r_cell_reg[385] = inform_R[448][7];				r_cell_reg[386] = inform_R[321][7];				r_cell_reg[387] = inform_R[449][7];				r_cell_reg[388] = inform_R[322][7];				r_cell_reg[389] = inform_R[450][7];				r_cell_reg[390] = inform_R[323][7];				r_cell_reg[391] = inform_R[451][7];				r_cell_reg[392] = inform_R[324][7];				r_cell_reg[393] = inform_R[452][7];				r_cell_reg[394] = inform_R[325][7];				r_cell_reg[395] = inform_R[453][7];				r_cell_reg[396] = inform_R[326][7];				r_cell_reg[397] = inform_R[454][7];				r_cell_reg[398] = inform_R[327][7];				r_cell_reg[399] = inform_R[455][7];				r_cell_reg[400] = inform_R[328][7];				r_cell_reg[401] = inform_R[456][7];				r_cell_reg[402] = inform_R[329][7];				r_cell_reg[403] = inform_R[457][7];				r_cell_reg[404] = inform_R[330][7];				r_cell_reg[405] = inform_R[458][7];				r_cell_reg[406] = inform_R[331][7];				r_cell_reg[407] = inform_R[459][7];				r_cell_reg[408] = inform_R[332][7];				r_cell_reg[409] = inform_R[460][7];				r_cell_reg[410] = inform_R[333][7];				r_cell_reg[411] = inform_R[461][7];				r_cell_reg[412] = inform_R[334][7];				r_cell_reg[413] = inform_R[462][7];				r_cell_reg[414] = inform_R[335][7];				r_cell_reg[415] = inform_R[463][7];				r_cell_reg[416] = inform_R[336][7];				r_cell_reg[417] = inform_R[464][7];				r_cell_reg[418] = inform_R[337][7];				r_cell_reg[419] = inform_R[465][7];				r_cell_reg[420] = inform_R[338][7];				r_cell_reg[421] = inform_R[466][7];				r_cell_reg[422] = inform_R[339][7];				r_cell_reg[423] = inform_R[467][7];				r_cell_reg[424] = inform_R[340][7];				r_cell_reg[425] = inform_R[468][7];				r_cell_reg[426] = inform_R[341][7];				r_cell_reg[427] = inform_R[469][7];				r_cell_reg[428] = inform_R[342][7];				r_cell_reg[429] = inform_R[470][7];				r_cell_reg[430] = inform_R[343][7];				r_cell_reg[431] = inform_R[471][7];				r_cell_reg[432] = inform_R[344][7];				r_cell_reg[433] = inform_R[472][7];				r_cell_reg[434] = inform_R[345][7];				r_cell_reg[435] = inform_R[473][7];				r_cell_reg[436] = inform_R[346][7];				r_cell_reg[437] = inform_R[474][7];				r_cell_reg[438] = inform_R[347][7];				r_cell_reg[439] = inform_R[475][7];				r_cell_reg[440] = inform_R[348][7];				r_cell_reg[441] = inform_R[476][7];				r_cell_reg[442] = inform_R[349][7];				r_cell_reg[443] = inform_R[477][7];				r_cell_reg[444] = inform_R[350][7];				r_cell_reg[445] = inform_R[478][7];				r_cell_reg[446] = inform_R[351][7];				r_cell_reg[447] = inform_R[479][7];				r_cell_reg[448] = inform_R[352][7];				r_cell_reg[449] = inform_R[480][7];				r_cell_reg[450] = inform_R[353][7];				r_cell_reg[451] = inform_R[481][7];				r_cell_reg[452] = inform_R[354][7];				r_cell_reg[453] = inform_R[482][7];				r_cell_reg[454] = inform_R[355][7];				r_cell_reg[455] = inform_R[483][7];				r_cell_reg[456] = inform_R[356][7];				r_cell_reg[457] = inform_R[484][7];				r_cell_reg[458] = inform_R[357][7];				r_cell_reg[459] = inform_R[485][7];				r_cell_reg[460] = inform_R[358][7];				r_cell_reg[461] = inform_R[486][7];				r_cell_reg[462] = inform_R[359][7];				r_cell_reg[463] = inform_R[487][7];				r_cell_reg[464] = inform_R[360][7];				r_cell_reg[465] = inform_R[488][7];				r_cell_reg[466] = inform_R[361][7];				r_cell_reg[467] = inform_R[489][7];				r_cell_reg[468] = inform_R[362][7];				r_cell_reg[469] = inform_R[490][7];				r_cell_reg[470] = inform_R[363][7];				r_cell_reg[471] = inform_R[491][7];				r_cell_reg[472] = inform_R[364][7];				r_cell_reg[473] = inform_R[492][7];				r_cell_reg[474] = inform_R[365][7];				r_cell_reg[475] = inform_R[493][7];				r_cell_reg[476] = inform_R[366][7];				r_cell_reg[477] = inform_R[494][7];				r_cell_reg[478] = inform_R[367][7];				r_cell_reg[479] = inform_R[495][7];				r_cell_reg[480] = inform_R[368][7];				r_cell_reg[481] = inform_R[496][7];				r_cell_reg[482] = inform_R[369][7];				r_cell_reg[483] = inform_R[497][7];				r_cell_reg[484] = inform_R[370][7];				r_cell_reg[485] = inform_R[498][7];				r_cell_reg[486] = inform_R[371][7];				r_cell_reg[487] = inform_R[499][7];				r_cell_reg[488] = inform_R[372][7];				r_cell_reg[489] = inform_R[500][7];				r_cell_reg[490] = inform_R[373][7];				r_cell_reg[491] = inform_R[501][7];				r_cell_reg[492] = inform_R[374][7];				r_cell_reg[493] = inform_R[502][7];				r_cell_reg[494] = inform_R[375][7];				r_cell_reg[495] = inform_R[503][7];				r_cell_reg[496] = inform_R[376][7];				r_cell_reg[497] = inform_R[504][7];				r_cell_reg[498] = inform_R[377][7];				r_cell_reg[499] = inform_R[505][7];				r_cell_reg[500] = inform_R[378][7];				r_cell_reg[501] = inform_R[506][7];				r_cell_reg[502] = inform_R[379][7];				r_cell_reg[503] = inform_R[507][7];				r_cell_reg[504] = inform_R[380][7];				r_cell_reg[505] = inform_R[508][7];				r_cell_reg[506] = inform_R[381][7];				r_cell_reg[507] = inform_R[509][7];				r_cell_reg[508] = inform_R[382][7];				r_cell_reg[509] = inform_R[510][7];				r_cell_reg[510] = inform_R[383][7];				r_cell_reg[511] = inform_R[511][7];				r_cell_reg[512] = inform_R[512][7];				r_cell_reg[513] = inform_R[640][7];				r_cell_reg[514] = inform_R[513][7];				r_cell_reg[515] = inform_R[641][7];				r_cell_reg[516] = inform_R[514][7];				r_cell_reg[517] = inform_R[642][7];				r_cell_reg[518] = inform_R[515][7];				r_cell_reg[519] = inform_R[643][7];				r_cell_reg[520] = inform_R[516][7];				r_cell_reg[521] = inform_R[644][7];				r_cell_reg[522] = inform_R[517][7];				r_cell_reg[523] = inform_R[645][7];				r_cell_reg[524] = inform_R[518][7];				r_cell_reg[525] = inform_R[646][7];				r_cell_reg[526] = inform_R[519][7];				r_cell_reg[527] = inform_R[647][7];				r_cell_reg[528] = inform_R[520][7];				r_cell_reg[529] = inform_R[648][7];				r_cell_reg[530] = inform_R[521][7];				r_cell_reg[531] = inform_R[649][7];				r_cell_reg[532] = inform_R[522][7];				r_cell_reg[533] = inform_R[650][7];				r_cell_reg[534] = inform_R[523][7];				r_cell_reg[535] = inform_R[651][7];				r_cell_reg[536] = inform_R[524][7];				r_cell_reg[537] = inform_R[652][7];				r_cell_reg[538] = inform_R[525][7];				r_cell_reg[539] = inform_R[653][7];				r_cell_reg[540] = inform_R[526][7];				r_cell_reg[541] = inform_R[654][7];				r_cell_reg[542] = inform_R[527][7];				r_cell_reg[543] = inform_R[655][7];				r_cell_reg[544] = inform_R[528][7];				r_cell_reg[545] = inform_R[656][7];				r_cell_reg[546] = inform_R[529][7];				r_cell_reg[547] = inform_R[657][7];				r_cell_reg[548] = inform_R[530][7];				r_cell_reg[549] = inform_R[658][7];				r_cell_reg[550] = inform_R[531][7];				r_cell_reg[551] = inform_R[659][7];				r_cell_reg[552] = inform_R[532][7];				r_cell_reg[553] = inform_R[660][7];				r_cell_reg[554] = inform_R[533][7];				r_cell_reg[555] = inform_R[661][7];				r_cell_reg[556] = inform_R[534][7];				r_cell_reg[557] = inform_R[662][7];				r_cell_reg[558] = inform_R[535][7];				r_cell_reg[559] = inform_R[663][7];				r_cell_reg[560] = inform_R[536][7];				r_cell_reg[561] = inform_R[664][7];				r_cell_reg[562] = inform_R[537][7];				r_cell_reg[563] = inform_R[665][7];				r_cell_reg[564] = inform_R[538][7];				r_cell_reg[565] = inform_R[666][7];				r_cell_reg[566] = inform_R[539][7];				r_cell_reg[567] = inform_R[667][7];				r_cell_reg[568] = inform_R[540][7];				r_cell_reg[569] = inform_R[668][7];				r_cell_reg[570] = inform_R[541][7];				r_cell_reg[571] = inform_R[669][7];				r_cell_reg[572] = inform_R[542][7];				r_cell_reg[573] = inform_R[670][7];				r_cell_reg[574] = inform_R[543][7];				r_cell_reg[575] = inform_R[671][7];				r_cell_reg[576] = inform_R[544][7];				r_cell_reg[577] = inform_R[672][7];				r_cell_reg[578] = inform_R[545][7];				r_cell_reg[579] = inform_R[673][7];				r_cell_reg[580] = inform_R[546][7];				r_cell_reg[581] = inform_R[674][7];				r_cell_reg[582] = inform_R[547][7];				r_cell_reg[583] = inform_R[675][7];				r_cell_reg[584] = inform_R[548][7];				r_cell_reg[585] = inform_R[676][7];				r_cell_reg[586] = inform_R[549][7];				r_cell_reg[587] = inform_R[677][7];				r_cell_reg[588] = inform_R[550][7];				r_cell_reg[589] = inform_R[678][7];				r_cell_reg[590] = inform_R[551][7];				r_cell_reg[591] = inform_R[679][7];				r_cell_reg[592] = inform_R[552][7];				r_cell_reg[593] = inform_R[680][7];				r_cell_reg[594] = inform_R[553][7];				r_cell_reg[595] = inform_R[681][7];				r_cell_reg[596] = inform_R[554][7];				r_cell_reg[597] = inform_R[682][7];				r_cell_reg[598] = inform_R[555][7];				r_cell_reg[599] = inform_R[683][7];				r_cell_reg[600] = inform_R[556][7];				r_cell_reg[601] = inform_R[684][7];				r_cell_reg[602] = inform_R[557][7];				r_cell_reg[603] = inform_R[685][7];				r_cell_reg[604] = inform_R[558][7];				r_cell_reg[605] = inform_R[686][7];				r_cell_reg[606] = inform_R[559][7];				r_cell_reg[607] = inform_R[687][7];				r_cell_reg[608] = inform_R[560][7];				r_cell_reg[609] = inform_R[688][7];				r_cell_reg[610] = inform_R[561][7];				r_cell_reg[611] = inform_R[689][7];				r_cell_reg[612] = inform_R[562][7];				r_cell_reg[613] = inform_R[690][7];				r_cell_reg[614] = inform_R[563][7];				r_cell_reg[615] = inform_R[691][7];				r_cell_reg[616] = inform_R[564][7];				r_cell_reg[617] = inform_R[692][7];				r_cell_reg[618] = inform_R[565][7];				r_cell_reg[619] = inform_R[693][7];				r_cell_reg[620] = inform_R[566][7];				r_cell_reg[621] = inform_R[694][7];				r_cell_reg[622] = inform_R[567][7];				r_cell_reg[623] = inform_R[695][7];				r_cell_reg[624] = inform_R[568][7];				r_cell_reg[625] = inform_R[696][7];				r_cell_reg[626] = inform_R[569][7];				r_cell_reg[627] = inform_R[697][7];				r_cell_reg[628] = inform_R[570][7];				r_cell_reg[629] = inform_R[698][7];				r_cell_reg[630] = inform_R[571][7];				r_cell_reg[631] = inform_R[699][7];				r_cell_reg[632] = inform_R[572][7];				r_cell_reg[633] = inform_R[700][7];				r_cell_reg[634] = inform_R[573][7];				r_cell_reg[635] = inform_R[701][7];				r_cell_reg[636] = inform_R[574][7];				r_cell_reg[637] = inform_R[702][7];				r_cell_reg[638] = inform_R[575][7];				r_cell_reg[639] = inform_R[703][7];				r_cell_reg[640] = inform_R[576][7];				r_cell_reg[641] = inform_R[704][7];				r_cell_reg[642] = inform_R[577][7];				r_cell_reg[643] = inform_R[705][7];				r_cell_reg[644] = inform_R[578][7];				r_cell_reg[645] = inform_R[706][7];				r_cell_reg[646] = inform_R[579][7];				r_cell_reg[647] = inform_R[707][7];				r_cell_reg[648] = inform_R[580][7];				r_cell_reg[649] = inform_R[708][7];				r_cell_reg[650] = inform_R[581][7];				r_cell_reg[651] = inform_R[709][7];				r_cell_reg[652] = inform_R[582][7];				r_cell_reg[653] = inform_R[710][7];				r_cell_reg[654] = inform_R[583][7];				r_cell_reg[655] = inform_R[711][7];				r_cell_reg[656] = inform_R[584][7];				r_cell_reg[657] = inform_R[712][7];				r_cell_reg[658] = inform_R[585][7];				r_cell_reg[659] = inform_R[713][7];				r_cell_reg[660] = inform_R[586][7];				r_cell_reg[661] = inform_R[714][7];				r_cell_reg[662] = inform_R[587][7];				r_cell_reg[663] = inform_R[715][7];				r_cell_reg[664] = inform_R[588][7];				r_cell_reg[665] = inform_R[716][7];				r_cell_reg[666] = inform_R[589][7];				r_cell_reg[667] = inform_R[717][7];				r_cell_reg[668] = inform_R[590][7];				r_cell_reg[669] = inform_R[718][7];				r_cell_reg[670] = inform_R[591][7];				r_cell_reg[671] = inform_R[719][7];				r_cell_reg[672] = inform_R[592][7];				r_cell_reg[673] = inform_R[720][7];				r_cell_reg[674] = inform_R[593][7];				r_cell_reg[675] = inform_R[721][7];				r_cell_reg[676] = inform_R[594][7];				r_cell_reg[677] = inform_R[722][7];				r_cell_reg[678] = inform_R[595][7];				r_cell_reg[679] = inform_R[723][7];				r_cell_reg[680] = inform_R[596][7];				r_cell_reg[681] = inform_R[724][7];				r_cell_reg[682] = inform_R[597][7];				r_cell_reg[683] = inform_R[725][7];				r_cell_reg[684] = inform_R[598][7];				r_cell_reg[685] = inform_R[726][7];				r_cell_reg[686] = inform_R[599][7];				r_cell_reg[687] = inform_R[727][7];				r_cell_reg[688] = inform_R[600][7];				r_cell_reg[689] = inform_R[728][7];				r_cell_reg[690] = inform_R[601][7];				r_cell_reg[691] = inform_R[729][7];				r_cell_reg[692] = inform_R[602][7];				r_cell_reg[693] = inform_R[730][7];				r_cell_reg[694] = inform_R[603][7];				r_cell_reg[695] = inform_R[731][7];				r_cell_reg[696] = inform_R[604][7];				r_cell_reg[697] = inform_R[732][7];				r_cell_reg[698] = inform_R[605][7];				r_cell_reg[699] = inform_R[733][7];				r_cell_reg[700] = inform_R[606][7];				r_cell_reg[701] = inform_R[734][7];				r_cell_reg[702] = inform_R[607][7];				r_cell_reg[703] = inform_R[735][7];				r_cell_reg[704] = inform_R[608][7];				r_cell_reg[705] = inform_R[736][7];				r_cell_reg[706] = inform_R[609][7];				r_cell_reg[707] = inform_R[737][7];				r_cell_reg[708] = inform_R[610][7];				r_cell_reg[709] = inform_R[738][7];				r_cell_reg[710] = inform_R[611][7];				r_cell_reg[711] = inform_R[739][7];				r_cell_reg[712] = inform_R[612][7];				r_cell_reg[713] = inform_R[740][7];				r_cell_reg[714] = inform_R[613][7];				r_cell_reg[715] = inform_R[741][7];				r_cell_reg[716] = inform_R[614][7];				r_cell_reg[717] = inform_R[742][7];				r_cell_reg[718] = inform_R[615][7];				r_cell_reg[719] = inform_R[743][7];				r_cell_reg[720] = inform_R[616][7];				r_cell_reg[721] = inform_R[744][7];				r_cell_reg[722] = inform_R[617][7];				r_cell_reg[723] = inform_R[745][7];				r_cell_reg[724] = inform_R[618][7];				r_cell_reg[725] = inform_R[746][7];				r_cell_reg[726] = inform_R[619][7];				r_cell_reg[727] = inform_R[747][7];				r_cell_reg[728] = inform_R[620][7];				r_cell_reg[729] = inform_R[748][7];				r_cell_reg[730] = inform_R[621][7];				r_cell_reg[731] = inform_R[749][7];				r_cell_reg[732] = inform_R[622][7];				r_cell_reg[733] = inform_R[750][7];				r_cell_reg[734] = inform_R[623][7];				r_cell_reg[735] = inform_R[751][7];				r_cell_reg[736] = inform_R[624][7];				r_cell_reg[737] = inform_R[752][7];				r_cell_reg[738] = inform_R[625][7];				r_cell_reg[739] = inform_R[753][7];				r_cell_reg[740] = inform_R[626][7];				r_cell_reg[741] = inform_R[754][7];				r_cell_reg[742] = inform_R[627][7];				r_cell_reg[743] = inform_R[755][7];				r_cell_reg[744] = inform_R[628][7];				r_cell_reg[745] = inform_R[756][7];				r_cell_reg[746] = inform_R[629][7];				r_cell_reg[747] = inform_R[757][7];				r_cell_reg[748] = inform_R[630][7];				r_cell_reg[749] = inform_R[758][7];				r_cell_reg[750] = inform_R[631][7];				r_cell_reg[751] = inform_R[759][7];				r_cell_reg[752] = inform_R[632][7];				r_cell_reg[753] = inform_R[760][7];				r_cell_reg[754] = inform_R[633][7];				r_cell_reg[755] = inform_R[761][7];				r_cell_reg[756] = inform_R[634][7];				r_cell_reg[757] = inform_R[762][7];				r_cell_reg[758] = inform_R[635][7];				r_cell_reg[759] = inform_R[763][7];				r_cell_reg[760] = inform_R[636][7];				r_cell_reg[761] = inform_R[764][7];				r_cell_reg[762] = inform_R[637][7];				r_cell_reg[763] = inform_R[765][7];				r_cell_reg[764] = inform_R[638][7];				r_cell_reg[765] = inform_R[766][7];				r_cell_reg[766] = inform_R[639][7];				r_cell_reg[767] = inform_R[767][7];				r_cell_reg[768] = inform_R[768][7];				r_cell_reg[769] = inform_R[896][7];				r_cell_reg[770] = inform_R[769][7];				r_cell_reg[771] = inform_R[897][7];				r_cell_reg[772] = inform_R[770][7];				r_cell_reg[773] = inform_R[898][7];				r_cell_reg[774] = inform_R[771][7];				r_cell_reg[775] = inform_R[899][7];				r_cell_reg[776] = inform_R[772][7];				r_cell_reg[777] = inform_R[900][7];				r_cell_reg[778] = inform_R[773][7];				r_cell_reg[779] = inform_R[901][7];				r_cell_reg[780] = inform_R[774][7];				r_cell_reg[781] = inform_R[902][7];				r_cell_reg[782] = inform_R[775][7];				r_cell_reg[783] = inform_R[903][7];				r_cell_reg[784] = inform_R[776][7];				r_cell_reg[785] = inform_R[904][7];				r_cell_reg[786] = inform_R[777][7];				r_cell_reg[787] = inform_R[905][7];				r_cell_reg[788] = inform_R[778][7];				r_cell_reg[789] = inform_R[906][7];				r_cell_reg[790] = inform_R[779][7];				r_cell_reg[791] = inform_R[907][7];				r_cell_reg[792] = inform_R[780][7];				r_cell_reg[793] = inform_R[908][7];				r_cell_reg[794] = inform_R[781][7];				r_cell_reg[795] = inform_R[909][7];				r_cell_reg[796] = inform_R[782][7];				r_cell_reg[797] = inform_R[910][7];				r_cell_reg[798] = inform_R[783][7];				r_cell_reg[799] = inform_R[911][7];				r_cell_reg[800] = inform_R[784][7];				r_cell_reg[801] = inform_R[912][7];				r_cell_reg[802] = inform_R[785][7];				r_cell_reg[803] = inform_R[913][7];				r_cell_reg[804] = inform_R[786][7];				r_cell_reg[805] = inform_R[914][7];				r_cell_reg[806] = inform_R[787][7];				r_cell_reg[807] = inform_R[915][7];				r_cell_reg[808] = inform_R[788][7];				r_cell_reg[809] = inform_R[916][7];				r_cell_reg[810] = inform_R[789][7];				r_cell_reg[811] = inform_R[917][7];				r_cell_reg[812] = inform_R[790][7];				r_cell_reg[813] = inform_R[918][7];				r_cell_reg[814] = inform_R[791][7];				r_cell_reg[815] = inform_R[919][7];				r_cell_reg[816] = inform_R[792][7];				r_cell_reg[817] = inform_R[920][7];				r_cell_reg[818] = inform_R[793][7];				r_cell_reg[819] = inform_R[921][7];				r_cell_reg[820] = inform_R[794][7];				r_cell_reg[821] = inform_R[922][7];				r_cell_reg[822] = inform_R[795][7];				r_cell_reg[823] = inform_R[923][7];				r_cell_reg[824] = inform_R[796][7];				r_cell_reg[825] = inform_R[924][7];				r_cell_reg[826] = inform_R[797][7];				r_cell_reg[827] = inform_R[925][7];				r_cell_reg[828] = inform_R[798][7];				r_cell_reg[829] = inform_R[926][7];				r_cell_reg[830] = inform_R[799][7];				r_cell_reg[831] = inform_R[927][7];				r_cell_reg[832] = inform_R[800][7];				r_cell_reg[833] = inform_R[928][7];				r_cell_reg[834] = inform_R[801][7];				r_cell_reg[835] = inform_R[929][7];				r_cell_reg[836] = inform_R[802][7];				r_cell_reg[837] = inform_R[930][7];				r_cell_reg[838] = inform_R[803][7];				r_cell_reg[839] = inform_R[931][7];				r_cell_reg[840] = inform_R[804][7];				r_cell_reg[841] = inform_R[932][7];				r_cell_reg[842] = inform_R[805][7];				r_cell_reg[843] = inform_R[933][7];				r_cell_reg[844] = inform_R[806][7];				r_cell_reg[845] = inform_R[934][7];				r_cell_reg[846] = inform_R[807][7];				r_cell_reg[847] = inform_R[935][7];				r_cell_reg[848] = inform_R[808][7];				r_cell_reg[849] = inform_R[936][7];				r_cell_reg[850] = inform_R[809][7];				r_cell_reg[851] = inform_R[937][7];				r_cell_reg[852] = inform_R[810][7];				r_cell_reg[853] = inform_R[938][7];				r_cell_reg[854] = inform_R[811][7];				r_cell_reg[855] = inform_R[939][7];				r_cell_reg[856] = inform_R[812][7];				r_cell_reg[857] = inform_R[940][7];				r_cell_reg[858] = inform_R[813][7];				r_cell_reg[859] = inform_R[941][7];				r_cell_reg[860] = inform_R[814][7];				r_cell_reg[861] = inform_R[942][7];				r_cell_reg[862] = inform_R[815][7];				r_cell_reg[863] = inform_R[943][7];				r_cell_reg[864] = inform_R[816][7];				r_cell_reg[865] = inform_R[944][7];				r_cell_reg[866] = inform_R[817][7];				r_cell_reg[867] = inform_R[945][7];				r_cell_reg[868] = inform_R[818][7];				r_cell_reg[869] = inform_R[946][7];				r_cell_reg[870] = inform_R[819][7];				r_cell_reg[871] = inform_R[947][7];				r_cell_reg[872] = inform_R[820][7];				r_cell_reg[873] = inform_R[948][7];				r_cell_reg[874] = inform_R[821][7];				r_cell_reg[875] = inform_R[949][7];				r_cell_reg[876] = inform_R[822][7];				r_cell_reg[877] = inform_R[950][7];				r_cell_reg[878] = inform_R[823][7];				r_cell_reg[879] = inform_R[951][7];				r_cell_reg[880] = inform_R[824][7];				r_cell_reg[881] = inform_R[952][7];				r_cell_reg[882] = inform_R[825][7];				r_cell_reg[883] = inform_R[953][7];				r_cell_reg[884] = inform_R[826][7];				r_cell_reg[885] = inform_R[954][7];				r_cell_reg[886] = inform_R[827][7];				r_cell_reg[887] = inform_R[955][7];				r_cell_reg[888] = inform_R[828][7];				r_cell_reg[889] = inform_R[956][7];				r_cell_reg[890] = inform_R[829][7];				r_cell_reg[891] = inform_R[957][7];				r_cell_reg[892] = inform_R[830][7];				r_cell_reg[893] = inform_R[958][7];				r_cell_reg[894] = inform_R[831][7];				r_cell_reg[895] = inform_R[959][7];				r_cell_reg[896] = inform_R[832][7];				r_cell_reg[897] = inform_R[960][7];				r_cell_reg[898] = inform_R[833][7];				r_cell_reg[899] = inform_R[961][7];				r_cell_reg[900] = inform_R[834][7];				r_cell_reg[901] = inform_R[962][7];				r_cell_reg[902] = inform_R[835][7];				r_cell_reg[903] = inform_R[963][7];				r_cell_reg[904] = inform_R[836][7];				r_cell_reg[905] = inform_R[964][7];				r_cell_reg[906] = inform_R[837][7];				r_cell_reg[907] = inform_R[965][7];				r_cell_reg[908] = inform_R[838][7];				r_cell_reg[909] = inform_R[966][7];				r_cell_reg[910] = inform_R[839][7];				r_cell_reg[911] = inform_R[967][7];				r_cell_reg[912] = inform_R[840][7];				r_cell_reg[913] = inform_R[968][7];				r_cell_reg[914] = inform_R[841][7];				r_cell_reg[915] = inform_R[969][7];				r_cell_reg[916] = inform_R[842][7];				r_cell_reg[917] = inform_R[970][7];				r_cell_reg[918] = inform_R[843][7];				r_cell_reg[919] = inform_R[971][7];				r_cell_reg[920] = inform_R[844][7];				r_cell_reg[921] = inform_R[972][7];				r_cell_reg[922] = inform_R[845][7];				r_cell_reg[923] = inform_R[973][7];				r_cell_reg[924] = inform_R[846][7];				r_cell_reg[925] = inform_R[974][7];				r_cell_reg[926] = inform_R[847][7];				r_cell_reg[927] = inform_R[975][7];				r_cell_reg[928] = inform_R[848][7];				r_cell_reg[929] = inform_R[976][7];				r_cell_reg[930] = inform_R[849][7];				r_cell_reg[931] = inform_R[977][7];				r_cell_reg[932] = inform_R[850][7];				r_cell_reg[933] = inform_R[978][7];				r_cell_reg[934] = inform_R[851][7];				r_cell_reg[935] = inform_R[979][7];				r_cell_reg[936] = inform_R[852][7];				r_cell_reg[937] = inform_R[980][7];				r_cell_reg[938] = inform_R[853][7];				r_cell_reg[939] = inform_R[981][7];				r_cell_reg[940] = inform_R[854][7];				r_cell_reg[941] = inform_R[982][7];				r_cell_reg[942] = inform_R[855][7];				r_cell_reg[943] = inform_R[983][7];				r_cell_reg[944] = inform_R[856][7];				r_cell_reg[945] = inform_R[984][7];				r_cell_reg[946] = inform_R[857][7];				r_cell_reg[947] = inform_R[985][7];				r_cell_reg[948] = inform_R[858][7];				r_cell_reg[949] = inform_R[986][7];				r_cell_reg[950] = inform_R[859][7];				r_cell_reg[951] = inform_R[987][7];				r_cell_reg[952] = inform_R[860][7];				r_cell_reg[953] = inform_R[988][7];				r_cell_reg[954] = inform_R[861][7];				r_cell_reg[955] = inform_R[989][7];				r_cell_reg[956] = inform_R[862][7];				r_cell_reg[957] = inform_R[990][7];				r_cell_reg[958] = inform_R[863][7];				r_cell_reg[959] = inform_R[991][7];				r_cell_reg[960] = inform_R[864][7];				r_cell_reg[961] = inform_R[992][7];				r_cell_reg[962] = inform_R[865][7];				r_cell_reg[963] = inform_R[993][7];				r_cell_reg[964] = inform_R[866][7];				r_cell_reg[965] = inform_R[994][7];				r_cell_reg[966] = inform_R[867][7];				r_cell_reg[967] = inform_R[995][7];				r_cell_reg[968] = inform_R[868][7];				r_cell_reg[969] = inform_R[996][7];				r_cell_reg[970] = inform_R[869][7];				r_cell_reg[971] = inform_R[997][7];				r_cell_reg[972] = inform_R[870][7];				r_cell_reg[973] = inform_R[998][7];				r_cell_reg[974] = inform_R[871][7];				r_cell_reg[975] = inform_R[999][7];				r_cell_reg[976] = inform_R[872][7];				r_cell_reg[977] = inform_R[1000][7];				r_cell_reg[978] = inform_R[873][7];				r_cell_reg[979] = inform_R[1001][7];				r_cell_reg[980] = inform_R[874][7];				r_cell_reg[981] = inform_R[1002][7];				r_cell_reg[982] = inform_R[875][7];				r_cell_reg[983] = inform_R[1003][7];				r_cell_reg[984] = inform_R[876][7];				r_cell_reg[985] = inform_R[1004][7];				r_cell_reg[986] = inform_R[877][7];				r_cell_reg[987] = inform_R[1005][7];				r_cell_reg[988] = inform_R[878][7];				r_cell_reg[989] = inform_R[1006][7];				r_cell_reg[990] = inform_R[879][7];				r_cell_reg[991] = inform_R[1007][7];				r_cell_reg[992] = inform_R[880][7];				r_cell_reg[993] = inform_R[1008][7];				r_cell_reg[994] = inform_R[881][7];				r_cell_reg[995] = inform_R[1009][7];				r_cell_reg[996] = inform_R[882][7];				r_cell_reg[997] = inform_R[1010][7];				r_cell_reg[998] = inform_R[883][7];				r_cell_reg[999] = inform_R[1011][7];				r_cell_reg[1000] = inform_R[884][7];				r_cell_reg[1001] = inform_R[1012][7];				r_cell_reg[1002] = inform_R[885][7];				r_cell_reg[1003] = inform_R[1013][7];				r_cell_reg[1004] = inform_R[886][7];				r_cell_reg[1005] = inform_R[1014][7];				r_cell_reg[1006] = inform_R[887][7];				r_cell_reg[1007] = inform_R[1015][7];				r_cell_reg[1008] = inform_R[888][7];				r_cell_reg[1009] = inform_R[1016][7];				r_cell_reg[1010] = inform_R[889][7];				r_cell_reg[1011] = inform_R[1017][7];				r_cell_reg[1012] = inform_R[890][7];				r_cell_reg[1013] = inform_R[1018][7];				r_cell_reg[1014] = inform_R[891][7];				r_cell_reg[1015] = inform_R[1019][7];				r_cell_reg[1016] = inform_R[892][7];				r_cell_reg[1017] = inform_R[1020][7];				r_cell_reg[1018] = inform_R[893][7];				r_cell_reg[1019] = inform_R[1021][7];				r_cell_reg[1020] = inform_R[894][7];				r_cell_reg[1021] = inform_R[1022][7];				r_cell_reg[1022] = inform_R[895][7];				r_cell_reg[1023] = inform_R[1023][7];				l_cell_reg[0] = inform_L[0][8];				l_cell_reg[1] = inform_L[128][8];				l_cell_reg[2] = inform_L[1][8];				l_cell_reg[3] = inform_L[129][8];				l_cell_reg[4] = inform_L[2][8];				l_cell_reg[5] = inform_L[130][8];				l_cell_reg[6] = inform_L[3][8];				l_cell_reg[7] = inform_L[131][8];				l_cell_reg[8] = inform_L[4][8];				l_cell_reg[9] = inform_L[132][8];				l_cell_reg[10] = inform_L[5][8];				l_cell_reg[11] = inform_L[133][8];				l_cell_reg[12] = inform_L[6][8];				l_cell_reg[13] = inform_L[134][8];				l_cell_reg[14] = inform_L[7][8];				l_cell_reg[15] = inform_L[135][8];				l_cell_reg[16] = inform_L[8][8];				l_cell_reg[17] = inform_L[136][8];				l_cell_reg[18] = inform_L[9][8];				l_cell_reg[19] = inform_L[137][8];				l_cell_reg[20] = inform_L[10][8];				l_cell_reg[21] = inform_L[138][8];				l_cell_reg[22] = inform_L[11][8];				l_cell_reg[23] = inform_L[139][8];				l_cell_reg[24] = inform_L[12][8];				l_cell_reg[25] = inform_L[140][8];				l_cell_reg[26] = inform_L[13][8];				l_cell_reg[27] = inform_L[141][8];				l_cell_reg[28] = inform_L[14][8];				l_cell_reg[29] = inform_L[142][8];				l_cell_reg[30] = inform_L[15][8];				l_cell_reg[31] = inform_L[143][8];				l_cell_reg[32] = inform_L[16][8];				l_cell_reg[33] = inform_L[144][8];				l_cell_reg[34] = inform_L[17][8];				l_cell_reg[35] = inform_L[145][8];				l_cell_reg[36] = inform_L[18][8];				l_cell_reg[37] = inform_L[146][8];				l_cell_reg[38] = inform_L[19][8];				l_cell_reg[39] = inform_L[147][8];				l_cell_reg[40] = inform_L[20][8];				l_cell_reg[41] = inform_L[148][8];				l_cell_reg[42] = inform_L[21][8];				l_cell_reg[43] = inform_L[149][8];				l_cell_reg[44] = inform_L[22][8];				l_cell_reg[45] = inform_L[150][8];				l_cell_reg[46] = inform_L[23][8];				l_cell_reg[47] = inform_L[151][8];				l_cell_reg[48] = inform_L[24][8];				l_cell_reg[49] = inform_L[152][8];				l_cell_reg[50] = inform_L[25][8];				l_cell_reg[51] = inform_L[153][8];				l_cell_reg[52] = inform_L[26][8];				l_cell_reg[53] = inform_L[154][8];				l_cell_reg[54] = inform_L[27][8];				l_cell_reg[55] = inform_L[155][8];				l_cell_reg[56] = inform_L[28][8];				l_cell_reg[57] = inform_L[156][8];				l_cell_reg[58] = inform_L[29][8];				l_cell_reg[59] = inform_L[157][8];				l_cell_reg[60] = inform_L[30][8];				l_cell_reg[61] = inform_L[158][8];				l_cell_reg[62] = inform_L[31][8];				l_cell_reg[63] = inform_L[159][8];				l_cell_reg[64] = inform_L[32][8];				l_cell_reg[65] = inform_L[160][8];				l_cell_reg[66] = inform_L[33][8];				l_cell_reg[67] = inform_L[161][8];				l_cell_reg[68] = inform_L[34][8];				l_cell_reg[69] = inform_L[162][8];				l_cell_reg[70] = inform_L[35][8];				l_cell_reg[71] = inform_L[163][8];				l_cell_reg[72] = inform_L[36][8];				l_cell_reg[73] = inform_L[164][8];				l_cell_reg[74] = inform_L[37][8];				l_cell_reg[75] = inform_L[165][8];				l_cell_reg[76] = inform_L[38][8];				l_cell_reg[77] = inform_L[166][8];				l_cell_reg[78] = inform_L[39][8];				l_cell_reg[79] = inform_L[167][8];				l_cell_reg[80] = inform_L[40][8];				l_cell_reg[81] = inform_L[168][8];				l_cell_reg[82] = inform_L[41][8];				l_cell_reg[83] = inform_L[169][8];				l_cell_reg[84] = inform_L[42][8];				l_cell_reg[85] = inform_L[170][8];				l_cell_reg[86] = inform_L[43][8];				l_cell_reg[87] = inform_L[171][8];				l_cell_reg[88] = inform_L[44][8];				l_cell_reg[89] = inform_L[172][8];				l_cell_reg[90] = inform_L[45][8];				l_cell_reg[91] = inform_L[173][8];				l_cell_reg[92] = inform_L[46][8];				l_cell_reg[93] = inform_L[174][8];				l_cell_reg[94] = inform_L[47][8];				l_cell_reg[95] = inform_L[175][8];				l_cell_reg[96] = inform_L[48][8];				l_cell_reg[97] = inform_L[176][8];				l_cell_reg[98] = inform_L[49][8];				l_cell_reg[99] = inform_L[177][8];				l_cell_reg[100] = inform_L[50][8];				l_cell_reg[101] = inform_L[178][8];				l_cell_reg[102] = inform_L[51][8];				l_cell_reg[103] = inform_L[179][8];				l_cell_reg[104] = inform_L[52][8];				l_cell_reg[105] = inform_L[180][8];				l_cell_reg[106] = inform_L[53][8];				l_cell_reg[107] = inform_L[181][8];				l_cell_reg[108] = inform_L[54][8];				l_cell_reg[109] = inform_L[182][8];				l_cell_reg[110] = inform_L[55][8];				l_cell_reg[111] = inform_L[183][8];				l_cell_reg[112] = inform_L[56][8];				l_cell_reg[113] = inform_L[184][8];				l_cell_reg[114] = inform_L[57][8];				l_cell_reg[115] = inform_L[185][8];				l_cell_reg[116] = inform_L[58][8];				l_cell_reg[117] = inform_L[186][8];				l_cell_reg[118] = inform_L[59][8];				l_cell_reg[119] = inform_L[187][8];				l_cell_reg[120] = inform_L[60][8];				l_cell_reg[121] = inform_L[188][8];				l_cell_reg[122] = inform_L[61][8];				l_cell_reg[123] = inform_L[189][8];				l_cell_reg[124] = inform_L[62][8];				l_cell_reg[125] = inform_L[190][8];				l_cell_reg[126] = inform_L[63][8];				l_cell_reg[127] = inform_L[191][8];				l_cell_reg[128] = inform_L[64][8];				l_cell_reg[129] = inform_L[192][8];				l_cell_reg[130] = inform_L[65][8];				l_cell_reg[131] = inform_L[193][8];				l_cell_reg[132] = inform_L[66][8];				l_cell_reg[133] = inform_L[194][8];				l_cell_reg[134] = inform_L[67][8];				l_cell_reg[135] = inform_L[195][8];				l_cell_reg[136] = inform_L[68][8];				l_cell_reg[137] = inform_L[196][8];				l_cell_reg[138] = inform_L[69][8];				l_cell_reg[139] = inform_L[197][8];				l_cell_reg[140] = inform_L[70][8];				l_cell_reg[141] = inform_L[198][8];				l_cell_reg[142] = inform_L[71][8];				l_cell_reg[143] = inform_L[199][8];				l_cell_reg[144] = inform_L[72][8];				l_cell_reg[145] = inform_L[200][8];				l_cell_reg[146] = inform_L[73][8];				l_cell_reg[147] = inform_L[201][8];				l_cell_reg[148] = inform_L[74][8];				l_cell_reg[149] = inform_L[202][8];				l_cell_reg[150] = inform_L[75][8];				l_cell_reg[151] = inform_L[203][8];				l_cell_reg[152] = inform_L[76][8];				l_cell_reg[153] = inform_L[204][8];				l_cell_reg[154] = inform_L[77][8];				l_cell_reg[155] = inform_L[205][8];				l_cell_reg[156] = inform_L[78][8];				l_cell_reg[157] = inform_L[206][8];				l_cell_reg[158] = inform_L[79][8];				l_cell_reg[159] = inform_L[207][8];				l_cell_reg[160] = inform_L[80][8];				l_cell_reg[161] = inform_L[208][8];				l_cell_reg[162] = inform_L[81][8];				l_cell_reg[163] = inform_L[209][8];				l_cell_reg[164] = inform_L[82][8];				l_cell_reg[165] = inform_L[210][8];				l_cell_reg[166] = inform_L[83][8];				l_cell_reg[167] = inform_L[211][8];				l_cell_reg[168] = inform_L[84][8];				l_cell_reg[169] = inform_L[212][8];				l_cell_reg[170] = inform_L[85][8];				l_cell_reg[171] = inform_L[213][8];				l_cell_reg[172] = inform_L[86][8];				l_cell_reg[173] = inform_L[214][8];				l_cell_reg[174] = inform_L[87][8];				l_cell_reg[175] = inform_L[215][8];				l_cell_reg[176] = inform_L[88][8];				l_cell_reg[177] = inform_L[216][8];				l_cell_reg[178] = inform_L[89][8];				l_cell_reg[179] = inform_L[217][8];				l_cell_reg[180] = inform_L[90][8];				l_cell_reg[181] = inform_L[218][8];				l_cell_reg[182] = inform_L[91][8];				l_cell_reg[183] = inform_L[219][8];				l_cell_reg[184] = inform_L[92][8];				l_cell_reg[185] = inform_L[220][8];				l_cell_reg[186] = inform_L[93][8];				l_cell_reg[187] = inform_L[221][8];				l_cell_reg[188] = inform_L[94][8];				l_cell_reg[189] = inform_L[222][8];				l_cell_reg[190] = inform_L[95][8];				l_cell_reg[191] = inform_L[223][8];				l_cell_reg[192] = inform_L[96][8];				l_cell_reg[193] = inform_L[224][8];				l_cell_reg[194] = inform_L[97][8];				l_cell_reg[195] = inform_L[225][8];				l_cell_reg[196] = inform_L[98][8];				l_cell_reg[197] = inform_L[226][8];				l_cell_reg[198] = inform_L[99][8];				l_cell_reg[199] = inform_L[227][8];				l_cell_reg[200] = inform_L[100][8];				l_cell_reg[201] = inform_L[228][8];				l_cell_reg[202] = inform_L[101][8];				l_cell_reg[203] = inform_L[229][8];				l_cell_reg[204] = inform_L[102][8];				l_cell_reg[205] = inform_L[230][8];				l_cell_reg[206] = inform_L[103][8];				l_cell_reg[207] = inform_L[231][8];				l_cell_reg[208] = inform_L[104][8];				l_cell_reg[209] = inform_L[232][8];				l_cell_reg[210] = inform_L[105][8];				l_cell_reg[211] = inform_L[233][8];				l_cell_reg[212] = inform_L[106][8];				l_cell_reg[213] = inform_L[234][8];				l_cell_reg[214] = inform_L[107][8];				l_cell_reg[215] = inform_L[235][8];				l_cell_reg[216] = inform_L[108][8];				l_cell_reg[217] = inform_L[236][8];				l_cell_reg[218] = inform_L[109][8];				l_cell_reg[219] = inform_L[237][8];				l_cell_reg[220] = inform_L[110][8];				l_cell_reg[221] = inform_L[238][8];				l_cell_reg[222] = inform_L[111][8];				l_cell_reg[223] = inform_L[239][8];				l_cell_reg[224] = inform_L[112][8];				l_cell_reg[225] = inform_L[240][8];				l_cell_reg[226] = inform_L[113][8];				l_cell_reg[227] = inform_L[241][8];				l_cell_reg[228] = inform_L[114][8];				l_cell_reg[229] = inform_L[242][8];				l_cell_reg[230] = inform_L[115][8];				l_cell_reg[231] = inform_L[243][8];				l_cell_reg[232] = inform_L[116][8];				l_cell_reg[233] = inform_L[244][8];				l_cell_reg[234] = inform_L[117][8];				l_cell_reg[235] = inform_L[245][8];				l_cell_reg[236] = inform_L[118][8];				l_cell_reg[237] = inform_L[246][8];				l_cell_reg[238] = inform_L[119][8];				l_cell_reg[239] = inform_L[247][8];				l_cell_reg[240] = inform_L[120][8];				l_cell_reg[241] = inform_L[248][8];				l_cell_reg[242] = inform_L[121][8];				l_cell_reg[243] = inform_L[249][8];				l_cell_reg[244] = inform_L[122][8];				l_cell_reg[245] = inform_L[250][8];				l_cell_reg[246] = inform_L[123][8];				l_cell_reg[247] = inform_L[251][8];				l_cell_reg[248] = inform_L[124][8];				l_cell_reg[249] = inform_L[252][8];				l_cell_reg[250] = inform_L[125][8];				l_cell_reg[251] = inform_L[253][8];				l_cell_reg[252] = inform_L[126][8];				l_cell_reg[253] = inform_L[254][8];				l_cell_reg[254] = inform_L[127][8];				l_cell_reg[255] = inform_L[255][8];				l_cell_reg[256] = inform_L[256][8];				l_cell_reg[257] = inform_L[384][8];				l_cell_reg[258] = inform_L[257][8];				l_cell_reg[259] = inform_L[385][8];				l_cell_reg[260] = inform_L[258][8];				l_cell_reg[261] = inform_L[386][8];				l_cell_reg[262] = inform_L[259][8];				l_cell_reg[263] = inform_L[387][8];				l_cell_reg[264] = inform_L[260][8];				l_cell_reg[265] = inform_L[388][8];				l_cell_reg[266] = inform_L[261][8];				l_cell_reg[267] = inform_L[389][8];				l_cell_reg[268] = inform_L[262][8];				l_cell_reg[269] = inform_L[390][8];				l_cell_reg[270] = inform_L[263][8];				l_cell_reg[271] = inform_L[391][8];				l_cell_reg[272] = inform_L[264][8];				l_cell_reg[273] = inform_L[392][8];				l_cell_reg[274] = inform_L[265][8];				l_cell_reg[275] = inform_L[393][8];				l_cell_reg[276] = inform_L[266][8];				l_cell_reg[277] = inform_L[394][8];				l_cell_reg[278] = inform_L[267][8];				l_cell_reg[279] = inform_L[395][8];				l_cell_reg[280] = inform_L[268][8];				l_cell_reg[281] = inform_L[396][8];				l_cell_reg[282] = inform_L[269][8];				l_cell_reg[283] = inform_L[397][8];				l_cell_reg[284] = inform_L[270][8];				l_cell_reg[285] = inform_L[398][8];				l_cell_reg[286] = inform_L[271][8];				l_cell_reg[287] = inform_L[399][8];				l_cell_reg[288] = inform_L[272][8];				l_cell_reg[289] = inform_L[400][8];				l_cell_reg[290] = inform_L[273][8];				l_cell_reg[291] = inform_L[401][8];				l_cell_reg[292] = inform_L[274][8];				l_cell_reg[293] = inform_L[402][8];				l_cell_reg[294] = inform_L[275][8];				l_cell_reg[295] = inform_L[403][8];				l_cell_reg[296] = inform_L[276][8];				l_cell_reg[297] = inform_L[404][8];				l_cell_reg[298] = inform_L[277][8];				l_cell_reg[299] = inform_L[405][8];				l_cell_reg[300] = inform_L[278][8];				l_cell_reg[301] = inform_L[406][8];				l_cell_reg[302] = inform_L[279][8];				l_cell_reg[303] = inform_L[407][8];				l_cell_reg[304] = inform_L[280][8];				l_cell_reg[305] = inform_L[408][8];				l_cell_reg[306] = inform_L[281][8];				l_cell_reg[307] = inform_L[409][8];				l_cell_reg[308] = inform_L[282][8];				l_cell_reg[309] = inform_L[410][8];				l_cell_reg[310] = inform_L[283][8];				l_cell_reg[311] = inform_L[411][8];				l_cell_reg[312] = inform_L[284][8];				l_cell_reg[313] = inform_L[412][8];				l_cell_reg[314] = inform_L[285][8];				l_cell_reg[315] = inform_L[413][8];				l_cell_reg[316] = inform_L[286][8];				l_cell_reg[317] = inform_L[414][8];				l_cell_reg[318] = inform_L[287][8];				l_cell_reg[319] = inform_L[415][8];				l_cell_reg[320] = inform_L[288][8];				l_cell_reg[321] = inform_L[416][8];				l_cell_reg[322] = inform_L[289][8];				l_cell_reg[323] = inform_L[417][8];				l_cell_reg[324] = inform_L[290][8];				l_cell_reg[325] = inform_L[418][8];				l_cell_reg[326] = inform_L[291][8];				l_cell_reg[327] = inform_L[419][8];				l_cell_reg[328] = inform_L[292][8];				l_cell_reg[329] = inform_L[420][8];				l_cell_reg[330] = inform_L[293][8];				l_cell_reg[331] = inform_L[421][8];				l_cell_reg[332] = inform_L[294][8];				l_cell_reg[333] = inform_L[422][8];				l_cell_reg[334] = inform_L[295][8];				l_cell_reg[335] = inform_L[423][8];				l_cell_reg[336] = inform_L[296][8];				l_cell_reg[337] = inform_L[424][8];				l_cell_reg[338] = inform_L[297][8];				l_cell_reg[339] = inform_L[425][8];				l_cell_reg[340] = inform_L[298][8];				l_cell_reg[341] = inform_L[426][8];				l_cell_reg[342] = inform_L[299][8];				l_cell_reg[343] = inform_L[427][8];				l_cell_reg[344] = inform_L[300][8];				l_cell_reg[345] = inform_L[428][8];				l_cell_reg[346] = inform_L[301][8];				l_cell_reg[347] = inform_L[429][8];				l_cell_reg[348] = inform_L[302][8];				l_cell_reg[349] = inform_L[430][8];				l_cell_reg[350] = inform_L[303][8];				l_cell_reg[351] = inform_L[431][8];				l_cell_reg[352] = inform_L[304][8];				l_cell_reg[353] = inform_L[432][8];				l_cell_reg[354] = inform_L[305][8];				l_cell_reg[355] = inform_L[433][8];				l_cell_reg[356] = inform_L[306][8];				l_cell_reg[357] = inform_L[434][8];				l_cell_reg[358] = inform_L[307][8];				l_cell_reg[359] = inform_L[435][8];				l_cell_reg[360] = inform_L[308][8];				l_cell_reg[361] = inform_L[436][8];				l_cell_reg[362] = inform_L[309][8];				l_cell_reg[363] = inform_L[437][8];				l_cell_reg[364] = inform_L[310][8];				l_cell_reg[365] = inform_L[438][8];				l_cell_reg[366] = inform_L[311][8];				l_cell_reg[367] = inform_L[439][8];				l_cell_reg[368] = inform_L[312][8];				l_cell_reg[369] = inform_L[440][8];				l_cell_reg[370] = inform_L[313][8];				l_cell_reg[371] = inform_L[441][8];				l_cell_reg[372] = inform_L[314][8];				l_cell_reg[373] = inform_L[442][8];				l_cell_reg[374] = inform_L[315][8];				l_cell_reg[375] = inform_L[443][8];				l_cell_reg[376] = inform_L[316][8];				l_cell_reg[377] = inform_L[444][8];				l_cell_reg[378] = inform_L[317][8];				l_cell_reg[379] = inform_L[445][8];				l_cell_reg[380] = inform_L[318][8];				l_cell_reg[381] = inform_L[446][8];				l_cell_reg[382] = inform_L[319][8];				l_cell_reg[383] = inform_L[447][8];				l_cell_reg[384] = inform_L[320][8];				l_cell_reg[385] = inform_L[448][8];				l_cell_reg[386] = inform_L[321][8];				l_cell_reg[387] = inform_L[449][8];				l_cell_reg[388] = inform_L[322][8];				l_cell_reg[389] = inform_L[450][8];				l_cell_reg[390] = inform_L[323][8];				l_cell_reg[391] = inform_L[451][8];				l_cell_reg[392] = inform_L[324][8];				l_cell_reg[393] = inform_L[452][8];				l_cell_reg[394] = inform_L[325][8];				l_cell_reg[395] = inform_L[453][8];				l_cell_reg[396] = inform_L[326][8];				l_cell_reg[397] = inform_L[454][8];				l_cell_reg[398] = inform_L[327][8];				l_cell_reg[399] = inform_L[455][8];				l_cell_reg[400] = inform_L[328][8];				l_cell_reg[401] = inform_L[456][8];				l_cell_reg[402] = inform_L[329][8];				l_cell_reg[403] = inform_L[457][8];				l_cell_reg[404] = inform_L[330][8];				l_cell_reg[405] = inform_L[458][8];				l_cell_reg[406] = inform_L[331][8];				l_cell_reg[407] = inform_L[459][8];				l_cell_reg[408] = inform_L[332][8];				l_cell_reg[409] = inform_L[460][8];				l_cell_reg[410] = inform_L[333][8];				l_cell_reg[411] = inform_L[461][8];				l_cell_reg[412] = inform_L[334][8];				l_cell_reg[413] = inform_L[462][8];				l_cell_reg[414] = inform_L[335][8];				l_cell_reg[415] = inform_L[463][8];				l_cell_reg[416] = inform_L[336][8];				l_cell_reg[417] = inform_L[464][8];				l_cell_reg[418] = inform_L[337][8];				l_cell_reg[419] = inform_L[465][8];				l_cell_reg[420] = inform_L[338][8];				l_cell_reg[421] = inform_L[466][8];				l_cell_reg[422] = inform_L[339][8];				l_cell_reg[423] = inform_L[467][8];				l_cell_reg[424] = inform_L[340][8];				l_cell_reg[425] = inform_L[468][8];				l_cell_reg[426] = inform_L[341][8];				l_cell_reg[427] = inform_L[469][8];				l_cell_reg[428] = inform_L[342][8];				l_cell_reg[429] = inform_L[470][8];				l_cell_reg[430] = inform_L[343][8];				l_cell_reg[431] = inform_L[471][8];				l_cell_reg[432] = inform_L[344][8];				l_cell_reg[433] = inform_L[472][8];				l_cell_reg[434] = inform_L[345][8];				l_cell_reg[435] = inform_L[473][8];				l_cell_reg[436] = inform_L[346][8];				l_cell_reg[437] = inform_L[474][8];				l_cell_reg[438] = inform_L[347][8];				l_cell_reg[439] = inform_L[475][8];				l_cell_reg[440] = inform_L[348][8];				l_cell_reg[441] = inform_L[476][8];				l_cell_reg[442] = inform_L[349][8];				l_cell_reg[443] = inform_L[477][8];				l_cell_reg[444] = inform_L[350][8];				l_cell_reg[445] = inform_L[478][8];				l_cell_reg[446] = inform_L[351][8];				l_cell_reg[447] = inform_L[479][8];				l_cell_reg[448] = inform_L[352][8];				l_cell_reg[449] = inform_L[480][8];				l_cell_reg[450] = inform_L[353][8];				l_cell_reg[451] = inform_L[481][8];				l_cell_reg[452] = inform_L[354][8];				l_cell_reg[453] = inform_L[482][8];				l_cell_reg[454] = inform_L[355][8];				l_cell_reg[455] = inform_L[483][8];				l_cell_reg[456] = inform_L[356][8];				l_cell_reg[457] = inform_L[484][8];				l_cell_reg[458] = inform_L[357][8];				l_cell_reg[459] = inform_L[485][8];				l_cell_reg[460] = inform_L[358][8];				l_cell_reg[461] = inform_L[486][8];				l_cell_reg[462] = inform_L[359][8];				l_cell_reg[463] = inform_L[487][8];				l_cell_reg[464] = inform_L[360][8];				l_cell_reg[465] = inform_L[488][8];				l_cell_reg[466] = inform_L[361][8];				l_cell_reg[467] = inform_L[489][8];				l_cell_reg[468] = inform_L[362][8];				l_cell_reg[469] = inform_L[490][8];				l_cell_reg[470] = inform_L[363][8];				l_cell_reg[471] = inform_L[491][8];				l_cell_reg[472] = inform_L[364][8];				l_cell_reg[473] = inform_L[492][8];				l_cell_reg[474] = inform_L[365][8];				l_cell_reg[475] = inform_L[493][8];				l_cell_reg[476] = inform_L[366][8];				l_cell_reg[477] = inform_L[494][8];				l_cell_reg[478] = inform_L[367][8];				l_cell_reg[479] = inform_L[495][8];				l_cell_reg[480] = inform_L[368][8];				l_cell_reg[481] = inform_L[496][8];				l_cell_reg[482] = inform_L[369][8];				l_cell_reg[483] = inform_L[497][8];				l_cell_reg[484] = inform_L[370][8];				l_cell_reg[485] = inform_L[498][8];				l_cell_reg[486] = inform_L[371][8];				l_cell_reg[487] = inform_L[499][8];				l_cell_reg[488] = inform_L[372][8];				l_cell_reg[489] = inform_L[500][8];				l_cell_reg[490] = inform_L[373][8];				l_cell_reg[491] = inform_L[501][8];				l_cell_reg[492] = inform_L[374][8];				l_cell_reg[493] = inform_L[502][8];				l_cell_reg[494] = inform_L[375][8];				l_cell_reg[495] = inform_L[503][8];				l_cell_reg[496] = inform_L[376][8];				l_cell_reg[497] = inform_L[504][8];				l_cell_reg[498] = inform_L[377][8];				l_cell_reg[499] = inform_L[505][8];				l_cell_reg[500] = inform_L[378][8];				l_cell_reg[501] = inform_L[506][8];				l_cell_reg[502] = inform_L[379][8];				l_cell_reg[503] = inform_L[507][8];				l_cell_reg[504] = inform_L[380][8];				l_cell_reg[505] = inform_L[508][8];				l_cell_reg[506] = inform_L[381][8];				l_cell_reg[507] = inform_L[509][8];				l_cell_reg[508] = inform_L[382][8];				l_cell_reg[509] = inform_L[510][8];				l_cell_reg[510] = inform_L[383][8];				l_cell_reg[511] = inform_L[511][8];				l_cell_reg[512] = inform_L[512][8];				l_cell_reg[513] = inform_L[640][8];				l_cell_reg[514] = inform_L[513][8];				l_cell_reg[515] = inform_L[641][8];				l_cell_reg[516] = inform_L[514][8];				l_cell_reg[517] = inform_L[642][8];				l_cell_reg[518] = inform_L[515][8];				l_cell_reg[519] = inform_L[643][8];				l_cell_reg[520] = inform_L[516][8];				l_cell_reg[521] = inform_L[644][8];				l_cell_reg[522] = inform_L[517][8];				l_cell_reg[523] = inform_L[645][8];				l_cell_reg[524] = inform_L[518][8];				l_cell_reg[525] = inform_L[646][8];				l_cell_reg[526] = inform_L[519][8];				l_cell_reg[527] = inform_L[647][8];				l_cell_reg[528] = inform_L[520][8];				l_cell_reg[529] = inform_L[648][8];				l_cell_reg[530] = inform_L[521][8];				l_cell_reg[531] = inform_L[649][8];				l_cell_reg[532] = inform_L[522][8];				l_cell_reg[533] = inform_L[650][8];				l_cell_reg[534] = inform_L[523][8];				l_cell_reg[535] = inform_L[651][8];				l_cell_reg[536] = inform_L[524][8];				l_cell_reg[537] = inform_L[652][8];				l_cell_reg[538] = inform_L[525][8];				l_cell_reg[539] = inform_L[653][8];				l_cell_reg[540] = inform_L[526][8];				l_cell_reg[541] = inform_L[654][8];				l_cell_reg[542] = inform_L[527][8];				l_cell_reg[543] = inform_L[655][8];				l_cell_reg[544] = inform_L[528][8];				l_cell_reg[545] = inform_L[656][8];				l_cell_reg[546] = inform_L[529][8];				l_cell_reg[547] = inform_L[657][8];				l_cell_reg[548] = inform_L[530][8];				l_cell_reg[549] = inform_L[658][8];				l_cell_reg[550] = inform_L[531][8];				l_cell_reg[551] = inform_L[659][8];				l_cell_reg[552] = inform_L[532][8];				l_cell_reg[553] = inform_L[660][8];				l_cell_reg[554] = inform_L[533][8];				l_cell_reg[555] = inform_L[661][8];				l_cell_reg[556] = inform_L[534][8];				l_cell_reg[557] = inform_L[662][8];				l_cell_reg[558] = inform_L[535][8];				l_cell_reg[559] = inform_L[663][8];				l_cell_reg[560] = inform_L[536][8];				l_cell_reg[561] = inform_L[664][8];				l_cell_reg[562] = inform_L[537][8];				l_cell_reg[563] = inform_L[665][8];				l_cell_reg[564] = inform_L[538][8];				l_cell_reg[565] = inform_L[666][8];				l_cell_reg[566] = inform_L[539][8];				l_cell_reg[567] = inform_L[667][8];				l_cell_reg[568] = inform_L[540][8];				l_cell_reg[569] = inform_L[668][8];				l_cell_reg[570] = inform_L[541][8];				l_cell_reg[571] = inform_L[669][8];				l_cell_reg[572] = inform_L[542][8];				l_cell_reg[573] = inform_L[670][8];				l_cell_reg[574] = inform_L[543][8];				l_cell_reg[575] = inform_L[671][8];				l_cell_reg[576] = inform_L[544][8];				l_cell_reg[577] = inform_L[672][8];				l_cell_reg[578] = inform_L[545][8];				l_cell_reg[579] = inform_L[673][8];				l_cell_reg[580] = inform_L[546][8];				l_cell_reg[581] = inform_L[674][8];				l_cell_reg[582] = inform_L[547][8];				l_cell_reg[583] = inform_L[675][8];				l_cell_reg[584] = inform_L[548][8];				l_cell_reg[585] = inform_L[676][8];				l_cell_reg[586] = inform_L[549][8];				l_cell_reg[587] = inform_L[677][8];				l_cell_reg[588] = inform_L[550][8];				l_cell_reg[589] = inform_L[678][8];				l_cell_reg[590] = inform_L[551][8];				l_cell_reg[591] = inform_L[679][8];				l_cell_reg[592] = inform_L[552][8];				l_cell_reg[593] = inform_L[680][8];				l_cell_reg[594] = inform_L[553][8];				l_cell_reg[595] = inform_L[681][8];				l_cell_reg[596] = inform_L[554][8];				l_cell_reg[597] = inform_L[682][8];				l_cell_reg[598] = inform_L[555][8];				l_cell_reg[599] = inform_L[683][8];				l_cell_reg[600] = inform_L[556][8];				l_cell_reg[601] = inform_L[684][8];				l_cell_reg[602] = inform_L[557][8];				l_cell_reg[603] = inform_L[685][8];				l_cell_reg[604] = inform_L[558][8];				l_cell_reg[605] = inform_L[686][8];				l_cell_reg[606] = inform_L[559][8];				l_cell_reg[607] = inform_L[687][8];				l_cell_reg[608] = inform_L[560][8];				l_cell_reg[609] = inform_L[688][8];				l_cell_reg[610] = inform_L[561][8];				l_cell_reg[611] = inform_L[689][8];				l_cell_reg[612] = inform_L[562][8];				l_cell_reg[613] = inform_L[690][8];				l_cell_reg[614] = inform_L[563][8];				l_cell_reg[615] = inform_L[691][8];				l_cell_reg[616] = inform_L[564][8];				l_cell_reg[617] = inform_L[692][8];				l_cell_reg[618] = inform_L[565][8];				l_cell_reg[619] = inform_L[693][8];				l_cell_reg[620] = inform_L[566][8];				l_cell_reg[621] = inform_L[694][8];				l_cell_reg[622] = inform_L[567][8];				l_cell_reg[623] = inform_L[695][8];				l_cell_reg[624] = inform_L[568][8];				l_cell_reg[625] = inform_L[696][8];				l_cell_reg[626] = inform_L[569][8];				l_cell_reg[627] = inform_L[697][8];				l_cell_reg[628] = inform_L[570][8];				l_cell_reg[629] = inform_L[698][8];				l_cell_reg[630] = inform_L[571][8];				l_cell_reg[631] = inform_L[699][8];				l_cell_reg[632] = inform_L[572][8];				l_cell_reg[633] = inform_L[700][8];				l_cell_reg[634] = inform_L[573][8];				l_cell_reg[635] = inform_L[701][8];				l_cell_reg[636] = inform_L[574][8];				l_cell_reg[637] = inform_L[702][8];				l_cell_reg[638] = inform_L[575][8];				l_cell_reg[639] = inform_L[703][8];				l_cell_reg[640] = inform_L[576][8];				l_cell_reg[641] = inform_L[704][8];				l_cell_reg[642] = inform_L[577][8];				l_cell_reg[643] = inform_L[705][8];				l_cell_reg[644] = inform_L[578][8];				l_cell_reg[645] = inform_L[706][8];				l_cell_reg[646] = inform_L[579][8];				l_cell_reg[647] = inform_L[707][8];				l_cell_reg[648] = inform_L[580][8];				l_cell_reg[649] = inform_L[708][8];				l_cell_reg[650] = inform_L[581][8];				l_cell_reg[651] = inform_L[709][8];				l_cell_reg[652] = inform_L[582][8];				l_cell_reg[653] = inform_L[710][8];				l_cell_reg[654] = inform_L[583][8];				l_cell_reg[655] = inform_L[711][8];				l_cell_reg[656] = inform_L[584][8];				l_cell_reg[657] = inform_L[712][8];				l_cell_reg[658] = inform_L[585][8];				l_cell_reg[659] = inform_L[713][8];				l_cell_reg[660] = inform_L[586][8];				l_cell_reg[661] = inform_L[714][8];				l_cell_reg[662] = inform_L[587][8];				l_cell_reg[663] = inform_L[715][8];				l_cell_reg[664] = inform_L[588][8];				l_cell_reg[665] = inform_L[716][8];				l_cell_reg[666] = inform_L[589][8];				l_cell_reg[667] = inform_L[717][8];				l_cell_reg[668] = inform_L[590][8];				l_cell_reg[669] = inform_L[718][8];				l_cell_reg[670] = inform_L[591][8];				l_cell_reg[671] = inform_L[719][8];				l_cell_reg[672] = inform_L[592][8];				l_cell_reg[673] = inform_L[720][8];				l_cell_reg[674] = inform_L[593][8];				l_cell_reg[675] = inform_L[721][8];				l_cell_reg[676] = inform_L[594][8];				l_cell_reg[677] = inform_L[722][8];				l_cell_reg[678] = inform_L[595][8];				l_cell_reg[679] = inform_L[723][8];				l_cell_reg[680] = inform_L[596][8];				l_cell_reg[681] = inform_L[724][8];				l_cell_reg[682] = inform_L[597][8];				l_cell_reg[683] = inform_L[725][8];				l_cell_reg[684] = inform_L[598][8];				l_cell_reg[685] = inform_L[726][8];				l_cell_reg[686] = inform_L[599][8];				l_cell_reg[687] = inform_L[727][8];				l_cell_reg[688] = inform_L[600][8];				l_cell_reg[689] = inform_L[728][8];				l_cell_reg[690] = inform_L[601][8];				l_cell_reg[691] = inform_L[729][8];				l_cell_reg[692] = inform_L[602][8];				l_cell_reg[693] = inform_L[730][8];				l_cell_reg[694] = inform_L[603][8];				l_cell_reg[695] = inform_L[731][8];				l_cell_reg[696] = inform_L[604][8];				l_cell_reg[697] = inform_L[732][8];				l_cell_reg[698] = inform_L[605][8];				l_cell_reg[699] = inform_L[733][8];				l_cell_reg[700] = inform_L[606][8];				l_cell_reg[701] = inform_L[734][8];				l_cell_reg[702] = inform_L[607][8];				l_cell_reg[703] = inform_L[735][8];				l_cell_reg[704] = inform_L[608][8];				l_cell_reg[705] = inform_L[736][8];				l_cell_reg[706] = inform_L[609][8];				l_cell_reg[707] = inform_L[737][8];				l_cell_reg[708] = inform_L[610][8];				l_cell_reg[709] = inform_L[738][8];				l_cell_reg[710] = inform_L[611][8];				l_cell_reg[711] = inform_L[739][8];				l_cell_reg[712] = inform_L[612][8];				l_cell_reg[713] = inform_L[740][8];				l_cell_reg[714] = inform_L[613][8];				l_cell_reg[715] = inform_L[741][8];				l_cell_reg[716] = inform_L[614][8];				l_cell_reg[717] = inform_L[742][8];				l_cell_reg[718] = inform_L[615][8];				l_cell_reg[719] = inform_L[743][8];				l_cell_reg[720] = inform_L[616][8];				l_cell_reg[721] = inform_L[744][8];				l_cell_reg[722] = inform_L[617][8];				l_cell_reg[723] = inform_L[745][8];				l_cell_reg[724] = inform_L[618][8];				l_cell_reg[725] = inform_L[746][8];				l_cell_reg[726] = inform_L[619][8];				l_cell_reg[727] = inform_L[747][8];				l_cell_reg[728] = inform_L[620][8];				l_cell_reg[729] = inform_L[748][8];				l_cell_reg[730] = inform_L[621][8];				l_cell_reg[731] = inform_L[749][8];				l_cell_reg[732] = inform_L[622][8];				l_cell_reg[733] = inform_L[750][8];				l_cell_reg[734] = inform_L[623][8];				l_cell_reg[735] = inform_L[751][8];				l_cell_reg[736] = inform_L[624][8];				l_cell_reg[737] = inform_L[752][8];				l_cell_reg[738] = inform_L[625][8];				l_cell_reg[739] = inform_L[753][8];				l_cell_reg[740] = inform_L[626][8];				l_cell_reg[741] = inform_L[754][8];				l_cell_reg[742] = inform_L[627][8];				l_cell_reg[743] = inform_L[755][8];				l_cell_reg[744] = inform_L[628][8];				l_cell_reg[745] = inform_L[756][8];				l_cell_reg[746] = inform_L[629][8];				l_cell_reg[747] = inform_L[757][8];				l_cell_reg[748] = inform_L[630][8];				l_cell_reg[749] = inform_L[758][8];				l_cell_reg[750] = inform_L[631][8];				l_cell_reg[751] = inform_L[759][8];				l_cell_reg[752] = inform_L[632][8];				l_cell_reg[753] = inform_L[760][8];				l_cell_reg[754] = inform_L[633][8];				l_cell_reg[755] = inform_L[761][8];				l_cell_reg[756] = inform_L[634][8];				l_cell_reg[757] = inform_L[762][8];				l_cell_reg[758] = inform_L[635][8];				l_cell_reg[759] = inform_L[763][8];				l_cell_reg[760] = inform_L[636][8];				l_cell_reg[761] = inform_L[764][8];				l_cell_reg[762] = inform_L[637][8];				l_cell_reg[763] = inform_L[765][8];				l_cell_reg[764] = inform_L[638][8];				l_cell_reg[765] = inform_L[766][8];				l_cell_reg[766] = inform_L[639][8];				l_cell_reg[767] = inform_L[767][8];				l_cell_reg[768] = inform_L[768][8];				l_cell_reg[769] = inform_L[896][8];				l_cell_reg[770] = inform_L[769][8];				l_cell_reg[771] = inform_L[897][8];				l_cell_reg[772] = inform_L[770][8];				l_cell_reg[773] = inform_L[898][8];				l_cell_reg[774] = inform_L[771][8];				l_cell_reg[775] = inform_L[899][8];				l_cell_reg[776] = inform_L[772][8];				l_cell_reg[777] = inform_L[900][8];				l_cell_reg[778] = inform_L[773][8];				l_cell_reg[779] = inform_L[901][8];				l_cell_reg[780] = inform_L[774][8];				l_cell_reg[781] = inform_L[902][8];				l_cell_reg[782] = inform_L[775][8];				l_cell_reg[783] = inform_L[903][8];				l_cell_reg[784] = inform_L[776][8];				l_cell_reg[785] = inform_L[904][8];				l_cell_reg[786] = inform_L[777][8];				l_cell_reg[787] = inform_L[905][8];				l_cell_reg[788] = inform_L[778][8];				l_cell_reg[789] = inform_L[906][8];				l_cell_reg[790] = inform_L[779][8];				l_cell_reg[791] = inform_L[907][8];				l_cell_reg[792] = inform_L[780][8];				l_cell_reg[793] = inform_L[908][8];				l_cell_reg[794] = inform_L[781][8];				l_cell_reg[795] = inform_L[909][8];				l_cell_reg[796] = inform_L[782][8];				l_cell_reg[797] = inform_L[910][8];				l_cell_reg[798] = inform_L[783][8];				l_cell_reg[799] = inform_L[911][8];				l_cell_reg[800] = inform_L[784][8];				l_cell_reg[801] = inform_L[912][8];				l_cell_reg[802] = inform_L[785][8];				l_cell_reg[803] = inform_L[913][8];				l_cell_reg[804] = inform_L[786][8];				l_cell_reg[805] = inform_L[914][8];				l_cell_reg[806] = inform_L[787][8];				l_cell_reg[807] = inform_L[915][8];				l_cell_reg[808] = inform_L[788][8];				l_cell_reg[809] = inform_L[916][8];				l_cell_reg[810] = inform_L[789][8];				l_cell_reg[811] = inform_L[917][8];				l_cell_reg[812] = inform_L[790][8];				l_cell_reg[813] = inform_L[918][8];				l_cell_reg[814] = inform_L[791][8];				l_cell_reg[815] = inform_L[919][8];				l_cell_reg[816] = inform_L[792][8];				l_cell_reg[817] = inform_L[920][8];				l_cell_reg[818] = inform_L[793][8];				l_cell_reg[819] = inform_L[921][8];				l_cell_reg[820] = inform_L[794][8];				l_cell_reg[821] = inform_L[922][8];				l_cell_reg[822] = inform_L[795][8];				l_cell_reg[823] = inform_L[923][8];				l_cell_reg[824] = inform_L[796][8];				l_cell_reg[825] = inform_L[924][8];				l_cell_reg[826] = inform_L[797][8];				l_cell_reg[827] = inform_L[925][8];				l_cell_reg[828] = inform_L[798][8];				l_cell_reg[829] = inform_L[926][8];				l_cell_reg[830] = inform_L[799][8];				l_cell_reg[831] = inform_L[927][8];				l_cell_reg[832] = inform_L[800][8];				l_cell_reg[833] = inform_L[928][8];				l_cell_reg[834] = inform_L[801][8];				l_cell_reg[835] = inform_L[929][8];				l_cell_reg[836] = inform_L[802][8];				l_cell_reg[837] = inform_L[930][8];				l_cell_reg[838] = inform_L[803][8];				l_cell_reg[839] = inform_L[931][8];				l_cell_reg[840] = inform_L[804][8];				l_cell_reg[841] = inform_L[932][8];				l_cell_reg[842] = inform_L[805][8];				l_cell_reg[843] = inform_L[933][8];				l_cell_reg[844] = inform_L[806][8];				l_cell_reg[845] = inform_L[934][8];				l_cell_reg[846] = inform_L[807][8];				l_cell_reg[847] = inform_L[935][8];				l_cell_reg[848] = inform_L[808][8];				l_cell_reg[849] = inform_L[936][8];				l_cell_reg[850] = inform_L[809][8];				l_cell_reg[851] = inform_L[937][8];				l_cell_reg[852] = inform_L[810][8];				l_cell_reg[853] = inform_L[938][8];				l_cell_reg[854] = inform_L[811][8];				l_cell_reg[855] = inform_L[939][8];				l_cell_reg[856] = inform_L[812][8];				l_cell_reg[857] = inform_L[940][8];				l_cell_reg[858] = inform_L[813][8];				l_cell_reg[859] = inform_L[941][8];				l_cell_reg[860] = inform_L[814][8];				l_cell_reg[861] = inform_L[942][8];				l_cell_reg[862] = inform_L[815][8];				l_cell_reg[863] = inform_L[943][8];				l_cell_reg[864] = inform_L[816][8];				l_cell_reg[865] = inform_L[944][8];				l_cell_reg[866] = inform_L[817][8];				l_cell_reg[867] = inform_L[945][8];				l_cell_reg[868] = inform_L[818][8];				l_cell_reg[869] = inform_L[946][8];				l_cell_reg[870] = inform_L[819][8];				l_cell_reg[871] = inform_L[947][8];				l_cell_reg[872] = inform_L[820][8];				l_cell_reg[873] = inform_L[948][8];				l_cell_reg[874] = inform_L[821][8];				l_cell_reg[875] = inform_L[949][8];				l_cell_reg[876] = inform_L[822][8];				l_cell_reg[877] = inform_L[950][8];				l_cell_reg[878] = inform_L[823][8];				l_cell_reg[879] = inform_L[951][8];				l_cell_reg[880] = inform_L[824][8];				l_cell_reg[881] = inform_L[952][8];				l_cell_reg[882] = inform_L[825][8];				l_cell_reg[883] = inform_L[953][8];				l_cell_reg[884] = inform_L[826][8];				l_cell_reg[885] = inform_L[954][8];				l_cell_reg[886] = inform_L[827][8];				l_cell_reg[887] = inform_L[955][8];				l_cell_reg[888] = inform_L[828][8];				l_cell_reg[889] = inform_L[956][8];				l_cell_reg[890] = inform_L[829][8];				l_cell_reg[891] = inform_L[957][8];				l_cell_reg[892] = inform_L[830][8];				l_cell_reg[893] = inform_L[958][8];				l_cell_reg[894] = inform_L[831][8];				l_cell_reg[895] = inform_L[959][8];				l_cell_reg[896] = inform_L[832][8];				l_cell_reg[897] = inform_L[960][8];				l_cell_reg[898] = inform_L[833][8];				l_cell_reg[899] = inform_L[961][8];				l_cell_reg[900] = inform_L[834][8];				l_cell_reg[901] = inform_L[962][8];				l_cell_reg[902] = inform_L[835][8];				l_cell_reg[903] = inform_L[963][8];				l_cell_reg[904] = inform_L[836][8];				l_cell_reg[905] = inform_L[964][8];				l_cell_reg[906] = inform_L[837][8];				l_cell_reg[907] = inform_L[965][8];				l_cell_reg[908] = inform_L[838][8];				l_cell_reg[909] = inform_L[966][8];				l_cell_reg[910] = inform_L[839][8];				l_cell_reg[911] = inform_L[967][8];				l_cell_reg[912] = inform_L[840][8];				l_cell_reg[913] = inform_L[968][8];				l_cell_reg[914] = inform_L[841][8];				l_cell_reg[915] = inform_L[969][8];				l_cell_reg[916] = inform_L[842][8];				l_cell_reg[917] = inform_L[970][8];				l_cell_reg[918] = inform_L[843][8];				l_cell_reg[919] = inform_L[971][8];				l_cell_reg[920] = inform_L[844][8];				l_cell_reg[921] = inform_L[972][8];				l_cell_reg[922] = inform_L[845][8];				l_cell_reg[923] = inform_L[973][8];				l_cell_reg[924] = inform_L[846][8];				l_cell_reg[925] = inform_L[974][8];				l_cell_reg[926] = inform_L[847][8];				l_cell_reg[927] = inform_L[975][8];				l_cell_reg[928] = inform_L[848][8];				l_cell_reg[929] = inform_L[976][8];				l_cell_reg[930] = inform_L[849][8];				l_cell_reg[931] = inform_L[977][8];				l_cell_reg[932] = inform_L[850][8];				l_cell_reg[933] = inform_L[978][8];				l_cell_reg[934] = inform_L[851][8];				l_cell_reg[935] = inform_L[979][8];				l_cell_reg[936] = inform_L[852][8];				l_cell_reg[937] = inform_L[980][8];				l_cell_reg[938] = inform_L[853][8];				l_cell_reg[939] = inform_L[981][8];				l_cell_reg[940] = inform_L[854][8];				l_cell_reg[941] = inform_L[982][8];				l_cell_reg[942] = inform_L[855][8];				l_cell_reg[943] = inform_L[983][8];				l_cell_reg[944] = inform_L[856][8];				l_cell_reg[945] = inform_L[984][8];				l_cell_reg[946] = inform_L[857][8];				l_cell_reg[947] = inform_L[985][8];				l_cell_reg[948] = inform_L[858][8];				l_cell_reg[949] = inform_L[986][8];				l_cell_reg[950] = inform_L[859][8];				l_cell_reg[951] = inform_L[987][8];				l_cell_reg[952] = inform_L[860][8];				l_cell_reg[953] = inform_L[988][8];				l_cell_reg[954] = inform_L[861][8];				l_cell_reg[955] = inform_L[989][8];				l_cell_reg[956] = inform_L[862][8];				l_cell_reg[957] = inform_L[990][8];				l_cell_reg[958] = inform_L[863][8];				l_cell_reg[959] = inform_L[991][8];				l_cell_reg[960] = inform_L[864][8];				l_cell_reg[961] = inform_L[992][8];				l_cell_reg[962] = inform_L[865][8];				l_cell_reg[963] = inform_L[993][8];				l_cell_reg[964] = inform_L[866][8];				l_cell_reg[965] = inform_L[994][8];				l_cell_reg[966] = inform_L[867][8];				l_cell_reg[967] = inform_L[995][8];				l_cell_reg[968] = inform_L[868][8];				l_cell_reg[969] = inform_L[996][8];				l_cell_reg[970] = inform_L[869][8];				l_cell_reg[971] = inform_L[997][8];				l_cell_reg[972] = inform_L[870][8];				l_cell_reg[973] = inform_L[998][8];				l_cell_reg[974] = inform_L[871][8];				l_cell_reg[975] = inform_L[999][8];				l_cell_reg[976] = inform_L[872][8];				l_cell_reg[977] = inform_L[1000][8];				l_cell_reg[978] = inform_L[873][8];				l_cell_reg[979] = inform_L[1001][8];				l_cell_reg[980] = inform_L[874][8];				l_cell_reg[981] = inform_L[1002][8];				l_cell_reg[982] = inform_L[875][8];				l_cell_reg[983] = inform_L[1003][8];				l_cell_reg[984] = inform_L[876][8];				l_cell_reg[985] = inform_L[1004][8];				l_cell_reg[986] = inform_L[877][8];				l_cell_reg[987] = inform_L[1005][8];				l_cell_reg[988] = inform_L[878][8];				l_cell_reg[989] = inform_L[1006][8];				l_cell_reg[990] = inform_L[879][8];				l_cell_reg[991] = inform_L[1007][8];				l_cell_reg[992] = inform_L[880][8];				l_cell_reg[993] = inform_L[1008][8];				l_cell_reg[994] = inform_L[881][8];				l_cell_reg[995] = inform_L[1009][8];				l_cell_reg[996] = inform_L[882][8];				l_cell_reg[997] = inform_L[1010][8];				l_cell_reg[998] = inform_L[883][8];				l_cell_reg[999] = inform_L[1011][8];				l_cell_reg[1000] = inform_L[884][8];				l_cell_reg[1001] = inform_L[1012][8];				l_cell_reg[1002] = inform_L[885][8];				l_cell_reg[1003] = inform_L[1013][8];				l_cell_reg[1004] = inform_L[886][8];				l_cell_reg[1005] = inform_L[1014][8];				l_cell_reg[1006] = inform_L[887][8];				l_cell_reg[1007] = inform_L[1015][8];				l_cell_reg[1008] = inform_L[888][8];				l_cell_reg[1009] = inform_L[1016][8];				l_cell_reg[1010] = inform_L[889][8];				l_cell_reg[1011] = inform_L[1017][8];				l_cell_reg[1012] = inform_L[890][8];				l_cell_reg[1013] = inform_L[1018][8];				l_cell_reg[1014] = inform_L[891][8];				l_cell_reg[1015] = inform_L[1019][8];				l_cell_reg[1016] = inform_L[892][8];				l_cell_reg[1017] = inform_L[1020][8];				l_cell_reg[1018] = inform_L[893][8];				l_cell_reg[1019] = inform_L[1021][8];				l_cell_reg[1020] = inform_L[894][8];				l_cell_reg[1021] = inform_L[1022][8];				l_cell_reg[1022] = inform_L[895][8];				l_cell_reg[1023] = inform_L[1023][8];			end
			9:			begin				r_cell_reg[0] = inform_R[0][8];				r_cell_reg[1] = inform_R[256][8];				r_cell_reg[2] = inform_R[1][8];				r_cell_reg[3] = inform_R[257][8];				r_cell_reg[4] = inform_R[2][8];				r_cell_reg[5] = inform_R[258][8];				r_cell_reg[6] = inform_R[3][8];				r_cell_reg[7] = inform_R[259][8];				r_cell_reg[8] = inform_R[4][8];				r_cell_reg[9] = inform_R[260][8];				r_cell_reg[10] = inform_R[5][8];				r_cell_reg[11] = inform_R[261][8];				r_cell_reg[12] = inform_R[6][8];				r_cell_reg[13] = inform_R[262][8];				r_cell_reg[14] = inform_R[7][8];				r_cell_reg[15] = inform_R[263][8];				r_cell_reg[16] = inform_R[8][8];				r_cell_reg[17] = inform_R[264][8];				r_cell_reg[18] = inform_R[9][8];				r_cell_reg[19] = inform_R[265][8];				r_cell_reg[20] = inform_R[10][8];				r_cell_reg[21] = inform_R[266][8];				r_cell_reg[22] = inform_R[11][8];				r_cell_reg[23] = inform_R[267][8];				r_cell_reg[24] = inform_R[12][8];				r_cell_reg[25] = inform_R[268][8];				r_cell_reg[26] = inform_R[13][8];				r_cell_reg[27] = inform_R[269][8];				r_cell_reg[28] = inform_R[14][8];				r_cell_reg[29] = inform_R[270][8];				r_cell_reg[30] = inform_R[15][8];				r_cell_reg[31] = inform_R[271][8];				r_cell_reg[32] = inform_R[16][8];				r_cell_reg[33] = inform_R[272][8];				r_cell_reg[34] = inform_R[17][8];				r_cell_reg[35] = inform_R[273][8];				r_cell_reg[36] = inform_R[18][8];				r_cell_reg[37] = inform_R[274][8];				r_cell_reg[38] = inform_R[19][8];				r_cell_reg[39] = inform_R[275][8];				r_cell_reg[40] = inform_R[20][8];				r_cell_reg[41] = inform_R[276][8];				r_cell_reg[42] = inform_R[21][8];				r_cell_reg[43] = inform_R[277][8];				r_cell_reg[44] = inform_R[22][8];				r_cell_reg[45] = inform_R[278][8];				r_cell_reg[46] = inform_R[23][8];				r_cell_reg[47] = inform_R[279][8];				r_cell_reg[48] = inform_R[24][8];				r_cell_reg[49] = inform_R[280][8];				r_cell_reg[50] = inform_R[25][8];				r_cell_reg[51] = inform_R[281][8];				r_cell_reg[52] = inform_R[26][8];				r_cell_reg[53] = inform_R[282][8];				r_cell_reg[54] = inform_R[27][8];				r_cell_reg[55] = inform_R[283][8];				r_cell_reg[56] = inform_R[28][8];				r_cell_reg[57] = inform_R[284][8];				r_cell_reg[58] = inform_R[29][8];				r_cell_reg[59] = inform_R[285][8];				r_cell_reg[60] = inform_R[30][8];				r_cell_reg[61] = inform_R[286][8];				r_cell_reg[62] = inform_R[31][8];				r_cell_reg[63] = inform_R[287][8];				r_cell_reg[64] = inform_R[32][8];				r_cell_reg[65] = inform_R[288][8];				r_cell_reg[66] = inform_R[33][8];				r_cell_reg[67] = inform_R[289][8];				r_cell_reg[68] = inform_R[34][8];				r_cell_reg[69] = inform_R[290][8];				r_cell_reg[70] = inform_R[35][8];				r_cell_reg[71] = inform_R[291][8];				r_cell_reg[72] = inform_R[36][8];				r_cell_reg[73] = inform_R[292][8];				r_cell_reg[74] = inform_R[37][8];				r_cell_reg[75] = inform_R[293][8];				r_cell_reg[76] = inform_R[38][8];				r_cell_reg[77] = inform_R[294][8];				r_cell_reg[78] = inform_R[39][8];				r_cell_reg[79] = inform_R[295][8];				r_cell_reg[80] = inform_R[40][8];				r_cell_reg[81] = inform_R[296][8];				r_cell_reg[82] = inform_R[41][8];				r_cell_reg[83] = inform_R[297][8];				r_cell_reg[84] = inform_R[42][8];				r_cell_reg[85] = inform_R[298][8];				r_cell_reg[86] = inform_R[43][8];				r_cell_reg[87] = inform_R[299][8];				r_cell_reg[88] = inform_R[44][8];				r_cell_reg[89] = inform_R[300][8];				r_cell_reg[90] = inform_R[45][8];				r_cell_reg[91] = inform_R[301][8];				r_cell_reg[92] = inform_R[46][8];				r_cell_reg[93] = inform_R[302][8];				r_cell_reg[94] = inform_R[47][8];				r_cell_reg[95] = inform_R[303][8];				r_cell_reg[96] = inform_R[48][8];				r_cell_reg[97] = inform_R[304][8];				r_cell_reg[98] = inform_R[49][8];				r_cell_reg[99] = inform_R[305][8];				r_cell_reg[100] = inform_R[50][8];				r_cell_reg[101] = inform_R[306][8];				r_cell_reg[102] = inform_R[51][8];				r_cell_reg[103] = inform_R[307][8];				r_cell_reg[104] = inform_R[52][8];				r_cell_reg[105] = inform_R[308][8];				r_cell_reg[106] = inform_R[53][8];				r_cell_reg[107] = inform_R[309][8];				r_cell_reg[108] = inform_R[54][8];				r_cell_reg[109] = inform_R[310][8];				r_cell_reg[110] = inform_R[55][8];				r_cell_reg[111] = inform_R[311][8];				r_cell_reg[112] = inform_R[56][8];				r_cell_reg[113] = inform_R[312][8];				r_cell_reg[114] = inform_R[57][8];				r_cell_reg[115] = inform_R[313][8];				r_cell_reg[116] = inform_R[58][8];				r_cell_reg[117] = inform_R[314][8];				r_cell_reg[118] = inform_R[59][8];				r_cell_reg[119] = inform_R[315][8];				r_cell_reg[120] = inform_R[60][8];				r_cell_reg[121] = inform_R[316][8];				r_cell_reg[122] = inform_R[61][8];				r_cell_reg[123] = inform_R[317][8];				r_cell_reg[124] = inform_R[62][8];				r_cell_reg[125] = inform_R[318][8];				r_cell_reg[126] = inform_R[63][8];				r_cell_reg[127] = inform_R[319][8];				r_cell_reg[128] = inform_R[64][8];				r_cell_reg[129] = inform_R[320][8];				r_cell_reg[130] = inform_R[65][8];				r_cell_reg[131] = inform_R[321][8];				r_cell_reg[132] = inform_R[66][8];				r_cell_reg[133] = inform_R[322][8];				r_cell_reg[134] = inform_R[67][8];				r_cell_reg[135] = inform_R[323][8];				r_cell_reg[136] = inform_R[68][8];				r_cell_reg[137] = inform_R[324][8];				r_cell_reg[138] = inform_R[69][8];				r_cell_reg[139] = inform_R[325][8];				r_cell_reg[140] = inform_R[70][8];				r_cell_reg[141] = inform_R[326][8];				r_cell_reg[142] = inform_R[71][8];				r_cell_reg[143] = inform_R[327][8];				r_cell_reg[144] = inform_R[72][8];				r_cell_reg[145] = inform_R[328][8];				r_cell_reg[146] = inform_R[73][8];				r_cell_reg[147] = inform_R[329][8];				r_cell_reg[148] = inform_R[74][8];				r_cell_reg[149] = inform_R[330][8];				r_cell_reg[150] = inform_R[75][8];				r_cell_reg[151] = inform_R[331][8];				r_cell_reg[152] = inform_R[76][8];				r_cell_reg[153] = inform_R[332][8];				r_cell_reg[154] = inform_R[77][8];				r_cell_reg[155] = inform_R[333][8];				r_cell_reg[156] = inform_R[78][8];				r_cell_reg[157] = inform_R[334][8];				r_cell_reg[158] = inform_R[79][8];				r_cell_reg[159] = inform_R[335][8];				r_cell_reg[160] = inform_R[80][8];				r_cell_reg[161] = inform_R[336][8];				r_cell_reg[162] = inform_R[81][8];				r_cell_reg[163] = inform_R[337][8];				r_cell_reg[164] = inform_R[82][8];				r_cell_reg[165] = inform_R[338][8];				r_cell_reg[166] = inform_R[83][8];				r_cell_reg[167] = inform_R[339][8];				r_cell_reg[168] = inform_R[84][8];				r_cell_reg[169] = inform_R[340][8];				r_cell_reg[170] = inform_R[85][8];				r_cell_reg[171] = inform_R[341][8];				r_cell_reg[172] = inform_R[86][8];				r_cell_reg[173] = inform_R[342][8];				r_cell_reg[174] = inform_R[87][8];				r_cell_reg[175] = inform_R[343][8];				r_cell_reg[176] = inform_R[88][8];				r_cell_reg[177] = inform_R[344][8];				r_cell_reg[178] = inform_R[89][8];				r_cell_reg[179] = inform_R[345][8];				r_cell_reg[180] = inform_R[90][8];				r_cell_reg[181] = inform_R[346][8];				r_cell_reg[182] = inform_R[91][8];				r_cell_reg[183] = inform_R[347][8];				r_cell_reg[184] = inform_R[92][8];				r_cell_reg[185] = inform_R[348][8];				r_cell_reg[186] = inform_R[93][8];				r_cell_reg[187] = inform_R[349][8];				r_cell_reg[188] = inform_R[94][8];				r_cell_reg[189] = inform_R[350][8];				r_cell_reg[190] = inform_R[95][8];				r_cell_reg[191] = inform_R[351][8];				r_cell_reg[192] = inform_R[96][8];				r_cell_reg[193] = inform_R[352][8];				r_cell_reg[194] = inform_R[97][8];				r_cell_reg[195] = inform_R[353][8];				r_cell_reg[196] = inform_R[98][8];				r_cell_reg[197] = inform_R[354][8];				r_cell_reg[198] = inform_R[99][8];				r_cell_reg[199] = inform_R[355][8];				r_cell_reg[200] = inform_R[100][8];				r_cell_reg[201] = inform_R[356][8];				r_cell_reg[202] = inform_R[101][8];				r_cell_reg[203] = inform_R[357][8];				r_cell_reg[204] = inform_R[102][8];				r_cell_reg[205] = inform_R[358][8];				r_cell_reg[206] = inform_R[103][8];				r_cell_reg[207] = inform_R[359][8];				r_cell_reg[208] = inform_R[104][8];				r_cell_reg[209] = inform_R[360][8];				r_cell_reg[210] = inform_R[105][8];				r_cell_reg[211] = inform_R[361][8];				r_cell_reg[212] = inform_R[106][8];				r_cell_reg[213] = inform_R[362][8];				r_cell_reg[214] = inform_R[107][8];				r_cell_reg[215] = inform_R[363][8];				r_cell_reg[216] = inform_R[108][8];				r_cell_reg[217] = inform_R[364][8];				r_cell_reg[218] = inform_R[109][8];				r_cell_reg[219] = inform_R[365][8];				r_cell_reg[220] = inform_R[110][8];				r_cell_reg[221] = inform_R[366][8];				r_cell_reg[222] = inform_R[111][8];				r_cell_reg[223] = inform_R[367][8];				r_cell_reg[224] = inform_R[112][8];				r_cell_reg[225] = inform_R[368][8];				r_cell_reg[226] = inform_R[113][8];				r_cell_reg[227] = inform_R[369][8];				r_cell_reg[228] = inform_R[114][8];				r_cell_reg[229] = inform_R[370][8];				r_cell_reg[230] = inform_R[115][8];				r_cell_reg[231] = inform_R[371][8];				r_cell_reg[232] = inform_R[116][8];				r_cell_reg[233] = inform_R[372][8];				r_cell_reg[234] = inform_R[117][8];				r_cell_reg[235] = inform_R[373][8];				r_cell_reg[236] = inform_R[118][8];				r_cell_reg[237] = inform_R[374][8];				r_cell_reg[238] = inform_R[119][8];				r_cell_reg[239] = inform_R[375][8];				r_cell_reg[240] = inform_R[120][8];				r_cell_reg[241] = inform_R[376][8];				r_cell_reg[242] = inform_R[121][8];				r_cell_reg[243] = inform_R[377][8];				r_cell_reg[244] = inform_R[122][8];				r_cell_reg[245] = inform_R[378][8];				r_cell_reg[246] = inform_R[123][8];				r_cell_reg[247] = inform_R[379][8];				r_cell_reg[248] = inform_R[124][8];				r_cell_reg[249] = inform_R[380][8];				r_cell_reg[250] = inform_R[125][8];				r_cell_reg[251] = inform_R[381][8];				r_cell_reg[252] = inform_R[126][8];				r_cell_reg[253] = inform_R[382][8];				r_cell_reg[254] = inform_R[127][8];				r_cell_reg[255] = inform_R[383][8];				r_cell_reg[256] = inform_R[128][8];				r_cell_reg[257] = inform_R[384][8];				r_cell_reg[258] = inform_R[129][8];				r_cell_reg[259] = inform_R[385][8];				r_cell_reg[260] = inform_R[130][8];				r_cell_reg[261] = inform_R[386][8];				r_cell_reg[262] = inform_R[131][8];				r_cell_reg[263] = inform_R[387][8];				r_cell_reg[264] = inform_R[132][8];				r_cell_reg[265] = inform_R[388][8];				r_cell_reg[266] = inform_R[133][8];				r_cell_reg[267] = inform_R[389][8];				r_cell_reg[268] = inform_R[134][8];				r_cell_reg[269] = inform_R[390][8];				r_cell_reg[270] = inform_R[135][8];				r_cell_reg[271] = inform_R[391][8];				r_cell_reg[272] = inform_R[136][8];				r_cell_reg[273] = inform_R[392][8];				r_cell_reg[274] = inform_R[137][8];				r_cell_reg[275] = inform_R[393][8];				r_cell_reg[276] = inform_R[138][8];				r_cell_reg[277] = inform_R[394][8];				r_cell_reg[278] = inform_R[139][8];				r_cell_reg[279] = inform_R[395][8];				r_cell_reg[280] = inform_R[140][8];				r_cell_reg[281] = inform_R[396][8];				r_cell_reg[282] = inform_R[141][8];				r_cell_reg[283] = inform_R[397][8];				r_cell_reg[284] = inform_R[142][8];				r_cell_reg[285] = inform_R[398][8];				r_cell_reg[286] = inform_R[143][8];				r_cell_reg[287] = inform_R[399][8];				r_cell_reg[288] = inform_R[144][8];				r_cell_reg[289] = inform_R[400][8];				r_cell_reg[290] = inform_R[145][8];				r_cell_reg[291] = inform_R[401][8];				r_cell_reg[292] = inform_R[146][8];				r_cell_reg[293] = inform_R[402][8];				r_cell_reg[294] = inform_R[147][8];				r_cell_reg[295] = inform_R[403][8];				r_cell_reg[296] = inform_R[148][8];				r_cell_reg[297] = inform_R[404][8];				r_cell_reg[298] = inform_R[149][8];				r_cell_reg[299] = inform_R[405][8];				r_cell_reg[300] = inform_R[150][8];				r_cell_reg[301] = inform_R[406][8];				r_cell_reg[302] = inform_R[151][8];				r_cell_reg[303] = inform_R[407][8];				r_cell_reg[304] = inform_R[152][8];				r_cell_reg[305] = inform_R[408][8];				r_cell_reg[306] = inform_R[153][8];				r_cell_reg[307] = inform_R[409][8];				r_cell_reg[308] = inform_R[154][8];				r_cell_reg[309] = inform_R[410][8];				r_cell_reg[310] = inform_R[155][8];				r_cell_reg[311] = inform_R[411][8];				r_cell_reg[312] = inform_R[156][8];				r_cell_reg[313] = inform_R[412][8];				r_cell_reg[314] = inform_R[157][8];				r_cell_reg[315] = inform_R[413][8];				r_cell_reg[316] = inform_R[158][8];				r_cell_reg[317] = inform_R[414][8];				r_cell_reg[318] = inform_R[159][8];				r_cell_reg[319] = inform_R[415][8];				r_cell_reg[320] = inform_R[160][8];				r_cell_reg[321] = inform_R[416][8];				r_cell_reg[322] = inform_R[161][8];				r_cell_reg[323] = inform_R[417][8];				r_cell_reg[324] = inform_R[162][8];				r_cell_reg[325] = inform_R[418][8];				r_cell_reg[326] = inform_R[163][8];				r_cell_reg[327] = inform_R[419][8];				r_cell_reg[328] = inform_R[164][8];				r_cell_reg[329] = inform_R[420][8];				r_cell_reg[330] = inform_R[165][8];				r_cell_reg[331] = inform_R[421][8];				r_cell_reg[332] = inform_R[166][8];				r_cell_reg[333] = inform_R[422][8];				r_cell_reg[334] = inform_R[167][8];				r_cell_reg[335] = inform_R[423][8];				r_cell_reg[336] = inform_R[168][8];				r_cell_reg[337] = inform_R[424][8];				r_cell_reg[338] = inform_R[169][8];				r_cell_reg[339] = inform_R[425][8];				r_cell_reg[340] = inform_R[170][8];				r_cell_reg[341] = inform_R[426][8];				r_cell_reg[342] = inform_R[171][8];				r_cell_reg[343] = inform_R[427][8];				r_cell_reg[344] = inform_R[172][8];				r_cell_reg[345] = inform_R[428][8];				r_cell_reg[346] = inform_R[173][8];				r_cell_reg[347] = inform_R[429][8];				r_cell_reg[348] = inform_R[174][8];				r_cell_reg[349] = inform_R[430][8];				r_cell_reg[350] = inform_R[175][8];				r_cell_reg[351] = inform_R[431][8];				r_cell_reg[352] = inform_R[176][8];				r_cell_reg[353] = inform_R[432][8];				r_cell_reg[354] = inform_R[177][8];				r_cell_reg[355] = inform_R[433][8];				r_cell_reg[356] = inform_R[178][8];				r_cell_reg[357] = inform_R[434][8];				r_cell_reg[358] = inform_R[179][8];				r_cell_reg[359] = inform_R[435][8];				r_cell_reg[360] = inform_R[180][8];				r_cell_reg[361] = inform_R[436][8];				r_cell_reg[362] = inform_R[181][8];				r_cell_reg[363] = inform_R[437][8];				r_cell_reg[364] = inform_R[182][8];				r_cell_reg[365] = inform_R[438][8];				r_cell_reg[366] = inform_R[183][8];				r_cell_reg[367] = inform_R[439][8];				r_cell_reg[368] = inform_R[184][8];				r_cell_reg[369] = inform_R[440][8];				r_cell_reg[370] = inform_R[185][8];				r_cell_reg[371] = inform_R[441][8];				r_cell_reg[372] = inform_R[186][8];				r_cell_reg[373] = inform_R[442][8];				r_cell_reg[374] = inform_R[187][8];				r_cell_reg[375] = inform_R[443][8];				r_cell_reg[376] = inform_R[188][8];				r_cell_reg[377] = inform_R[444][8];				r_cell_reg[378] = inform_R[189][8];				r_cell_reg[379] = inform_R[445][8];				r_cell_reg[380] = inform_R[190][8];				r_cell_reg[381] = inform_R[446][8];				r_cell_reg[382] = inform_R[191][8];				r_cell_reg[383] = inform_R[447][8];				r_cell_reg[384] = inform_R[192][8];				r_cell_reg[385] = inform_R[448][8];				r_cell_reg[386] = inform_R[193][8];				r_cell_reg[387] = inform_R[449][8];				r_cell_reg[388] = inform_R[194][8];				r_cell_reg[389] = inform_R[450][8];				r_cell_reg[390] = inform_R[195][8];				r_cell_reg[391] = inform_R[451][8];				r_cell_reg[392] = inform_R[196][8];				r_cell_reg[393] = inform_R[452][8];				r_cell_reg[394] = inform_R[197][8];				r_cell_reg[395] = inform_R[453][8];				r_cell_reg[396] = inform_R[198][8];				r_cell_reg[397] = inform_R[454][8];				r_cell_reg[398] = inform_R[199][8];				r_cell_reg[399] = inform_R[455][8];				r_cell_reg[400] = inform_R[200][8];				r_cell_reg[401] = inform_R[456][8];				r_cell_reg[402] = inform_R[201][8];				r_cell_reg[403] = inform_R[457][8];				r_cell_reg[404] = inform_R[202][8];				r_cell_reg[405] = inform_R[458][8];				r_cell_reg[406] = inform_R[203][8];				r_cell_reg[407] = inform_R[459][8];				r_cell_reg[408] = inform_R[204][8];				r_cell_reg[409] = inform_R[460][8];				r_cell_reg[410] = inform_R[205][8];				r_cell_reg[411] = inform_R[461][8];				r_cell_reg[412] = inform_R[206][8];				r_cell_reg[413] = inform_R[462][8];				r_cell_reg[414] = inform_R[207][8];				r_cell_reg[415] = inform_R[463][8];				r_cell_reg[416] = inform_R[208][8];				r_cell_reg[417] = inform_R[464][8];				r_cell_reg[418] = inform_R[209][8];				r_cell_reg[419] = inform_R[465][8];				r_cell_reg[420] = inform_R[210][8];				r_cell_reg[421] = inform_R[466][8];				r_cell_reg[422] = inform_R[211][8];				r_cell_reg[423] = inform_R[467][8];				r_cell_reg[424] = inform_R[212][8];				r_cell_reg[425] = inform_R[468][8];				r_cell_reg[426] = inform_R[213][8];				r_cell_reg[427] = inform_R[469][8];				r_cell_reg[428] = inform_R[214][8];				r_cell_reg[429] = inform_R[470][8];				r_cell_reg[430] = inform_R[215][8];				r_cell_reg[431] = inform_R[471][8];				r_cell_reg[432] = inform_R[216][8];				r_cell_reg[433] = inform_R[472][8];				r_cell_reg[434] = inform_R[217][8];				r_cell_reg[435] = inform_R[473][8];				r_cell_reg[436] = inform_R[218][8];				r_cell_reg[437] = inform_R[474][8];				r_cell_reg[438] = inform_R[219][8];				r_cell_reg[439] = inform_R[475][8];				r_cell_reg[440] = inform_R[220][8];				r_cell_reg[441] = inform_R[476][8];				r_cell_reg[442] = inform_R[221][8];				r_cell_reg[443] = inform_R[477][8];				r_cell_reg[444] = inform_R[222][8];				r_cell_reg[445] = inform_R[478][8];				r_cell_reg[446] = inform_R[223][8];				r_cell_reg[447] = inform_R[479][8];				r_cell_reg[448] = inform_R[224][8];				r_cell_reg[449] = inform_R[480][8];				r_cell_reg[450] = inform_R[225][8];				r_cell_reg[451] = inform_R[481][8];				r_cell_reg[452] = inform_R[226][8];				r_cell_reg[453] = inform_R[482][8];				r_cell_reg[454] = inform_R[227][8];				r_cell_reg[455] = inform_R[483][8];				r_cell_reg[456] = inform_R[228][8];				r_cell_reg[457] = inform_R[484][8];				r_cell_reg[458] = inform_R[229][8];				r_cell_reg[459] = inform_R[485][8];				r_cell_reg[460] = inform_R[230][8];				r_cell_reg[461] = inform_R[486][8];				r_cell_reg[462] = inform_R[231][8];				r_cell_reg[463] = inform_R[487][8];				r_cell_reg[464] = inform_R[232][8];				r_cell_reg[465] = inform_R[488][8];				r_cell_reg[466] = inform_R[233][8];				r_cell_reg[467] = inform_R[489][8];				r_cell_reg[468] = inform_R[234][8];				r_cell_reg[469] = inform_R[490][8];				r_cell_reg[470] = inform_R[235][8];				r_cell_reg[471] = inform_R[491][8];				r_cell_reg[472] = inform_R[236][8];				r_cell_reg[473] = inform_R[492][8];				r_cell_reg[474] = inform_R[237][8];				r_cell_reg[475] = inform_R[493][8];				r_cell_reg[476] = inform_R[238][8];				r_cell_reg[477] = inform_R[494][8];				r_cell_reg[478] = inform_R[239][8];				r_cell_reg[479] = inform_R[495][8];				r_cell_reg[480] = inform_R[240][8];				r_cell_reg[481] = inform_R[496][8];				r_cell_reg[482] = inform_R[241][8];				r_cell_reg[483] = inform_R[497][8];				r_cell_reg[484] = inform_R[242][8];				r_cell_reg[485] = inform_R[498][8];				r_cell_reg[486] = inform_R[243][8];				r_cell_reg[487] = inform_R[499][8];				r_cell_reg[488] = inform_R[244][8];				r_cell_reg[489] = inform_R[500][8];				r_cell_reg[490] = inform_R[245][8];				r_cell_reg[491] = inform_R[501][8];				r_cell_reg[492] = inform_R[246][8];				r_cell_reg[493] = inform_R[502][8];				r_cell_reg[494] = inform_R[247][8];				r_cell_reg[495] = inform_R[503][8];				r_cell_reg[496] = inform_R[248][8];				r_cell_reg[497] = inform_R[504][8];				r_cell_reg[498] = inform_R[249][8];				r_cell_reg[499] = inform_R[505][8];				r_cell_reg[500] = inform_R[250][8];				r_cell_reg[501] = inform_R[506][8];				r_cell_reg[502] = inform_R[251][8];				r_cell_reg[503] = inform_R[507][8];				r_cell_reg[504] = inform_R[252][8];				r_cell_reg[505] = inform_R[508][8];				r_cell_reg[506] = inform_R[253][8];				r_cell_reg[507] = inform_R[509][8];				r_cell_reg[508] = inform_R[254][8];				r_cell_reg[509] = inform_R[510][8];				r_cell_reg[510] = inform_R[255][8];				r_cell_reg[511] = inform_R[511][8];				r_cell_reg[512] = inform_R[512][8];				r_cell_reg[513] = inform_R[768][8];				r_cell_reg[514] = inform_R[513][8];				r_cell_reg[515] = inform_R[769][8];				r_cell_reg[516] = inform_R[514][8];				r_cell_reg[517] = inform_R[770][8];				r_cell_reg[518] = inform_R[515][8];				r_cell_reg[519] = inform_R[771][8];				r_cell_reg[520] = inform_R[516][8];				r_cell_reg[521] = inform_R[772][8];				r_cell_reg[522] = inform_R[517][8];				r_cell_reg[523] = inform_R[773][8];				r_cell_reg[524] = inform_R[518][8];				r_cell_reg[525] = inform_R[774][8];				r_cell_reg[526] = inform_R[519][8];				r_cell_reg[527] = inform_R[775][8];				r_cell_reg[528] = inform_R[520][8];				r_cell_reg[529] = inform_R[776][8];				r_cell_reg[530] = inform_R[521][8];				r_cell_reg[531] = inform_R[777][8];				r_cell_reg[532] = inform_R[522][8];				r_cell_reg[533] = inform_R[778][8];				r_cell_reg[534] = inform_R[523][8];				r_cell_reg[535] = inform_R[779][8];				r_cell_reg[536] = inform_R[524][8];				r_cell_reg[537] = inform_R[780][8];				r_cell_reg[538] = inform_R[525][8];				r_cell_reg[539] = inform_R[781][8];				r_cell_reg[540] = inform_R[526][8];				r_cell_reg[541] = inform_R[782][8];				r_cell_reg[542] = inform_R[527][8];				r_cell_reg[543] = inform_R[783][8];				r_cell_reg[544] = inform_R[528][8];				r_cell_reg[545] = inform_R[784][8];				r_cell_reg[546] = inform_R[529][8];				r_cell_reg[547] = inform_R[785][8];				r_cell_reg[548] = inform_R[530][8];				r_cell_reg[549] = inform_R[786][8];				r_cell_reg[550] = inform_R[531][8];				r_cell_reg[551] = inform_R[787][8];				r_cell_reg[552] = inform_R[532][8];				r_cell_reg[553] = inform_R[788][8];				r_cell_reg[554] = inform_R[533][8];				r_cell_reg[555] = inform_R[789][8];				r_cell_reg[556] = inform_R[534][8];				r_cell_reg[557] = inform_R[790][8];				r_cell_reg[558] = inform_R[535][8];				r_cell_reg[559] = inform_R[791][8];				r_cell_reg[560] = inform_R[536][8];				r_cell_reg[561] = inform_R[792][8];				r_cell_reg[562] = inform_R[537][8];				r_cell_reg[563] = inform_R[793][8];				r_cell_reg[564] = inform_R[538][8];				r_cell_reg[565] = inform_R[794][8];				r_cell_reg[566] = inform_R[539][8];				r_cell_reg[567] = inform_R[795][8];				r_cell_reg[568] = inform_R[540][8];				r_cell_reg[569] = inform_R[796][8];				r_cell_reg[570] = inform_R[541][8];				r_cell_reg[571] = inform_R[797][8];				r_cell_reg[572] = inform_R[542][8];				r_cell_reg[573] = inform_R[798][8];				r_cell_reg[574] = inform_R[543][8];				r_cell_reg[575] = inform_R[799][8];				r_cell_reg[576] = inform_R[544][8];				r_cell_reg[577] = inform_R[800][8];				r_cell_reg[578] = inform_R[545][8];				r_cell_reg[579] = inform_R[801][8];				r_cell_reg[580] = inform_R[546][8];				r_cell_reg[581] = inform_R[802][8];				r_cell_reg[582] = inform_R[547][8];				r_cell_reg[583] = inform_R[803][8];				r_cell_reg[584] = inform_R[548][8];				r_cell_reg[585] = inform_R[804][8];				r_cell_reg[586] = inform_R[549][8];				r_cell_reg[587] = inform_R[805][8];				r_cell_reg[588] = inform_R[550][8];				r_cell_reg[589] = inform_R[806][8];				r_cell_reg[590] = inform_R[551][8];				r_cell_reg[591] = inform_R[807][8];				r_cell_reg[592] = inform_R[552][8];				r_cell_reg[593] = inform_R[808][8];				r_cell_reg[594] = inform_R[553][8];				r_cell_reg[595] = inform_R[809][8];				r_cell_reg[596] = inform_R[554][8];				r_cell_reg[597] = inform_R[810][8];				r_cell_reg[598] = inform_R[555][8];				r_cell_reg[599] = inform_R[811][8];				r_cell_reg[600] = inform_R[556][8];				r_cell_reg[601] = inform_R[812][8];				r_cell_reg[602] = inform_R[557][8];				r_cell_reg[603] = inform_R[813][8];				r_cell_reg[604] = inform_R[558][8];				r_cell_reg[605] = inform_R[814][8];				r_cell_reg[606] = inform_R[559][8];				r_cell_reg[607] = inform_R[815][8];				r_cell_reg[608] = inform_R[560][8];				r_cell_reg[609] = inform_R[816][8];				r_cell_reg[610] = inform_R[561][8];				r_cell_reg[611] = inform_R[817][8];				r_cell_reg[612] = inform_R[562][8];				r_cell_reg[613] = inform_R[818][8];				r_cell_reg[614] = inform_R[563][8];				r_cell_reg[615] = inform_R[819][8];				r_cell_reg[616] = inform_R[564][8];				r_cell_reg[617] = inform_R[820][8];				r_cell_reg[618] = inform_R[565][8];				r_cell_reg[619] = inform_R[821][8];				r_cell_reg[620] = inform_R[566][8];				r_cell_reg[621] = inform_R[822][8];				r_cell_reg[622] = inform_R[567][8];				r_cell_reg[623] = inform_R[823][8];				r_cell_reg[624] = inform_R[568][8];				r_cell_reg[625] = inform_R[824][8];				r_cell_reg[626] = inform_R[569][8];				r_cell_reg[627] = inform_R[825][8];				r_cell_reg[628] = inform_R[570][8];				r_cell_reg[629] = inform_R[826][8];				r_cell_reg[630] = inform_R[571][8];				r_cell_reg[631] = inform_R[827][8];				r_cell_reg[632] = inform_R[572][8];				r_cell_reg[633] = inform_R[828][8];				r_cell_reg[634] = inform_R[573][8];				r_cell_reg[635] = inform_R[829][8];				r_cell_reg[636] = inform_R[574][8];				r_cell_reg[637] = inform_R[830][8];				r_cell_reg[638] = inform_R[575][8];				r_cell_reg[639] = inform_R[831][8];				r_cell_reg[640] = inform_R[576][8];				r_cell_reg[641] = inform_R[832][8];				r_cell_reg[642] = inform_R[577][8];				r_cell_reg[643] = inform_R[833][8];				r_cell_reg[644] = inform_R[578][8];				r_cell_reg[645] = inform_R[834][8];				r_cell_reg[646] = inform_R[579][8];				r_cell_reg[647] = inform_R[835][8];				r_cell_reg[648] = inform_R[580][8];				r_cell_reg[649] = inform_R[836][8];				r_cell_reg[650] = inform_R[581][8];				r_cell_reg[651] = inform_R[837][8];				r_cell_reg[652] = inform_R[582][8];				r_cell_reg[653] = inform_R[838][8];				r_cell_reg[654] = inform_R[583][8];				r_cell_reg[655] = inform_R[839][8];				r_cell_reg[656] = inform_R[584][8];				r_cell_reg[657] = inform_R[840][8];				r_cell_reg[658] = inform_R[585][8];				r_cell_reg[659] = inform_R[841][8];				r_cell_reg[660] = inform_R[586][8];				r_cell_reg[661] = inform_R[842][8];				r_cell_reg[662] = inform_R[587][8];				r_cell_reg[663] = inform_R[843][8];				r_cell_reg[664] = inform_R[588][8];				r_cell_reg[665] = inform_R[844][8];				r_cell_reg[666] = inform_R[589][8];				r_cell_reg[667] = inform_R[845][8];				r_cell_reg[668] = inform_R[590][8];				r_cell_reg[669] = inform_R[846][8];				r_cell_reg[670] = inform_R[591][8];				r_cell_reg[671] = inform_R[847][8];				r_cell_reg[672] = inform_R[592][8];				r_cell_reg[673] = inform_R[848][8];				r_cell_reg[674] = inform_R[593][8];				r_cell_reg[675] = inform_R[849][8];				r_cell_reg[676] = inform_R[594][8];				r_cell_reg[677] = inform_R[850][8];				r_cell_reg[678] = inform_R[595][8];				r_cell_reg[679] = inform_R[851][8];				r_cell_reg[680] = inform_R[596][8];				r_cell_reg[681] = inform_R[852][8];				r_cell_reg[682] = inform_R[597][8];				r_cell_reg[683] = inform_R[853][8];				r_cell_reg[684] = inform_R[598][8];				r_cell_reg[685] = inform_R[854][8];				r_cell_reg[686] = inform_R[599][8];				r_cell_reg[687] = inform_R[855][8];				r_cell_reg[688] = inform_R[600][8];				r_cell_reg[689] = inform_R[856][8];				r_cell_reg[690] = inform_R[601][8];				r_cell_reg[691] = inform_R[857][8];				r_cell_reg[692] = inform_R[602][8];				r_cell_reg[693] = inform_R[858][8];				r_cell_reg[694] = inform_R[603][8];				r_cell_reg[695] = inform_R[859][8];				r_cell_reg[696] = inform_R[604][8];				r_cell_reg[697] = inform_R[860][8];				r_cell_reg[698] = inform_R[605][8];				r_cell_reg[699] = inform_R[861][8];				r_cell_reg[700] = inform_R[606][8];				r_cell_reg[701] = inform_R[862][8];				r_cell_reg[702] = inform_R[607][8];				r_cell_reg[703] = inform_R[863][8];				r_cell_reg[704] = inform_R[608][8];				r_cell_reg[705] = inform_R[864][8];				r_cell_reg[706] = inform_R[609][8];				r_cell_reg[707] = inform_R[865][8];				r_cell_reg[708] = inform_R[610][8];				r_cell_reg[709] = inform_R[866][8];				r_cell_reg[710] = inform_R[611][8];				r_cell_reg[711] = inform_R[867][8];				r_cell_reg[712] = inform_R[612][8];				r_cell_reg[713] = inform_R[868][8];				r_cell_reg[714] = inform_R[613][8];				r_cell_reg[715] = inform_R[869][8];				r_cell_reg[716] = inform_R[614][8];				r_cell_reg[717] = inform_R[870][8];				r_cell_reg[718] = inform_R[615][8];				r_cell_reg[719] = inform_R[871][8];				r_cell_reg[720] = inform_R[616][8];				r_cell_reg[721] = inform_R[872][8];				r_cell_reg[722] = inform_R[617][8];				r_cell_reg[723] = inform_R[873][8];				r_cell_reg[724] = inform_R[618][8];				r_cell_reg[725] = inform_R[874][8];				r_cell_reg[726] = inform_R[619][8];				r_cell_reg[727] = inform_R[875][8];				r_cell_reg[728] = inform_R[620][8];				r_cell_reg[729] = inform_R[876][8];				r_cell_reg[730] = inform_R[621][8];				r_cell_reg[731] = inform_R[877][8];				r_cell_reg[732] = inform_R[622][8];				r_cell_reg[733] = inform_R[878][8];				r_cell_reg[734] = inform_R[623][8];				r_cell_reg[735] = inform_R[879][8];				r_cell_reg[736] = inform_R[624][8];				r_cell_reg[737] = inform_R[880][8];				r_cell_reg[738] = inform_R[625][8];				r_cell_reg[739] = inform_R[881][8];				r_cell_reg[740] = inform_R[626][8];				r_cell_reg[741] = inform_R[882][8];				r_cell_reg[742] = inform_R[627][8];				r_cell_reg[743] = inform_R[883][8];				r_cell_reg[744] = inform_R[628][8];				r_cell_reg[745] = inform_R[884][8];				r_cell_reg[746] = inform_R[629][8];				r_cell_reg[747] = inform_R[885][8];				r_cell_reg[748] = inform_R[630][8];				r_cell_reg[749] = inform_R[886][8];				r_cell_reg[750] = inform_R[631][8];				r_cell_reg[751] = inform_R[887][8];				r_cell_reg[752] = inform_R[632][8];				r_cell_reg[753] = inform_R[888][8];				r_cell_reg[754] = inform_R[633][8];				r_cell_reg[755] = inform_R[889][8];				r_cell_reg[756] = inform_R[634][8];				r_cell_reg[757] = inform_R[890][8];				r_cell_reg[758] = inform_R[635][8];				r_cell_reg[759] = inform_R[891][8];				r_cell_reg[760] = inform_R[636][8];				r_cell_reg[761] = inform_R[892][8];				r_cell_reg[762] = inform_R[637][8];				r_cell_reg[763] = inform_R[893][8];				r_cell_reg[764] = inform_R[638][8];				r_cell_reg[765] = inform_R[894][8];				r_cell_reg[766] = inform_R[639][8];				r_cell_reg[767] = inform_R[895][8];				r_cell_reg[768] = inform_R[640][8];				r_cell_reg[769] = inform_R[896][8];				r_cell_reg[770] = inform_R[641][8];				r_cell_reg[771] = inform_R[897][8];				r_cell_reg[772] = inform_R[642][8];				r_cell_reg[773] = inform_R[898][8];				r_cell_reg[774] = inform_R[643][8];				r_cell_reg[775] = inform_R[899][8];				r_cell_reg[776] = inform_R[644][8];				r_cell_reg[777] = inform_R[900][8];				r_cell_reg[778] = inform_R[645][8];				r_cell_reg[779] = inform_R[901][8];				r_cell_reg[780] = inform_R[646][8];				r_cell_reg[781] = inform_R[902][8];				r_cell_reg[782] = inform_R[647][8];				r_cell_reg[783] = inform_R[903][8];				r_cell_reg[784] = inform_R[648][8];				r_cell_reg[785] = inform_R[904][8];				r_cell_reg[786] = inform_R[649][8];				r_cell_reg[787] = inform_R[905][8];				r_cell_reg[788] = inform_R[650][8];				r_cell_reg[789] = inform_R[906][8];				r_cell_reg[790] = inform_R[651][8];				r_cell_reg[791] = inform_R[907][8];				r_cell_reg[792] = inform_R[652][8];				r_cell_reg[793] = inform_R[908][8];				r_cell_reg[794] = inform_R[653][8];				r_cell_reg[795] = inform_R[909][8];				r_cell_reg[796] = inform_R[654][8];				r_cell_reg[797] = inform_R[910][8];				r_cell_reg[798] = inform_R[655][8];				r_cell_reg[799] = inform_R[911][8];				r_cell_reg[800] = inform_R[656][8];				r_cell_reg[801] = inform_R[912][8];				r_cell_reg[802] = inform_R[657][8];				r_cell_reg[803] = inform_R[913][8];				r_cell_reg[804] = inform_R[658][8];				r_cell_reg[805] = inform_R[914][8];				r_cell_reg[806] = inform_R[659][8];				r_cell_reg[807] = inform_R[915][8];				r_cell_reg[808] = inform_R[660][8];				r_cell_reg[809] = inform_R[916][8];				r_cell_reg[810] = inform_R[661][8];				r_cell_reg[811] = inform_R[917][8];				r_cell_reg[812] = inform_R[662][8];				r_cell_reg[813] = inform_R[918][8];				r_cell_reg[814] = inform_R[663][8];				r_cell_reg[815] = inform_R[919][8];				r_cell_reg[816] = inform_R[664][8];				r_cell_reg[817] = inform_R[920][8];				r_cell_reg[818] = inform_R[665][8];				r_cell_reg[819] = inform_R[921][8];				r_cell_reg[820] = inform_R[666][8];				r_cell_reg[821] = inform_R[922][8];				r_cell_reg[822] = inform_R[667][8];				r_cell_reg[823] = inform_R[923][8];				r_cell_reg[824] = inform_R[668][8];				r_cell_reg[825] = inform_R[924][8];				r_cell_reg[826] = inform_R[669][8];				r_cell_reg[827] = inform_R[925][8];				r_cell_reg[828] = inform_R[670][8];				r_cell_reg[829] = inform_R[926][8];				r_cell_reg[830] = inform_R[671][8];				r_cell_reg[831] = inform_R[927][8];				r_cell_reg[832] = inform_R[672][8];				r_cell_reg[833] = inform_R[928][8];				r_cell_reg[834] = inform_R[673][8];				r_cell_reg[835] = inform_R[929][8];				r_cell_reg[836] = inform_R[674][8];				r_cell_reg[837] = inform_R[930][8];				r_cell_reg[838] = inform_R[675][8];				r_cell_reg[839] = inform_R[931][8];				r_cell_reg[840] = inform_R[676][8];				r_cell_reg[841] = inform_R[932][8];				r_cell_reg[842] = inform_R[677][8];				r_cell_reg[843] = inform_R[933][8];				r_cell_reg[844] = inform_R[678][8];				r_cell_reg[845] = inform_R[934][8];				r_cell_reg[846] = inform_R[679][8];				r_cell_reg[847] = inform_R[935][8];				r_cell_reg[848] = inform_R[680][8];				r_cell_reg[849] = inform_R[936][8];				r_cell_reg[850] = inform_R[681][8];				r_cell_reg[851] = inform_R[937][8];				r_cell_reg[852] = inform_R[682][8];				r_cell_reg[853] = inform_R[938][8];				r_cell_reg[854] = inform_R[683][8];				r_cell_reg[855] = inform_R[939][8];				r_cell_reg[856] = inform_R[684][8];				r_cell_reg[857] = inform_R[940][8];				r_cell_reg[858] = inform_R[685][8];				r_cell_reg[859] = inform_R[941][8];				r_cell_reg[860] = inform_R[686][8];				r_cell_reg[861] = inform_R[942][8];				r_cell_reg[862] = inform_R[687][8];				r_cell_reg[863] = inform_R[943][8];				r_cell_reg[864] = inform_R[688][8];				r_cell_reg[865] = inform_R[944][8];				r_cell_reg[866] = inform_R[689][8];				r_cell_reg[867] = inform_R[945][8];				r_cell_reg[868] = inform_R[690][8];				r_cell_reg[869] = inform_R[946][8];				r_cell_reg[870] = inform_R[691][8];				r_cell_reg[871] = inform_R[947][8];				r_cell_reg[872] = inform_R[692][8];				r_cell_reg[873] = inform_R[948][8];				r_cell_reg[874] = inform_R[693][8];				r_cell_reg[875] = inform_R[949][8];				r_cell_reg[876] = inform_R[694][8];				r_cell_reg[877] = inform_R[950][8];				r_cell_reg[878] = inform_R[695][8];				r_cell_reg[879] = inform_R[951][8];				r_cell_reg[880] = inform_R[696][8];				r_cell_reg[881] = inform_R[952][8];				r_cell_reg[882] = inform_R[697][8];				r_cell_reg[883] = inform_R[953][8];				r_cell_reg[884] = inform_R[698][8];				r_cell_reg[885] = inform_R[954][8];				r_cell_reg[886] = inform_R[699][8];				r_cell_reg[887] = inform_R[955][8];				r_cell_reg[888] = inform_R[700][8];				r_cell_reg[889] = inform_R[956][8];				r_cell_reg[890] = inform_R[701][8];				r_cell_reg[891] = inform_R[957][8];				r_cell_reg[892] = inform_R[702][8];				r_cell_reg[893] = inform_R[958][8];				r_cell_reg[894] = inform_R[703][8];				r_cell_reg[895] = inform_R[959][8];				r_cell_reg[896] = inform_R[704][8];				r_cell_reg[897] = inform_R[960][8];				r_cell_reg[898] = inform_R[705][8];				r_cell_reg[899] = inform_R[961][8];				r_cell_reg[900] = inform_R[706][8];				r_cell_reg[901] = inform_R[962][8];				r_cell_reg[902] = inform_R[707][8];				r_cell_reg[903] = inform_R[963][8];				r_cell_reg[904] = inform_R[708][8];				r_cell_reg[905] = inform_R[964][8];				r_cell_reg[906] = inform_R[709][8];				r_cell_reg[907] = inform_R[965][8];				r_cell_reg[908] = inform_R[710][8];				r_cell_reg[909] = inform_R[966][8];				r_cell_reg[910] = inform_R[711][8];				r_cell_reg[911] = inform_R[967][8];				r_cell_reg[912] = inform_R[712][8];				r_cell_reg[913] = inform_R[968][8];				r_cell_reg[914] = inform_R[713][8];				r_cell_reg[915] = inform_R[969][8];				r_cell_reg[916] = inform_R[714][8];				r_cell_reg[917] = inform_R[970][8];				r_cell_reg[918] = inform_R[715][8];				r_cell_reg[919] = inform_R[971][8];				r_cell_reg[920] = inform_R[716][8];				r_cell_reg[921] = inform_R[972][8];				r_cell_reg[922] = inform_R[717][8];				r_cell_reg[923] = inform_R[973][8];				r_cell_reg[924] = inform_R[718][8];				r_cell_reg[925] = inform_R[974][8];				r_cell_reg[926] = inform_R[719][8];				r_cell_reg[927] = inform_R[975][8];				r_cell_reg[928] = inform_R[720][8];				r_cell_reg[929] = inform_R[976][8];				r_cell_reg[930] = inform_R[721][8];				r_cell_reg[931] = inform_R[977][8];				r_cell_reg[932] = inform_R[722][8];				r_cell_reg[933] = inform_R[978][8];				r_cell_reg[934] = inform_R[723][8];				r_cell_reg[935] = inform_R[979][8];				r_cell_reg[936] = inform_R[724][8];				r_cell_reg[937] = inform_R[980][8];				r_cell_reg[938] = inform_R[725][8];				r_cell_reg[939] = inform_R[981][8];				r_cell_reg[940] = inform_R[726][8];				r_cell_reg[941] = inform_R[982][8];				r_cell_reg[942] = inform_R[727][8];				r_cell_reg[943] = inform_R[983][8];				r_cell_reg[944] = inform_R[728][8];				r_cell_reg[945] = inform_R[984][8];				r_cell_reg[946] = inform_R[729][8];				r_cell_reg[947] = inform_R[985][8];				r_cell_reg[948] = inform_R[730][8];				r_cell_reg[949] = inform_R[986][8];				r_cell_reg[950] = inform_R[731][8];				r_cell_reg[951] = inform_R[987][8];				r_cell_reg[952] = inform_R[732][8];				r_cell_reg[953] = inform_R[988][8];				r_cell_reg[954] = inform_R[733][8];				r_cell_reg[955] = inform_R[989][8];				r_cell_reg[956] = inform_R[734][8];				r_cell_reg[957] = inform_R[990][8];				r_cell_reg[958] = inform_R[735][8];				r_cell_reg[959] = inform_R[991][8];				r_cell_reg[960] = inform_R[736][8];				r_cell_reg[961] = inform_R[992][8];				r_cell_reg[962] = inform_R[737][8];				r_cell_reg[963] = inform_R[993][8];				r_cell_reg[964] = inform_R[738][8];				r_cell_reg[965] = inform_R[994][8];				r_cell_reg[966] = inform_R[739][8];				r_cell_reg[967] = inform_R[995][8];				r_cell_reg[968] = inform_R[740][8];				r_cell_reg[969] = inform_R[996][8];				r_cell_reg[970] = inform_R[741][8];				r_cell_reg[971] = inform_R[997][8];				r_cell_reg[972] = inform_R[742][8];				r_cell_reg[973] = inform_R[998][8];				r_cell_reg[974] = inform_R[743][8];				r_cell_reg[975] = inform_R[999][8];				r_cell_reg[976] = inform_R[744][8];				r_cell_reg[977] = inform_R[1000][8];				r_cell_reg[978] = inform_R[745][8];				r_cell_reg[979] = inform_R[1001][8];				r_cell_reg[980] = inform_R[746][8];				r_cell_reg[981] = inform_R[1002][8];				r_cell_reg[982] = inform_R[747][8];				r_cell_reg[983] = inform_R[1003][8];				r_cell_reg[984] = inform_R[748][8];				r_cell_reg[985] = inform_R[1004][8];				r_cell_reg[986] = inform_R[749][8];				r_cell_reg[987] = inform_R[1005][8];				r_cell_reg[988] = inform_R[750][8];				r_cell_reg[989] = inform_R[1006][8];				r_cell_reg[990] = inform_R[751][8];				r_cell_reg[991] = inform_R[1007][8];				r_cell_reg[992] = inform_R[752][8];				r_cell_reg[993] = inform_R[1008][8];				r_cell_reg[994] = inform_R[753][8];				r_cell_reg[995] = inform_R[1009][8];				r_cell_reg[996] = inform_R[754][8];				r_cell_reg[997] = inform_R[1010][8];				r_cell_reg[998] = inform_R[755][8];				r_cell_reg[999] = inform_R[1011][8];				r_cell_reg[1000] = inform_R[756][8];				r_cell_reg[1001] = inform_R[1012][8];				r_cell_reg[1002] = inform_R[757][8];				r_cell_reg[1003] = inform_R[1013][8];				r_cell_reg[1004] = inform_R[758][8];				r_cell_reg[1005] = inform_R[1014][8];				r_cell_reg[1006] = inform_R[759][8];				r_cell_reg[1007] = inform_R[1015][8];				r_cell_reg[1008] = inform_R[760][8];				r_cell_reg[1009] = inform_R[1016][8];				r_cell_reg[1010] = inform_R[761][8];				r_cell_reg[1011] = inform_R[1017][8];				r_cell_reg[1012] = inform_R[762][8];				r_cell_reg[1013] = inform_R[1018][8];				r_cell_reg[1014] = inform_R[763][8];				r_cell_reg[1015] = inform_R[1019][8];				r_cell_reg[1016] = inform_R[764][8];				r_cell_reg[1017] = inform_R[1020][8];				r_cell_reg[1018] = inform_R[765][8];				r_cell_reg[1019] = inform_R[1021][8];				r_cell_reg[1020] = inform_R[766][8];				r_cell_reg[1021] = inform_R[1022][8];				r_cell_reg[1022] = inform_R[767][8];				r_cell_reg[1023] = inform_R[1023][8];				l_cell_reg[0] = inform_L[0][9];				l_cell_reg[1] = inform_L[256][9];				l_cell_reg[2] = inform_L[1][9];				l_cell_reg[3] = inform_L[257][9];				l_cell_reg[4] = inform_L[2][9];				l_cell_reg[5] = inform_L[258][9];				l_cell_reg[6] = inform_L[3][9];				l_cell_reg[7] = inform_L[259][9];				l_cell_reg[8] = inform_L[4][9];				l_cell_reg[9] = inform_L[260][9];				l_cell_reg[10] = inform_L[5][9];				l_cell_reg[11] = inform_L[261][9];				l_cell_reg[12] = inform_L[6][9];				l_cell_reg[13] = inform_L[262][9];				l_cell_reg[14] = inform_L[7][9];				l_cell_reg[15] = inform_L[263][9];				l_cell_reg[16] = inform_L[8][9];				l_cell_reg[17] = inform_L[264][9];				l_cell_reg[18] = inform_L[9][9];				l_cell_reg[19] = inform_L[265][9];				l_cell_reg[20] = inform_L[10][9];				l_cell_reg[21] = inform_L[266][9];				l_cell_reg[22] = inform_L[11][9];				l_cell_reg[23] = inform_L[267][9];				l_cell_reg[24] = inform_L[12][9];				l_cell_reg[25] = inform_L[268][9];				l_cell_reg[26] = inform_L[13][9];				l_cell_reg[27] = inform_L[269][9];				l_cell_reg[28] = inform_L[14][9];				l_cell_reg[29] = inform_L[270][9];				l_cell_reg[30] = inform_L[15][9];				l_cell_reg[31] = inform_L[271][9];				l_cell_reg[32] = inform_L[16][9];				l_cell_reg[33] = inform_L[272][9];				l_cell_reg[34] = inform_L[17][9];				l_cell_reg[35] = inform_L[273][9];				l_cell_reg[36] = inform_L[18][9];				l_cell_reg[37] = inform_L[274][9];				l_cell_reg[38] = inform_L[19][9];				l_cell_reg[39] = inform_L[275][9];				l_cell_reg[40] = inform_L[20][9];				l_cell_reg[41] = inform_L[276][9];				l_cell_reg[42] = inform_L[21][9];				l_cell_reg[43] = inform_L[277][9];				l_cell_reg[44] = inform_L[22][9];				l_cell_reg[45] = inform_L[278][9];				l_cell_reg[46] = inform_L[23][9];				l_cell_reg[47] = inform_L[279][9];				l_cell_reg[48] = inform_L[24][9];				l_cell_reg[49] = inform_L[280][9];				l_cell_reg[50] = inform_L[25][9];				l_cell_reg[51] = inform_L[281][9];				l_cell_reg[52] = inform_L[26][9];				l_cell_reg[53] = inform_L[282][9];				l_cell_reg[54] = inform_L[27][9];				l_cell_reg[55] = inform_L[283][9];				l_cell_reg[56] = inform_L[28][9];				l_cell_reg[57] = inform_L[284][9];				l_cell_reg[58] = inform_L[29][9];				l_cell_reg[59] = inform_L[285][9];				l_cell_reg[60] = inform_L[30][9];				l_cell_reg[61] = inform_L[286][9];				l_cell_reg[62] = inform_L[31][9];				l_cell_reg[63] = inform_L[287][9];				l_cell_reg[64] = inform_L[32][9];				l_cell_reg[65] = inform_L[288][9];				l_cell_reg[66] = inform_L[33][9];				l_cell_reg[67] = inform_L[289][9];				l_cell_reg[68] = inform_L[34][9];				l_cell_reg[69] = inform_L[290][9];				l_cell_reg[70] = inform_L[35][9];				l_cell_reg[71] = inform_L[291][9];				l_cell_reg[72] = inform_L[36][9];				l_cell_reg[73] = inform_L[292][9];				l_cell_reg[74] = inform_L[37][9];				l_cell_reg[75] = inform_L[293][9];				l_cell_reg[76] = inform_L[38][9];				l_cell_reg[77] = inform_L[294][9];				l_cell_reg[78] = inform_L[39][9];				l_cell_reg[79] = inform_L[295][9];				l_cell_reg[80] = inform_L[40][9];				l_cell_reg[81] = inform_L[296][9];				l_cell_reg[82] = inform_L[41][9];				l_cell_reg[83] = inform_L[297][9];				l_cell_reg[84] = inform_L[42][9];				l_cell_reg[85] = inform_L[298][9];				l_cell_reg[86] = inform_L[43][9];				l_cell_reg[87] = inform_L[299][9];				l_cell_reg[88] = inform_L[44][9];				l_cell_reg[89] = inform_L[300][9];				l_cell_reg[90] = inform_L[45][9];				l_cell_reg[91] = inform_L[301][9];				l_cell_reg[92] = inform_L[46][9];				l_cell_reg[93] = inform_L[302][9];				l_cell_reg[94] = inform_L[47][9];				l_cell_reg[95] = inform_L[303][9];				l_cell_reg[96] = inform_L[48][9];				l_cell_reg[97] = inform_L[304][9];				l_cell_reg[98] = inform_L[49][9];				l_cell_reg[99] = inform_L[305][9];				l_cell_reg[100] = inform_L[50][9];				l_cell_reg[101] = inform_L[306][9];				l_cell_reg[102] = inform_L[51][9];				l_cell_reg[103] = inform_L[307][9];				l_cell_reg[104] = inform_L[52][9];				l_cell_reg[105] = inform_L[308][9];				l_cell_reg[106] = inform_L[53][9];				l_cell_reg[107] = inform_L[309][9];				l_cell_reg[108] = inform_L[54][9];				l_cell_reg[109] = inform_L[310][9];				l_cell_reg[110] = inform_L[55][9];				l_cell_reg[111] = inform_L[311][9];				l_cell_reg[112] = inform_L[56][9];				l_cell_reg[113] = inform_L[312][9];				l_cell_reg[114] = inform_L[57][9];				l_cell_reg[115] = inform_L[313][9];				l_cell_reg[116] = inform_L[58][9];				l_cell_reg[117] = inform_L[314][9];				l_cell_reg[118] = inform_L[59][9];				l_cell_reg[119] = inform_L[315][9];				l_cell_reg[120] = inform_L[60][9];				l_cell_reg[121] = inform_L[316][9];				l_cell_reg[122] = inform_L[61][9];				l_cell_reg[123] = inform_L[317][9];				l_cell_reg[124] = inform_L[62][9];				l_cell_reg[125] = inform_L[318][9];				l_cell_reg[126] = inform_L[63][9];				l_cell_reg[127] = inform_L[319][9];				l_cell_reg[128] = inform_L[64][9];				l_cell_reg[129] = inform_L[320][9];				l_cell_reg[130] = inform_L[65][9];				l_cell_reg[131] = inform_L[321][9];				l_cell_reg[132] = inform_L[66][9];				l_cell_reg[133] = inform_L[322][9];				l_cell_reg[134] = inform_L[67][9];				l_cell_reg[135] = inform_L[323][9];				l_cell_reg[136] = inform_L[68][9];				l_cell_reg[137] = inform_L[324][9];				l_cell_reg[138] = inform_L[69][9];				l_cell_reg[139] = inform_L[325][9];				l_cell_reg[140] = inform_L[70][9];				l_cell_reg[141] = inform_L[326][9];				l_cell_reg[142] = inform_L[71][9];				l_cell_reg[143] = inform_L[327][9];				l_cell_reg[144] = inform_L[72][9];				l_cell_reg[145] = inform_L[328][9];				l_cell_reg[146] = inform_L[73][9];				l_cell_reg[147] = inform_L[329][9];				l_cell_reg[148] = inform_L[74][9];				l_cell_reg[149] = inform_L[330][9];				l_cell_reg[150] = inform_L[75][9];				l_cell_reg[151] = inform_L[331][9];				l_cell_reg[152] = inform_L[76][9];				l_cell_reg[153] = inform_L[332][9];				l_cell_reg[154] = inform_L[77][9];				l_cell_reg[155] = inform_L[333][9];				l_cell_reg[156] = inform_L[78][9];				l_cell_reg[157] = inform_L[334][9];				l_cell_reg[158] = inform_L[79][9];				l_cell_reg[159] = inform_L[335][9];				l_cell_reg[160] = inform_L[80][9];				l_cell_reg[161] = inform_L[336][9];				l_cell_reg[162] = inform_L[81][9];				l_cell_reg[163] = inform_L[337][9];				l_cell_reg[164] = inform_L[82][9];				l_cell_reg[165] = inform_L[338][9];				l_cell_reg[166] = inform_L[83][9];				l_cell_reg[167] = inform_L[339][9];				l_cell_reg[168] = inform_L[84][9];				l_cell_reg[169] = inform_L[340][9];				l_cell_reg[170] = inform_L[85][9];				l_cell_reg[171] = inform_L[341][9];				l_cell_reg[172] = inform_L[86][9];				l_cell_reg[173] = inform_L[342][9];				l_cell_reg[174] = inform_L[87][9];				l_cell_reg[175] = inform_L[343][9];				l_cell_reg[176] = inform_L[88][9];				l_cell_reg[177] = inform_L[344][9];				l_cell_reg[178] = inform_L[89][9];				l_cell_reg[179] = inform_L[345][9];				l_cell_reg[180] = inform_L[90][9];				l_cell_reg[181] = inform_L[346][9];				l_cell_reg[182] = inform_L[91][9];				l_cell_reg[183] = inform_L[347][9];				l_cell_reg[184] = inform_L[92][9];				l_cell_reg[185] = inform_L[348][9];				l_cell_reg[186] = inform_L[93][9];				l_cell_reg[187] = inform_L[349][9];				l_cell_reg[188] = inform_L[94][9];				l_cell_reg[189] = inform_L[350][9];				l_cell_reg[190] = inform_L[95][9];				l_cell_reg[191] = inform_L[351][9];				l_cell_reg[192] = inform_L[96][9];				l_cell_reg[193] = inform_L[352][9];				l_cell_reg[194] = inform_L[97][9];				l_cell_reg[195] = inform_L[353][9];				l_cell_reg[196] = inform_L[98][9];				l_cell_reg[197] = inform_L[354][9];				l_cell_reg[198] = inform_L[99][9];				l_cell_reg[199] = inform_L[355][9];				l_cell_reg[200] = inform_L[100][9];				l_cell_reg[201] = inform_L[356][9];				l_cell_reg[202] = inform_L[101][9];				l_cell_reg[203] = inform_L[357][9];				l_cell_reg[204] = inform_L[102][9];				l_cell_reg[205] = inform_L[358][9];				l_cell_reg[206] = inform_L[103][9];				l_cell_reg[207] = inform_L[359][9];				l_cell_reg[208] = inform_L[104][9];				l_cell_reg[209] = inform_L[360][9];				l_cell_reg[210] = inform_L[105][9];				l_cell_reg[211] = inform_L[361][9];				l_cell_reg[212] = inform_L[106][9];				l_cell_reg[213] = inform_L[362][9];				l_cell_reg[214] = inform_L[107][9];				l_cell_reg[215] = inform_L[363][9];				l_cell_reg[216] = inform_L[108][9];				l_cell_reg[217] = inform_L[364][9];				l_cell_reg[218] = inform_L[109][9];				l_cell_reg[219] = inform_L[365][9];				l_cell_reg[220] = inform_L[110][9];				l_cell_reg[221] = inform_L[366][9];				l_cell_reg[222] = inform_L[111][9];				l_cell_reg[223] = inform_L[367][9];				l_cell_reg[224] = inform_L[112][9];				l_cell_reg[225] = inform_L[368][9];				l_cell_reg[226] = inform_L[113][9];				l_cell_reg[227] = inform_L[369][9];				l_cell_reg[228] = inform_L[114][9];				l_cell_reg[229] = inform_L[370][9];				l_cell_reg[230] = inform_L[115][9];				l_cell_reg[231] = inform_L[371][9];				l_cell_reg[232] = inform_L[116][9];				l_cell_reg[233] = inform_L[372][9];				l_cell_reg[234] = inform_L[117][9];				l_cell_reg[235] = inform_L[373][9];				l_cell_reg[236] = inform_L[118][9];				l_cell_reg[237] = inform_L[374][9];				l_cell_reg[238] = inform_L[119][9];				l_cell_reg[239] = inform_L[375][9];				l_cell_reg[240] = inform_L[120][9];				l_cell_reg[241] = inform_L[376][9];				l_cell_reg[242] = inform_L[121][9];				l_cell_reg[243] = inform_L[377][9];				l_cell_reg[244] = inform_L[122][9];				l_cell_reg[245] = inform_L[378][9];				l_cell_reg[246] = inform_L[123][9];				l_cell_reg[247] = inform_L[379][9];				l_cell_reg[248] = inform_L[124][9];				l_cell_reg[249] = inform_L[380][9];				l_cell_reg[250] = inform_L[125][9];				l_cell_reg[251] = inform_L[381][9];				l_cell_reg[252] = inform_L[126][9];				l_cell_reg[253] = inform_L[382][9];				l_cell_reg[254] = inform_L[127][9];				l_cell_reg[255] = inform_L[383][9];				l_cell_reg[256] = inform_L[128][9];				l_cell_reg[257] = inform_L[384][9];				l_cell_reg[258] = inform_L[129][9];				l_cell_reg[259] = inform_L[385][9];				l_cell_reg[260] = inform_L[130][9];				l_cell_reg[261] = inform_L[386][9];				l_cell_reg[262] = inform_L[131][9];				l_cell_reg[263] = inform_L[387][9];				l_cell_reg[264] = inform_L[132][9];				l_cell_reg[265] = inform_L[388][9];				l_cell_reg[266] = inform_L[133][9];				l_cell_reg[267] = inform_L[389][9];				l_cell_reg[268] = inform_L[134][9];				l_cell_reg[269] = inform_L[390][9];				l_cell_reg[270] = inform_L[135][9];				l_cell_reg[271] = inform_L[391][9];				l_cell_reg[272] = inform_L[136][9];				l_cell_reg[273] = inform_L[392][9];				l_cell_reg[274] = inform_L[137][9];				l_cell_reg[275] = inform_L[393][9];				l_cell_reg[276] = inform_L[138][9];				l_cell_reg[277] = inform_L[394][9];				l_cell_reg[278] = inform_L[139][9];				l_cell_reg[279] = inform_L[395][9];				l_cell_reg[280] = inform_L[140][9];				l_cell_reg[281] = inform_L[396][9];				l_cell_reg[282] = inform_L[141][9];				l_cell_reg[283] = inform_L[397][9];				l_cell_reg[284] = inform_L[142][9];				l_cell_reg[285] = inform_L[398][9];				l_cell_reg[286] = inform_L[143][9];				l_cell_reg[287] = inform_L[399][9];				l_cell_reg[288] = inform_L[144][9];				l_cell_reg[289] = inform_L[400][9];				l_cell_reg[290] = inform_L[145][9];				l_cell_reg[291] = inform_L[401][9];				l_cell_reg[292] = inform_L[146][9];				l_cell_reg[293] = inform_L[402][9];				l_cell_reg[294] = inform_L[147][9];				l_cell_reg[295] = inform_L[403][9];				l_cell_reg[296] = inform_L[148][9];				l_cell_reg[297] = inform_L[404][9];				l_cell_reg[298] = inform_L[149][9];				l_cell_reg[299] = inform_L[405][9];				l_cell_reg[300] = inform_L[150][9];				l_cell_reg[301] = inform_L[406][9];				l_cell_reg[302] = inform_L[151][9];				l_cell_reg[303] = inform_L[407][9];				l_cell_reg[304] = inform_L[152][9];				l_cell_reg[305] = inform_L[408][9];				l_cell_reg[306] = inform_L[153][9];				l_cell_reg[307] = inform_L[409][9];				l_cell_reg[308] = inform_L[154][9];				l_cell_reg[309] = inform_L[410][9];				l_cell_reg[310] = inform_L[155][9];				l_cell_reg[311] = inform_L[411][9];				l_cell_reg[312] = inform_L[156][9];				l_cell_reg[313] = inform_L[412][9];				l_cell_reg[314] = inform_L[157][9];				l_cell_reg[315] = inform_L[413][9];				l_cell_reg[316] = inform_L[158][9];				l_cell_reg[317] = inform_L[414][9];				l_cell_reg[318] = inform_L[159][9];				l_cell_reg[319] = inform_L[415][9];				l_cell_reg[320] = inform_L[160][9];				l_cell_reg[321] = inform_L[416][9];				l_cell_reg[322] = inform_L[161][9];				l_cell_reg[323] = inform_L[417][9];				l_cell_reg[324] = inform_L[162][9];				l_cell_reg[325] = inform_L[418][9];				l_cell_reg[326] = inform_L[163][9];				l_cell_reg[327] = inform_L[419][9];				l_cell_reg[328] = inform_L[164][9];				l_cell_reg[329] = inform_L[420][9];				l_cell_reg[330] = inform_L[165][9];				l_cell_reg[331] = inform_L[421][9];				l_cell_reg[332] = inform_L[166][9];				l_cell_reg[333] = inform_L[422][9];				l_cell_reg[334] = inform_L[167][9];				l_cell_reg[335] = inform_L[423][9];				l_cell_reg[336] = inform_L[168][9];				l_cell_reg[337] = inform_L[424][9];				l_cell_reg[338] = inform_L[169][9];				l_cell_reg[339] = inform_L[425][9];				l_cell_reg[340] = inform_L[170][9];				l_cell_reg[341] = inform_L[426][9];				l_cell_reg[342] = inform_L[171][9];				l_cell_reg[343] = inform_L[427][9];				l_cell_reg[344] = inform_L[172][9];				l_cell_reg[345] = inform_L[428][9];				l_cell_reg[346] = inform_L[173][9];				l_cell_reg[347] = inform_L[429][9];				l_cell_reg[348] = inform_L[174][9];				l_cell_reg[349] = inform_L[430][9];				l_cell_reg[350] = inform_L[175][9];				l_cell_reg[351] = inform_L[431][9];				l_cell_reg[352] = inform_L[176][9];				l_cell_reg[353] = inform_L[432][9];				l_cell_reg[354] = inform_L[177][9];				l_cell_reg[355] = inform_L[433][9];				l_cell_reg[356] = inform_L[178][9];				l_cell_reg[357] = inform_L[434][9];				l_cell_reg[358] = inform_L[179][9];				l_cell_reg[359] = inform_L[435][9];				l_cell_reg[360] = inform_L[180][9];				l_cell_reg[361] = inform_L[436][9];				l_cell_reg[362] = inform_L[181][9];				l_cell_reg[363] = inform_L[437][9];				l_cell_reg[364] = inform_L[182][9];				l_cell_reg[365] = inform_L[438][9];				l_cell_reg[366] = inform_L[183][9];				l_cell_reg[367] = inform_L[439][9];				l_cell_reg[368] = inform_L[184][9];				l_cell_reg[369] = inform_L[440][9];				l_cell_reg[370] = inform_L[185][9];				l_cell_reg[371] = inform_L[441][9];				l_cell_reg[372] = inform_L[186][9];				l_cell_reg[373] = inform_L[442][9];				l_cell_reg[374] = inform_L[187][9];				l_cell_reg[375] = inform_L[443][9];				l_cell_reg[376] = inform_L[188][9];				l_cell_reg[377] = inform_L[444][9];				l_cell_reg[378] = inform_L[189][9];				l_cell_reg[379] = inform_L[445][9];				l_cell_reg[380] = inform_L[190][9];				l_cell_reg[381] = inform_L[446][9];				l_cell_reg[382] = inform_L[191][9];				l_cell_reg[383] = inform_L[447][9];				l_cell_reg[384] = inform_L[192][9];				l_cell_reg[385] = inform_L[448][9];				l_cell_reg[386] = inform_L[193][9];				l_cell_reg[387] = inform_L[449][9];				l_cell_reg[388] = inform_L[194][9];				l_cell_reg[389] = inform_L[450][9];				l_cell_reg[390] = inform_L[195][9];				l_cell_reg[391] = inform_L[451][9];				l_cell_reg[392] = inform_L[196][9];				l_cell_reg[393] = inform_L[452][9];				l_cell_reg[394] = inform_L[197][9];				l_cell_reg[395] = inform_L[453][9];				l_cell_reg[396] = inform_L[198][9];				l_cell_reg[397] = inform_L[454][9];				l_cell_reg[398] = inform_L[199][9];				l_cell_reg[399] = inform_L[455][9];				l_cell_reg[400] = inform_L[200][9];				l_cell_reg[401] = inform_L[456][9];				l_cell_reg[402] = inform_L[201][9];				l_cell_reg[403] = inform_L[457][9];				l_cell_reg[404] = inform_L[202][9];				l_cell_reg[405] = inform_L[458][9];				l_cell_reg[406] = inform_L[203][9];				l_cell_reg[407] = inform_L[459][9];				l_cell_reg[408] = inform_L[204][9];				l_cell_reg[409] = inform_L[460][9];				l_cell_reg[410] = inform_L[205][9];				l_cell_reg[411] = inform_L[461][9];				l_cell_reg[412] = inform_L[206][9];				l_cell_reg[413] = inform_L[462][9];				l_cell_reg[414] = inform_L[207][9];				l_cell_reg[415] = inform_L[463][9];				l_cell_reg[416] = inform_L[208][9];				l_cell_reg[417] = inform_L[464][9];				l_cell_reg[418] = inform_L[209][9];				l_cell_reg[419] = inform_L[465][9];				l_cell_reg[420] = inform_L[210][9];				l_cell_reg[421] = inform_L[466][9];				l_cell_reg[422] = inform_L[211][9];				l_cell_reg[423] = inform_L[467][9];				l_cell_reg[424] = inform_L[212][9];				l_cell_reg[425] = inform_L[468][9];				l_cell_reg[426] = inform_L[213][9];				l_cell_reg[427] = inform_L[469][9];				l_cell_reg[428] = inform_L[214][9];				l_cell_reg[429] = inform_L[470][9];				l_cell_reg[430] = inform_L[215][9];				l_cell_reg[431] = inform_L[471][9];				l_cell_reg[432] = inform_L[216][9];				l_cell_reg[433] = inform_L[472][9];				l_cell_reg[434] = inform_L[217][9];				l_cell_reg[435] = inform_L[473][9];				l_cell_reg[436] = inform_L[218][9];				l_cell_reg[437] = inform_L[474][9];				l_cell_reg[438] = inform_L[219][9];				l_cell_reg[439] = inform_L[475][9];				l_cell_reg[440] = inform_L[220][9];				l_cell_reg[441] = inform_L[476][9];				l_cell_reg[442] = inform_L[221][9];				l_cell_reg[443] = inform_L[477][9];				l_cell_reg[444] = inform_L[222][9];				l_cell_reg[445] = inform_L[478][9];				l_cell_reg[446] = inform_L[223][9];				l_cell_reg[447] = inform_L[479][9];				l_cell_reg[448] = inform_L[224][9];				l_cell_reg[449] = inform_L[480][9];				l_cell_reg[450] = inform_L[225][9];				l_cell_reg[451] = inform_L[481][9];				l_cell_reg[452] = inform_L[226][9];				l_cell_reg[453] = inform_L[482][9];				l_cell_reg[454] = inform_L[227][9];				l_cell_reg[455] = inform_L[483][9];				l_cell_reg[456] = inform_L[228][9];				l_cell_reg[457] = inform_L[484][9];				l_cell_reg[458] = inform_L[229][9];				l_cell_reg[459] = inform_L[485][9];				l_cell_reg[460] = inform_L[230][9];				l_cell_reg[461] = inform_L[486][9];				l_cell_reg[462] = inform_L[231][9];				l_cell_reg[463] = inform_L[487][9];				l_cell_reg[464] = inform_L[232][9];				l_cell_reg[465] = inform_L[488][9];				l_cell_reg[466] = inform_L[233][9];				l_cell_reg[467] = inform_L[489][9];				l_cell_reg[468] = inform_L[234][9];				l_cell_reg[469] = inform_L[490][9];				l_cell_reg[470] = inform_L[235][9];				l_cell_reg[471] = inform_L[491][9];				l_cell_reg[472] = inform_L[236][9];				l_cell_reg[473] = inform_L[492][9];				l_cell_reg[474] = inform_L[237][9];				l_cell_reg[475] = inform_L[493][9];				l_cell_reg[476] = inform_L[238][9];				l_cell_reg[477] = inform_L[494][9];				l_cell_reg[478] = inform_L[239][9];				l_cell_reg[479] = inform_L[495][9];				l_cell_reg[480] = inform_L[240][9];				l_cell_reg[481] = inform_L[496][9];				l_cell_reg[482] = inform_L[241][9];				l_cell_reg[483] = inform_L[497][9];				l_cell_reg[484] = inform_L[242][9];				l_cell_reg[485] = inform_L[498][9];				l_cell_reg[486] = inform_L[243][9];				l_cell_reg[487] = inform_L[499][9];				l_cell_reg[488] = inform_L[244][9];				l_cell_reg[489] = inform_L[500][9];				l_cell_reg[490] = inform_L[245][9];				l_cell_reg[491] = inform_L[501][9];				l_cell_reg[492] = inform_L[246][9];				l_cell_reg[493] = inform_L[502][9];				l_cell_reg[494] = inform_L[247][9];				l_cell_reg[495] = inform_L[503][9];				l_cell_reg[496] = inform_L[248][9];				l_cell_reg[497] = inform_L[504][9];				l_cell_reg[498] = inform_L[249][9];				l_cell_reg[499] = inform_L[505][9];				l_cell_reg[500] = inform_L[250][9];				l_cell_reg[501] = inform_L[506][9];				l_cell_reg[502] = inform_L[251][9];				l_cell_reg[503] = inform_L[507][9];				l_cell_reg[504] = inform_L[252][9];				l_cell_reg[505] = inform_L[508][9];				l_cell_reg[506] = inform_L[253][9];				l_cell_reg[507] = inform_L[509][9];				l_cell_reg[508] = inform_L[254][9];				l_cell_reg[509] = inform_L[510][9];				l_cell_reg[510] = inform_L[255][9];				l_cell_reg[511] = inform_L[511][9];				l_cell_reg[512] = inform_L[512][9];				l_cell_reg[513] = inform_L[768][9];				l_cell_reg[514] = inform_L[513][9];				l_cell_reg[515] = inform_L[769][9];				l_cell_reg[516] = inform_L[514][9];				l_cell_reg[517] = inform_L[770][9];				l_cell_reg[518] = inform_L[515][9];				l_cell_reg[519] = inform_L[771][9];				l_cell_reg[520] = inform_L[516][9];				l_cell_reg[521] = inform_L[772][9];				l_cell_reg[522] = inform_L[517][9];				l_cell_reg[523] = inform_L[773][9];				l_cell_reg[524] = inform_L[518][9];				l_cell_reg[525] = inform_L[774][9];				l_cell_reg[526] = inform_L[519][9];				l_cell_reg[527] = inform_L[775][9];				l_cell_reg[528] = inform_L[520][9];				l_cell_reg[529] = inform_L[776][9];				l_cell_reg[530] = inform_L[521][9];				l_cell_reg[531] = inform_L[777][9];				l_cell_reg[532] = inform_L[522][9];				l_cell_reg[533] = inform_L[778][9];				l_cell_reg[534] = inform_L[523][9];				l_cell_reg[535] = inform_L[779][9];				l_cell_reg[536] = inform_L[524][9];				l_cell_reg[537] = inform_L[780][9];				l_cell_reg[538] = inform_L[525][9];				l_cell_reg[539] = inform_L[781][9];				l_cell_reg[540] = inform_L[526][9];				l_cell_reg[541] = inform_L[782][9];				l_cell_reg[542] = inform_L[527][9];				l_cell_reg[543] = inform_L[783][9];				l_cell_reg[544] = inform_L[528][9];				l_cell_reg[545] = inform_L[784][9];				l_cell_reg[546] = inform_L[529][9];				l_cell_reg[547] = inform_L[785][9];				l_cell_reg[548] = inform_L[530][9];				l_cell_reg[549] = inform_L[786][9];				l_cell_reg[550] = inform_L[531][9];				l_cell_reg[551] = inform_L[787][9];				l_cell_reg[552] = inform_L[532][9];				l_cell_reg[553] = inform_L[788][9];				l_cell_reg[554] = inform_L[533][9];				l_cell_reg[555] = inform_L[789][9];				l_cell_reg[556] = inform_L[534][9];				l_cell_reg[557] = inform_L[790][9];				l_cell_reg[558] = inform_L[535][9];				l_cell_reg[559] = inform_L[791][9];				l_cell_reg[560] = inform_L[536][9];				l_cell_reg[561] = inform_L[792][9];				l_cell_reg[562] = inform_L[537][9];				l_cell_reg[563] = inform_L[793][9];				l_cell_reg[564] = inform_L[538][9];				l_cell_reg[565] = inform_L[794][9];				l_cell_reg[566] = inform_L[539][9];				l_cell_reg[567] = inform_L[795][9];				l_cell_reg[568] = inform_L[540][9];				l_cell_reg[569] = inform_L[796][9];				l_cell_reg[570] = inform_L[541][9];				l_cell_reg[571] = inform_L[797][9];				l_cell_reg[572] = inform_L[542][9];				l_cell_reg[573] = inform_L[798][9];				l_cell_reg[574] = inform_L[543][9];				l_cell_reg[575] = inform_L[799][9];				l_cell_reg[576] = inform_L[544][9];				l_cell_reg[577] = inform_L[800][9];				l_cell_reg[578] = inform_L[545][9];				l_cell_reg[579] = inform_L[801][9];				l_cell_reg[580] = inform_L[546][9];				l_cell_reg[581] = inform_L[802][9];				l_cell_reg[582] = inform_L[547][9];				l_cell_reg[583] = inform_L[803][9];				l_cell_reg[584] = inform_L[548][9];				l_cell_reg[585] = inform_L[804][9];				l_cell_reg[586] = inform_L[549][9];				l_cell_reg[587] = inform_L[805][9];				l_cell_reg[588] = inform_L[550][9];				l_cell_reg[589] = inform_L[806][9];				l_cell_reg[590] = inform_L[551][9];				l_cell_reg[591] = inform_L[807][9];				l_cell_reg[592] = inform_L[552][9];				l_cell_reg[593] = inform_L[808][9];				l_cell_reg[594] = inform_L[553][9];				l_cell_reg[595] = inform_L[809][9];				l_cell_reg[596] = inform_L[554][9];				l_cell_reg[597] = inform_L[810][9];				l_cell_reg[598] = inform_L[555][9];				l_cell_reg[599] = inform_L[811][9];				l_cell_reg[600] = inform_L[556][9];				l_cell_reg[601] = inform_L[812][9];				l_cell_reg[602] = inform_L[557][9];				l_cell_reg[603] = inform_L[813][9];				l_cell_reg[604] = inform_L[558][9];				l_cell_reg[605] = inform_L[814][9];				l_cell_reg[606] = inform_L[559][9];				l_cell_reg[607] = inform_L[815][9];				l_cell_reg[608] = inform_L[560][9];				l_cell_reg[609] = inform_L[816][9];				l_cell_reg[610] = inform_L[561][9];				l_cell_reg[611] = inform_L[817][9];				l_cell_reg[612] = inform_L[562][9];				l_cell_reg[613] = inform_L[818][9];				l_cell_reg[614] = inform_L[563][9];				l_cell_reg[615] = inform_L[819][9];				l_cell_reg[616] = inform_L[564][9];				l_cell_reg[617] = inform_L[820][9];				l_cell_reg[618] = inform_L[565][9];				l_cell_reg[619] = inform_L[821][9];				l_cell_reg[620] = inform_L[566][9];				l_cell_reg[621] = inform_L[822][9];				l_cell_reg[622] = inform_L[567][9];				l_cell_reg[623] = inform_L[823][9];				l_cell_reg[624] = inform_L[568][9];				l_cell_reg[625] = inform_L[824][9];				l_cell_reg[626] = inform_L[569][9];				l_cell_reg[627] = inform_L[825][9];				l_cell_reg[628] = inform_L[570][9];				l_cell_reg[629] = inform_L[826][9];				l_cell_reg[630] = inform_L[571][9];				l_cell_reg[631] = inform_L[827][9];				l_cell_reg[632] = inform_L[572][9];				l_cell_reg[633] = inform_L[828][9];				l_cell_reg[634] = inform_L[573][9];				l_cell_reg[635] = inform_L[829][9];				l_cell_reg[636] = inform_L[574][9];				l_cell_reg[637] = inform_L[830][9];				l_cell_reg[638] = inform_L[575][9];				l_cell_reg[639] = inform_L[831][9];				l_cell_reg[640] = inform_L[576][9];				l_cell_reg[641] = inform_L[832][9];				l_cell_reg[642] = inform_L[577][9];				l_cell_reg[643] = inform_L[833][9];				l_cell_reg[644] = inform_L[578][9];				l_cell_reg[645] = inform_L[834][9];				l_cell_reg[646] = inform_L[579][9];				l_cell_reg[647] = inform_L[835][9];				l_cell_reg[648] = inform_L[580][9];				l_cell_reg[649] = inform_L[836][9];				l_cell_reg[650] = inform_L[581][9];				l_cell_reg[651] = inform_L[837][9];				l_cell_reg[652] = inform_L[582][9];				l_cell_reg[653] = inform_L[838][9];				l_cell_reg[654] = inform_L[583][9];				l_cell_reg[655] = inform_L[839][9];				l_cell_reg[656] = inform_L[584][9];				l_cell_reg[657] = inform_L[840][9];				l_cell_reg[658] = inform_L[585][9];				l_cell_reg[659] = inform_L[841][9];				l_cell_reg[660] = inform_L[586][9];				l_cell_reg[661] = inform_L[842][9];				l_cell_reg[662] = inform_L[587][9];				l_cell_reg[663] = inform_L[843][9];				l_cell_reg[664] = inform_L[588][9];				l_cell_reg[665] = inform_L[844][9];				l_cell_reg[666] = inform_L[589][9];				l_cell_reg[667] = inform_L[845][9];				l_cell_reg[668] = inform_L[590][9];				l_cell_reg[669] = inform_L[846][9];				l_cell_reg[670] = inform_L[591][9];				l_cell_reg[671] = inform_L[847][9];				l_cell_reg[672] = inform_L[592][9];				l_cell_reg[673] = inform_L[848][9];				l_cell_reg[674] = inform_L[593][9];				l_cell_reg[675] = inform_L[849][9];				l_cell_reg[676] = inform_L[594][9];				l_cell_reg[677] = inform_L[850][9];				l_cell_reg[678] = inform_L[595][9];				l_cell_reg[679] = inform_L[851][9];				l_cell_reg[680] = inform_L[596][9];				l_cell_reg[681] = inform_L[852][9];				l_cell_reg[682] = inform_L[597][9];				l_cell_reg[683] = inform_L[853][9];				l_cell_reg[684] = inform_L[598][9];				l_cell_reg[685] = inform_L[854][9];				l_cell_reg[686] = inform_L[599][9];				l_cell_reg[687] = inform_L[855][9];				l_cell_reg[688] = inform_L[600][9];				l_cell_reg[689] = inform_L[856][9];				l_cell_reg[690] = inform_L[601][9];				l_cell_reg[691] = inform_L[857][9];				l_cell_reg[692] = inform_L[602][9];				l_cell_reg[693] = inform_L[858][9];				l_cell_reg[694] = inform_L[603][9];				l_cell_reg[695] = inform_L[859][9];				l_cell_reg[696] = inform_L[604][9];				l_cell_reg[697] = inform_L[860][9];				l_cell_reg[698] = inform_L[605][9];				l_cell_reg[699] = inform_L[861][9];				l_cell_reg[700] = inform_L[606][9];				l_cell_reg[701] = inform_L[862][9];				l_cell_reg[702] = inform_L[607][9];				l_cell_reg[703] = inform_L[863][9];				l_cell_reg[704] = inform_L[608][9];				l_cell_reg[705] = inform_L[864][9];				l_cell_reg[706] = inform_L[609][9];				l_cell_reg[707] = inform_L[865][9];				l_cell_reg[708] = inform_L[610][9];				l_cell_reg[709] = inform_L[866][9];				l_cell_reg[710] = inform_L[611][9];				l_cell_reg[711] = inform_L[867][9];				l_cell_reg[712] = inform_L[612][9];				l_cell_reg[713] = inform_L[868][9];				l_cell_reg[714] = inform_L[613][9];				l_cell_reg[715] = inform_L[869][9];				l_cell_reg[716] = inform_L[614][9];				l_cell_reg[717] = inform_L[870][9];				l_cell_reg[718] = inform_L[615][9];				l_cell_reg[719] = inform_L[871][9];				l_cell_reg[720] = inform_L[616][9];				l_cell_reg[721] = inform_L[872][9];				l_cell_reg[722] = inform_L[617][9];				l_cell_reg[723] = inform_L[873][9];				l_cell_reg[724] = inform_L[618][9];				l_cell_reg[725] = inform_L[874][9];				l_cell_reg[726] = inform_L[619][9];				l_cell_reg[727] = inform_L[875][9];				l_cell_reg[728] = inform_L[620][9];				l_cell_reg[729] = inform_L[876][9];				l_cell_reg[730] = inform_L[621][9];				l_cell_reg[731] = inform_L[877][9];				l_cell_reg[732] = inform_L[622][9];				l_cell_reg[733] = inform_L[878][9];				l_cell_reg[734] = inform_L[623][9];				l_cell_reg[735] = inform_L[879][9];				l_cell_reg[736] = inform_L[624][9];				l_cell_reg[737] = inform_L[880][9];				l_cell_reg[738] = inform_L[625][9];				l_cell_reg[739] = inform_L[881][9];				l_cell_reg[740] = inform_L[626][9];				l_cell_reg[741] = inform_L[882][9];				l_cell_reg[742] = inform_L[627][9];				l_cell_reg[743] = inform_L[883][9];				l_cell_reg[744] = inform_L[628][9];				l_cell_reg[745] = inform_L[884][9];				l_cell_reg[746] = inform_L[629][9];				l_cell_reg[747] = inform_L[885][9];				l_cell_reg[748] = inform_L[630][9];				l_cell_reg[749] = inform_L[886][9];				l_cell_reg[750] = inform_L[631][9];				l_cell_reg[751] = inform_L[887][9];				l_cell_reg[752] = inform_L[632][9];				l_cell_reg[753] = inform_L[888][9];				l_cell_reg[754] = inform_L[633][9];				l_cell_reg[755] = inform_L[889][9];				l_cell_reg[756] = inform_L[634][9];				l_cell_reg[757] = inform_L[890][9];				l_cell_reg[758] = inform_L[635][9];				l_cell_reg[759] = inform_L[891][9];				l_cell_reg[760] = inform_L[636][9];				l_cell_reg[761] = inform_L[892][9];				l_cell_reg[762] = inform_L[637][9];				l_cell_reg[763] = inform_L[893][9];				l_cell_reg[764] = inform_L[638][9];				l_cell_reg[765] = inform_L[894][9];				l_cell_reg[766] = inform_L[639][9];				l_cell_reg[767] = inform_L[895][9];				l_cell_reg[768] = inform_L[640][9];				l_cell_reg[769] = inform_L[896][9];				l_cell_reg[770] = inform_L[641][9];				l_cell_reg[771] = inform_L[897][9];				l_cell_reg[772] = inform_L[642][9];				l_cell_reg[773] = inform_L[898][9];				l_cell_reg[774] = inform_L[643][9];				l_cell_reg[775] = inform_L[899][9];				l_cell_reg[776] = inform_L[644][9];				l_cell_reg[777] = inform_L[900][9];				l_cell_reg[778] = inform_L[645][9];				l_cell_reg[779] = inform_L[901][9];				l_cell_reg[780] = inform_L[646][9];				l_cell_reg[781] = inform_L[902][9];				l_cell_reg[782] = inform_L[647][9];				l_cell_reg[783] = inform_L[903][9];				l_cell_reg[784] = inform_L[648][9];				l_cell_reg[785] = inform_L[904][9];				l_cell_reg[786] = inform_L[649][9];				l_cell_reg[787] = inform_L[905][9];				l_cell_reg[788] = inform_L[650][9];				l_cell_reg[789] = inform_L[906][9];				l_cell_reg[790] = inform_L[651][9];				l_cell_reg[791] = inform_L[907][9];				l_cell_reg[792] = inform_L[652][9];				l_cell_reg[793] = inform_L[908][9];				l_cell_reg[794] = inform_L[653][9];				l_cell_reg[795] = inform_L[909][9];				l_cell_reg[796] = inform_L[654][9];				l_cell_reg[797] = inform_L[910][9];				l_cell_reg[798] = inform_L[655][9];				l_cell_reg[799] = inform_L[911][9];				l_cell_reg[800] = inform_L[656][9];				l_cell_reg[801] = inform_L[912][9];				l_cell_reg[802] = inform_L[657][9];				l_cell_reg[803] = inform_L[913][9];				l_cell_reg[804] = inform_L[658][9];				l_cell_reg[805] = inform_L[914][9];				l_cell_reg[806] = inform_L[659][9];				l_cell_reg[807] = inform_L[915][9];				l_cell_reg[808] = inform_L[660][9];				l_cell_reg[809] = inform_L[916][9];				l_cell_reg[810] = inform_L[661][9];				l_cell_reg[811] = inform_L[917][9];				l_cell_reg[812] = inform_L[662][9];				l_cell_reg[813] = inform_L[918][9];				l_cell_reg[814] = inform_L[663][9];				l_cell_reg[815] = inform_L[919][9];				l_cell_reg[816] = inform_L[664][9];				l_cell_reg[817] = inform_L[920][9];				l_cell_reg[818] = inform_L[665][9];				l_cell_reg[819] = inform_L[921][9];				l_cell_reg[820] = inform_L[666][9];				l_cell_reg[821] = inform_L[922][9];				l_cell_reg[822] = inform_L[667][9];				l_cell_reg[823] = inform_L[923][9];				l_cell_reg[824] = inform_L[668][9];				l_cell_reg[825] = inform_L[924][9];				l_cell_reg[826] = inform_L[669][9];				l_cell_reg[827] = inform_L[925][9];				l_cell_reg[828] = inform_L[670][9];				l_cell_reg[829] = inform_L[926][9];				l_cell_reg[830] = inform_L[671][9];				l_cell_reg[831] = inform_L[927][9];				l_cell_reg[832] = inform_L[672][9];				l_cell_reg[833] = inform_L[928][9];				l_cell_reg[834] = inform_L[673][9];				l_cell_reg[835] = inform_L[929][9];				l_cell_reg[836] = inform_L[674][9];				l_cell_reg[837] = inform_L[930][9];				l_cell_reg[838] = inform_L[675][9];				l_cell_reg[839] = inform_L[931][9];				l_cell_reg[840] = inform_L[676][9];				l_cell_reg[841] = inform_L[932][9];				l_cell_reg[842] = inform_L[677][9];				l_cell_reg[843] = inform_L[933][9];				l_cell_reg[844] = inform_L[678][9];				l_cell_reg[845] = inform_L[934][9];				l_cell_reg[846] = inform_L[679][9];				l_cell_reg[847] = inform_L[935][9];				l_cell_reg[848] = inform_L[680][9];				l_cell_reg[849] = inform_L[936][9];				l_cell_reg[850] = inform_L[681][9];				l_cell_reg[851] = inform_L[937][9];				l_cell_reg[852] = inform_L[682][9];				l_cell_reg[853] = inform_L[938][9];				l_cell_reg[854] = inform_L[683][9];				l_cell_reg[855] = inform_L[939][9];				l_cell_reg[856] = inform_L[684][9];				l_cell_reg[857] = inform_L[940][9];				l_cell_reg[858] = inform_L[685][9];				l_cell_reg[859] = inform_L[941][9];				l_cell_reg[860] = inform_L[686][9];				l_cell_reg[861] = inform_L[942][9];				l_cell_reg[862] = inform_L[687][9];				l_cell_reg[863] = inform_L[943][9];				l_cell_reg[864] = inform_L[688][9];				l_cell_reg[865] = inform_L[944][9];				l_cell_reg[866] = inform_L[689][9];				l_cell_reg[867] = inform_L[945][9];				l_cell_reg[868] = inform_L[690][9];				l_cell_reg[869] = inform_L[946][9];				l_cell_reg[870] = inform_L[691][9];				l_cell_reg[871] = inform_L[947][9];				l_cell_reg[872] = inform_L[692][9];				l_cell_reg[873] = inform_L[948][9];				l_cell_reg[874] = inform_L[693][9];				l_cell_reg[875] = inform_L[949][9];				l_cell_reg[876] = inform_L[694][9];				l_cell_reg[877] = inform_L[950][9];				l_cell_reg[878] = inform_L[695][9];				l_cell_reg[879] = inform_L[951][9];				l_cell_reg[880] = inform_L[696][9];				l_cell_reg[881] = inform_L[952][9];				l_cell_reg[882] = inform_L[697][9];				l_cell_reg[883] = inform_L[953][9];				l_cell_reg[884] = inform_L[698][9];				l_cell_reg[885] = inform_L[954][9];				l_cell_reg[886] = inform_L[699][9];				l_cell_reg[887] = inform_L[955][9];				l_cell_reg[888] = inform_L[700][9];				l_cell_reg[889] = inform_L[956][9];				l_cell_reg[890] = inform_L[701][9];				l_cell_reg[891] = inform_L[957][9];				l_cell_reg[892] = inform_L[702][9];				l_cell_reg[893] = inform_L[958][9];				l_cell_reg[894] = inform_L[703][9];				l_cell_reg[895] = inform_L[959][9];				l_cell_reg[896] = inform_L[704][9];				l_cell_reg[897] = inform_L[960][9];				l_cell_reg[898] = inform_L[705][9];				l_cell_reg[899] = inform_L[961][9];				l_cell_reg[900] = inform_L[706][9];				l_cell_reg[901] = inform_L[962][9];				l_cell_reg[902] = inform_L[707][9];				l_cell_reg[903] = inform_L[963][9];				l_cell_reg[904] = inform_L[708][9];				l_cell_reg[905] = inform_L[964][9];				l_cell_reg[906] = inform_L[709][9];				l_cell_reg[907] = inform_L[965][9];				l_cell_reg[908] = inform_L[710][9];				l_cell_reg[909] = inform_L[966][9];				l_cell_reg[910] = inform_L[711][9];				l_cell_reg[911] = inform_L[967][9];				l_cell_reg[912] = inform_L[712][9];				l_cell_reg[913] = inform_L[968][9];				l_cell_reg[914] = inform_L[713][9];				l_cell_reg[915] = inform_L[969][9];				l_cell_reg[916] = inform_L[714][9];				l_cell_reg[917] = inform_L[970][9];				l_cell_reg[918] = inform_L[715][9];				l_cell_reg[919] = inform_L[971][9];				l_cell_reg[920] = inform_L[716][9];				l_cell_reg[921] = inform_L[972][9];				l_cell_reg[922] = inform_L[717][9];				l_cell_reg[923] = inform_L[973][9];				l_cell_reg[924] = inform_L[718][9];				l_cell_reg[925] = inform_L[974][9];				l_cell_reg[926] = inform_L[719][9];				l_cell_reg[927] = inform_L[975][9];				l_cell_reg[928] = inform_L[720][9];				l_cell_reg[929] = inform_L[976][9];				l_cell_reg[930] = inform_L[721][9];				l_cell_reg[931] = inform_L[977][9];				l_cell_reg[932] = inform_L[722][9];				l_cell_reg[933] = inform_L[978][9];				l_cell_reg[934] = inform_L[723][9];				l_cell_reg[935] = inform_L[979][9];				l_cell_reg[936] = inform_L[724][9];				l_cell_reg[937] = inform_L[980][9];				l_cell_reg[938] = inform_L[725][9];				l_cell_reg[939] = inform_L[981][9];				l_cell_reg[940] = inform_L[726][9];				l_cell_reg[941] = inform_L[982][9];				l_cell_reg[942] = inform_L[727][9];				l_cell_reg[943] = inform_L[983][9];				l_cell_reg[944] = inform_L[728][9];				l_cell_reg[945] = inform_L[984][9];				l_cell_reg[946] = inform_L[729][9];				l_cell_reg[947] = inform_L[985][9];				l_cell_reg[948] = inform_L[730][9];				l_cell_reg[949] = inform_L[986][9];				l_cell_reg[950] = inform_L[731][9];				l_cell_reg[951] = inform_L[987][9];				l_cell_reg[952] = inform_L[732][9];				l_cell_reg[953] = inform_L[988][9];				l_cell_reg[954] = inform_L[733][9];				l_cell_reg[955] = inform_L[989][9];				l_cell_reg[956] = inform_L[734][9];				l_cell_reg[957] = inform_L[990][9];				l_cell_reg[958] = inform_L[735][9];				l_cell_reg[959] = inform_L[991][9];				l_cell_reg[960] = inform_L[736][9];				l_cell_reg[961] = inform_L[992][9];				l_cell_reg[962] = inform_L[737][9];				l_cell_reg[963] = inform_L[993][9];				l_cell_reg[964] = inform_L[738][9];				l_cell_reg[965] = inform_L[994][9];				l_cell_reg[966] = inform_L[739][9];				l_cell_reg[967] = inform_L[995][9];				l_cell_reg[968] = inform_L[740][9];				l_cell_reg[969] = inform_L[996][9];				l_cell_reg[970] = inform_L[741][9];				l_cell_reg[971] = inform_L[997][9];				l_cell_reg[972] = inform_L[742][9];				l_cell_reg[973] = inform_L[998][9];				l_cell_reg[974] = inform_L[743][9];				l_cell_reg[975] = inform_L[999][9];				l_cell_reg[976] = inform_L[744][9];				l_cell_reg[977] = inform_L[1000][9];				l_cell_reg[978] = inform_L[745][9];				l_cell_reg[979] = inform_L[1001][9];				l_cell_reg[980] = inform_L[746][9];				l_cell_reg[981] = inform_L[1002][9];				l_cell_reg[982] = inform_L[747][9];				l_cell_reg[983] = inform_L[1003][9];				l_cell_reg[984] = inform_L[748][9];				l_cell_reg[985] = inform_L[1004][9];				l_cell_reg[986] = inform_L[749][9];				l_cell_reg[987] = inform_L[1005][9];				l_cell_reg[988] = inform_L[750][9];				l_cell_reg[989] = inform_L[1006][9];				l_cell_reg[990] = inform_L[751][9];				l_cell_reg[991] = inform_L[1007][9];				l_cell_reg[992] = inform_L[752][9];				l_cell_reg[993] = inform_L[1008][9];				l_cell_reg[994] = inform_L[753][9];				l_cell_reg[995] = inform_L[1009][9];				l_cell_reg[996] = inform_L[754][9];				l_cell_reg[997] = inform_L[1010][9];				l_cell_reg[998] = inform_L[755][9];				l_cell_reg[999] = inform_L[1011][9];				l_cell_reg[1000] = inform_L[756][9];				l_cell_reg[1001] = inform_L[1012][9];				l_cell_reg[1002] = inform_L[757][9];				l_cell_reg[1003] = inform_L[1013][9];				l_cell_reg[1004] = inform_L[758][9];				l_cell_reg[1005] = inform_L[1014][9];				l_cell_reg[1006] = inform_L[759][9];				l_cell_reg[1007] = inform_L[1015][9];				l_cell_reg[1008] = inform_L[760][9];				l_cell_reg[1009] = inform_L[1016][9];				l_cell_reg[1010] = inform_L[761][9];				l_cell_reg[1011] = inform_L[1017][9];				l_cell_reg[1012] = inform_L[762][9];				l_cell_reg[1013] = inform_L[1018][9];				l_cell_reg[1014] = inform_L[763][9];				l_cell_reg[1015] = inform_L[1019][9];				l_cell_reg[1016] = inform_L[764][9];				l_cell_reg[1017] = inform_L[1020][9];				l_cell_reg[1018] = inform_L[765][9];				l_cell_reg[1019] = inform_L[1021][9];				l_cell_reg[1020] = inform_L[766][9];				l_cell_reg[1021] = inform_L[1022][9];				l_cell_reg[1022] = inform_L[767][9];				l_cell_reg[1023] = inform_L[1023][9];			end
			10:			begin				r_cell_reg[0] = inform_R[0][9];				r_cell_reg[1] = inform_R[512][9];				r_cell_reg[2] = inform_R[1][9];				r_cell_reg[3] = inform_R[513][9];				r_cell_reg[4] = inform_R[2][9];				r_cell_reg[5] = inform_R[514][9];				r_cell_reg[6] = inform_R[3][9];				r_cell_reg[7] = inform_R[515][9];				r_cell_reg[8] = inform_R[4][9];				r_cell_reg[9] = inform_R[516][9];				r_cell_reg[10] = inform_R[5][9];				r_cell_reg[11] = inform_R[517][9];				r_cell_reg[12] = inform_R[6][9];				r_cell_reg[13] = inform_R[518][9];				r_cell_reg[14] = inform_R[7][9];				r_cell_reg[15] = inform_R[519][9];				r_cell_reg[16] = inform_R[8][9];				r_cell_reg[17] = inform_R[520][9];				r_cell_reg[18] = inform_R[9][9];				r_cell_reg[19] = inform_R[521][9];				r_cell_reg[20] = inform_R[10][9];				r_cell_reg[21] = inform_R[522][9];				r_cell_reg[22] = inform_R[11][9];				r_cell_reg[23] = inform_R[523][9];				r_cell_reg[24] = inform_R[12][9];				r_cell_reg[25] = inform_R[524][9];				r_cell_reg[26] = inform_R[13][9];				r_cell_reg[27] = inform_R[525][9];				r_cell_reg[28] = inform_R[14][9];				r_cell_reg[29] = inform_R[526][9];				r_cell_reg[30] = inform_R[15][9];				r_cell_reg[31] = inform_R[527][9];				r_cell_reg[32] = inform_R[16][9];				r_cell_reg[33] = inform_R[528][9];				r_cell_reg[34] = inform_R[17][9];				r_cell_reg[35] = inform_R[529][9];				r_cell_reg[36] = inform_R[18][9];				r_cell_reg[37] = inform_R[530][9];				r_cell_reg[38] = inform_R[19][9];				r_cell_reg[39] = inform_R[531][9];				r_cell_reg[40] = inform_R[20][9];				r_cell_reg[41] = inform_R[532][9];				r_cell_reg[42] = inform_R[21][9];				r_cell_reg[43] = inform_R[533][9];				r_cell_reg[44] = inform_R[22][9];				r_cell_reg[45] = inform_R[534][9];				r_cell_reg[46] = inform_R[23][9];				r_cell_reg[47] = inform_R[535][9];				r_cell_reg[48] = inform_R[24][9];				r_cell_reg[49] = inform_R[536][9];				r_cell_reg[50] = inform_R[25][9];				r_cell_reg[51] = inform_R[537][9];				r_cell_reg[52] = inform_R[26][9];				r_cell_reg[53] = inform_R[538][9];				r_cell_reg[54] = inform_R[27][9];				r_cell_reg[55] = inform_R[539][9];				r_cell_reg[56] = inform_R[28][9];				r_cell_reg[57] = inform_R[540][9];				r_cell_reg[58] = inform_R[29][9];				r_cell_reg[59] = inform_R[541][9];				r_cell_reg[60] = inform_R[30][9];				r_cell_reg[61] = inform_R[542][9];				r_cell_reg[62] = inform_R[31][9];				r_cell_reg[63] = inform_R[543][9];				r_cell_reg[64] = inform_R[32][9];				r_cell_reg[65] = inform_R[544][9];				r_cell_reg[66] = inform_R[33][9];				r_cell_reg[67] = inform_R[545][9];				r_cell_reg[68] = inform_R[34][9];				r_cell_reg[69] = inform_R[546][9];				r_cell_reg[70] = inform_R[35][9];				r_cell_reg[71] = inform_R[547][9];				r_cell_reg[72] = inform_R[36][9];				r_cell_reg[73] = inform_R[548][9];				r_cell_reg[74] = inform_R[37][9];				r_cell_reg[75] = inform_R[549][9];				r_cell_reg[76] = inform_R[38][9];				r_cell_reg[77] = inform_R[550][9];				r_cell_reg[78] = inform_R[39][9];				r_cell_reg[79] = inform_R[551][9];				r_cell_reg[80] = inform_R[40][9];				r_cell_reg[81] = inform_R[552][9];				r_cell_reg[82] = inform_R[41][9];				r_cell_reg[83] = inform_R[553][9];				r_cell_reg[84] = inform_R[42][9];				r_cell_reg[85] = inform_R[554][9];				r_cell_reg[86] = inform_R[43][9];				r_cell_reg[87] = inform_R[555][9];				r_cell_reg[88] = inform_R[44][9];				r_cell_reg[89] = inform_R[556][9];				r_cell_reg[90] = inform_R[45][9];				r_cell_reg[91] = inform_R[557][9];				r_cell_reg[92] = inform_R[46][9];				r_cell_reg[93] = inform_R[558][9];				r_cell_reg[94] = inform_R[47][9];				r_cell_reg[95] = inform_R[559][9];				r_cell_reg[96] = inform_R[48][9];				r_cell_reg[97] = inform_R[560][9];				r_cell_reg[98] = inform_R[49][9];				r_cell_reg[99] = inform_R[561][9];				r_cell_reg[100] = inform_R[50][9];				r_cell_reg[101] = inform_R[562][9];				r_cell_reg[102] = inform_R[51][9];				r_cell_reg[103] = inform_R[563][9];				r_cell_reg[104] = inform_R[52][9];				r_cell_reg[105] = inform_R[564][9];				r_cell_reg[106] = inform_R[53][9];				r_cell_reg[107] = inform_R[565][9];				r_cell_reg[108] = inform_R[54][9];				r_cell_reg[109] = inform_R[566][9];				r_cell_reg[110] = inform_R[55][9];				r_cell_reg[111] = inform_R[567][9];				r_cell_reg[112] = inform_R[56][9];				r_cell_reg[113] = inform_R[568][9];				r_cell_reg[114] = inform_R[57][9];				r_cell_reg[115] = inform_R[569][9];				r_cell_reg[116] = inform_R[58][9];				r_cell_reg[117] = inform_R[570][9];				r_cell_reg[118] = inform_R[59][9];				r_cell_reg[119] = inform_R[571][9];				r_cell_reg[120] = inform_R[60][9];				r_cell_reg[121] = inform_R[572][9];				r_cell_reg[122] = inform_R[61][9];				r_cell_reg[123] = inform_R[573][9];				r_cell_reg[124] = inform_R[62][9];				r_cell_reg[125] = inform_R[574][9];				r_cell_reg[126] = inform_R[63][9];				r_cell_reg[127] = inform_R[575][9];				r_cell_reg[128] = inform_R[64][9];				r_cell_reg[129] = inform_R[576][9];				r_cell_reg[130] = inform_R[65][9];				r_cell_reg[131] = inform_R[577][9];				r_cell_reg[132] = inform_R[66][9];				r_cell_reg[133] = inform_R[578][9];				r_cell_reg[134] = inform_R[67][9];				r_cell_reg[135] = inform_R[579][9];				r_cell_reg[136] = inform_R[68][9];				r_cell_reg[137] = inform_R[580][9];				r_cell_reg[138] = inform_R[69][9];				r_cell_reg[139] = inform_R[581][9];				r_cell_reg[140] = inform_R[70][9];				r_cell_reg[141] = inform_R[582][9];				r_cell_reg[142] = inform_R[71][9];				r_cell_reg[143] = inform_R[583][9];				r_cell_reg[144] = inform_R[72][9];				r_cell_reg[145] = inform_R[584][9];				r_cell_reg[146] = inform_R[73][9];				r_cell_reg[147] = inform_R[585][9];				r_cell_reg[148] = inform_R[74][9];				r_cell_reg[149] = inform_R[586][9];				r_cell_reg[150] = inform_R[75][9];				r_cell_reg[151] = inform_R[587][9];				r_cell_reg[152] = inform_R[76][9];				r_cell_reg[153] = inform_R[588][9];				r_cell_reg[154] = inform_R[77][9];				r_cell_reg[155] = inform_R[589][9];				r_cell_reg[156] = inform_R[78][9];				r_cell_reg[157] = inform_R[590][9];				r_cell_reg[158] = inform_R[79][9];				r_cell_reg[159] = inform_R[591][9];				r_cell_reg[160] = inform_R[80][9];				r_cell_reg[161] = inform_R[592][9];				r_cell_reg[162] = inform_R[81][9];				r_cell_reg[163] = inform_R[593][9];				r_cell_reg[164] = inform_R[82][9];				r_cell_reg[165] = inform_R[594][9];				r_cell_reg[166] = inform_R[83][9];				r_cell_reg[167] = inform_R[595][9];				r_cell_reg[168] = inform_R[84][9];				r_cell_reg[169] = inform_R[596][9];				r_cell_reg[170] = inform_R[85][9];				r_cell_reg[171] = inform_R[597][9];				r_cell_reg[172] = inform_R[86][9];				r_cell_reg[173] = inform_R[598][9];				r_cell_reg[174] = inform_R[87][9];				r_cell_reg[175] = inform_R[599][9];				r_cell_reg[176] = inform_R[88][9];				r_cell_reg[177] = inform_R[600][9];				r_cell_reg[178] = inform_R[89][9];				r_cell_reg[179] = inform_R[601][9];				r_cell_reg[180] = inform_R[90][9];				r_cell_reg[181] = inform_R[602][9];				r_cell_reg[182] = inform_R[91][9];				r_cell_reg[183] = inform_R[603][9];				r_cell_reg[184] = inform_R[92][9];				r_cell_reg[185] = inform_R[604][9];				r_cell_reg[186] = inform_R[93][9];				r_cell_reg[187] = inform_R[605][9];				r_cell_reg[188] = inform_R[94][9];				r_cell_reg[189] = inform_R[606][9];				r_cell_reg[190] = inform_R[95][9];				r_cell_reg[191] = inform_R[607][9];				r_cell_reg[192] = inform_R[96][9];				r_cell_reg[193] = inform_R[608][9];				r_cell_reg[194] = inform_R[97][9];				r_cell_reg[195] = inform_R[609][9];				r_cell_reg[196] = inform_R[98][9];				r_cell_reg[197] = inform_R[610][9];				r_cell_reg[198] = inform_R[99][9];				r_cell_reg[199] = inform_R[611][9];				r_cell_reg[200] = inform_R[100][9];				r_cell_reg[201] = inform_R[612][9];				r_cell_reg[202] = inform_R[101][9];				r_cell_reg[203] = inform_R[613][9];				r_cell_reg[204] = inform_R[102][9];				r_cell_reg[205] = inform_R[614][9];				r_cell_reg[206] = inform_R[103][9];				r_cell_reg[207] = inform_R[615][9];				r_cell_reg[208] = inform_R[104][9];				r_cell_reg[209] = inform_R[616][9];				r_cell_reg[210] = inform_R[105][9];				r_cell_reg[211] = inform_R[617][9];				r_cell_reg[212] = inform_R[106][9];				r_cell_reg[213] = inform_R[618][9];				r_cell_reg[214] = inform_R[107][9];				r_cell_reg[215] = inform_R[619][9];				r_cell_reg[216] = inform_R[108][9];				r_cell_reg[217] = inform_R[620][9];				r_cell_reg[218] = inform_R[109][9];				r_cell_reg[219] = inform_R[621][9];				r_cell_reg[220] = inform_R[110][9];				r_cell_reg[221] = inform_R[622][9];				r_cell_reg[222] = inform_R[111][9];				r_cell_reg[223] = inform_R[623][9];				r_cell_reg[224] = inform_R[112][9];				r_cell_reg[225] = inform_R[624][9];				r_cell_reg[226] = inform_R[113][9];				r_cell_reg[227] = inform_R[625][9];				r_cell_reg[228] = inform_R[114][9];				r_cell_reg[229] = inform_R[626][9];				r_cell_reg[230] = inform_R[115][9];				r_cell_reg[231] = inform_R[627][9];				r_cell_reg[232] = inform_R[116][9];				r_cell_reg[233] = inform_R[628][9];				r_cell_reg[234] = inform_R[117][9];				r_cell_reg[235] = inform_R[629][9];				r_cell_reg[236] = inform_R[118][9];				r_cell_reg[237] = inform_R[630][9];				r_cell_reg[238] = inform_R[119][9];				r_cell_reg[239] = inform_R[631][9];				r_cell_reg[240] = inform_R[120][9];				r_cell_reg[241] = inform_R[632][9];				r_cell_reg[242] = inform_R[121][9];				r_cell_reg[243] = inform_R[633][9];				r_cell_reg[244] = inform_R[122][9];				r_cell_reg[245] = inform_R[634][9];				r_cell_reg[246] = inform_R[123][9];				r_cell_reg[247] = inform_R[635][9];				r_cell_reg[248] = inform_R[124][9];				r_cell_reg[249] = inform_R[636][9];				r_cell_reg[250] = inform_R[125][9];				r_cell_reg[251] = inform_R[637][9];				r_cell_reg[252] = inform_R[126][9];				r_cell_reg[253] = inform_R[638][9];				r_cell_reg[254] = inform_R[127][9];				r_cell_reg[255] = inform_R[639][9];				r_cell_reg[256] = inform_R[128][9];				r_cell_reg[257] = inform_R[640][9];				r_cell_reg[258] = inform_R[129][9];				r_cell_reg[259] = inform_R[641][9];				r_cell_reg[260] = inform_R[130][9];				r_cell_reg[261] = inform_R[642][9];				r_cell_reg[262] = inform_R[131][9];				r_cell_reg[263] = inform_R[643][9];				r_cell_reg[264] = inform_R[132][9];				r_cell_reg[265] = inform_R[644][9];				r_cell_reg[266] = inform_R[133][9];				r_cell_reg[267] = inform_R[645][9];				r_cell_reg[268] = inform_R[134][9];				r_cell_reg[269] = inform_R[646][9];				r_cell_reg[270] = inform_R[135][9];				r_cell_reg[271] = inform_R[647][9];				r_cell_reg[272] = inform_R[136][9];				r_cell_reg[273] = inform_R[648][9];				r_cell_reg[274] = inform_R[137][9];				r_cell_reg[275] = inform_R[649][9];				r_cell_reg[276] = inform_R[138][9];				r_cell_reg[277] = inform_R[650][9];				r_cell_reg[278] = inform_R[139][9];				r_cell_reg[279] = inform_R[651][9];				r_cell_reg[280] = inform_R[140][9];				r_cell_reg[281] = inform_R[652][9];				r_cell_reg[282] = inform_R[141][9];				r_cell_reg[283] = inform_R[653][9];				r_cell_reg[284] = inform_R[142][9];				r_cell_reg[285] = inform_R[654][9];				r_cell_reg[286] = inform_R[143][9];				r_cell_reg[287] = inform_R[655][9];				r_cell_reg[288] = inform_R[144][9];				r_cell_reg[289] = inform_R[656][9];				r_cell_reg[290] = inform_R[145][9];				r_cell_reg[291] = inform_R[657][9];				r_cell_reg[292] = inform_R[146][9];				r_cell_reg[293] = inform_R[658][9];				r_cell_reg[294] = inform_R[147][9];				r_cell_reg[295] = inform_R[659][9];				r_cell_reg[296] = inform_R[148][9];				r_cell_reg[297] = inform_R[660][9];				r_cell_reg[298] = inform_R[149][9];				r_cell_reg[299] = inform_R[661][9];				r_cell_reg[300] = inform_R[150][9];				r_cell_reg[301] = inform_R[662][9];				r_cell_reg[302] = inform_R[151][9];				r_cell_reg[303] = inform_R[663][9];				r_cell_reg[304] = inform_R[152][9];				r_cell_reg[305] = inform_R[664][9];				r_cell_reg[306] = inform_R[153][9];				r_cell_reg[307] = inform_R[665][9];				r_cell_reg[308] = inform_R[154][9];				r_cell_reg[309] = inform_R[666][9];				r_cell_reg[310] = inform_R[155][9];				r_cell_reg[311] = inform_R[667][9];				r_cell_reg[312] = inform_R[156][9];				r_cell_reg[313] = inform_R[668][9];				r_cell_reg[314] = inform_R[157][9];				r_cell_reg[315] = inform_R[669][9];				r_cell_reg[316] = inform_R[158][9];				r_cell_reg[317] = inform_R[670][9];				r_cell_reg[318] = inform_R[159][9];				r_cell_reg[319] = inform_R[671][9];				r_cell_reg[320] = inform_R[160][9];				r_cell_reg[321] = inform_R[672][9];				r_cell_reg[322] = inform_R[161][9];				r_cell_reg[323] = inform_R[673][9];				r_cell_reg[324] = inform_R[162][9];				r_cell_reg[325] = inform_R[674][9];				r_cell_reg[326] = inform_R[163][9];				r_cell_reg[327] = inform_R[675][9];				r_cell_reg[328] = inform_R[164][9];				r_cell_reg[329] = inform_R[676][9];				r_cell_reg[330] = inform_R[165][9];				r_cell_reg[331] = inform_R[677][9];				r_cell_reg[332] = inform_R[166][9];				r_cell_reg[333] = inform_R[678][9];				r_cell_reg[334] = inform_R[167][9];				r_cell_reg[335] = inform_R[679][9];				r_cell_reg[336] = inform_R[168][9];				r_cell_reg[337] = inform_R[680][9];				r_cell_reg[338] = inform_R[169][9];				r_cell_reg[339] = inform_R[681][9];				r_cell_reg[340] = inform_R[170][9];				r_cell_reg[341] = inform_R[682][9];				r_cell_reg[342] = inform_R[171][9];				r_cell_reg[343] = inform_R[683][9];				r_cell_reg[344] = inform_R[172][9];				r_cell_reg[345] = inform_R[684][9];				r_cell_reg[346] = inform_R[173][9];				r_cell_reg[347] = inform_R[685][9];				r_cell_reg[348] = inform_R[174][9];				r_cell_reg[349] = inform_R[686][9];				r_cell_reg[350] = inform_R[175][9];				r_cell_reg[351] = inform_R[687][9];				r_cell_reg[352] = inform_R[176][9];				r_cell_reg[353] = inform_R[688][9];				r_cell_reg[354] = inform_R[177][9];				r_cell_reg[355] = inform_R[689][9];				r_cell_reg[356] = inform_R[178][9];				r_cell_reg[357] = inform_R[690][9];				r_cell_reg[358] = inform_R[179][9];				r_cell_reg[359] = inform_R[691][9];				r_cell_reg[360] = inform_R[180][9];				r_cell_reg[361] = inform_R[692][9];				r_cell_reg[362] = inform_R[181][9];				r_cell_reg[363] = inform_R[693][9];				r_cell_reg[364] = inform_R[182][9];				r_cell_reg[365] = inform_R[694][9];				r_cell_reg[366] = inform_R[183][9];				r_cell_reg[367] = inform_R[695][9];				r_cell_reg[368] = inform_R[184][9];				r_cell_reg[369] = inform_R[696][9];				r_cell_reg[370] = inform_R[185][9];				r_cell_reg[371] = inform_R[697][9];				r_cell_reg[372] = inform_R[186][9];				r_cell_reg[373] = inform_R[698][9];				r_cell_reg[374] = inform_R[187][9];				r_cell_reg[375] = inform_R[699][9];				r_cell_reg[376] = inform_R[188][9];				r_cell_reg[377] = inform_R[700][9];				r_cell_reg[378] = inform_R[189][9];				r_cell_reg[379] = inform_R[701][9];				r_cell_reg[380] = inform_R[190][9];				r_cell_reg[381] = inform_R[702][9];				r_cell_reg[382] = inform_R[191][9];				r_cell_reg[383] = inform_R[703][9];				r_cell_reg[384] = inform_R[192][9];				r_cell_reg[385] = inform_R[704][9];				r_cell_reg[386] = inform_R[193][9];				r_cell_reg[387] = inform_R[705][9];				r_cell_reg[388] = inform_R[194][9];				r_cell_reg[389] = inform_R[706][9];				r_cell_reg[390] = inform_R[195][9];				r_cell_reg[391] = inform_R[707][9];				r_cell_reg[392] = inform_R[196][9];				r_cell_reg[393] = inform_R[708][9];				r_cell_reg[394] = inform_R[197][9];				r_cell_reg[395] = inform_R[709][9];				r_cell_reg[396] = inform_R[198][9];				r_cell_reg[397] = inform_R[710][9];				r_cell_reg[398] = inform_R[199][9];				r_cell_reg[399] = inform_R[711][9];				r_cell_reg[400] = inform_R[200][9];				r_cell_reg[401] = inform_R[712][9];				r_cell_reg[402] = inform_R[201][9];				r_cell_reg[403] = inform_R[713][9];				r_cell_reg[404] = inform_R[202][9];				r_cell_reg[405] = inform_R[714][9];				r_cell_reg[406] = inform_R[203][9];				r_cell_reg[407] = inform_R[715][9];				r_cell_reg[408] = inform_R[204][9];				r_cell_reg[409] = inform_R[716][9];				r_cell_reg[410] = inform_R[205][9];				r_cell_reg[411] = inform_R[717][9];				r_cell_reg[412] = inform_R[206][9];				r_cell_reg[413] = inform_R[718][9];				r_cell_reg[414] = inform_R[207][9];				r_cell_reg[415] = inform_R[719][9];				r_cell_reg[416] = inform_R[208][9];				r_cell_reg[417] = inform_R[720][9];				r_cell_reg[418] = inform_R[209][9];				r_cell_reg[419] = inform_R[721][9];				r_cell_reg[420] = inform_R[210][9];				r_cell_reg[421] = inform_R[722][9];				r_cell_reg[422] = inform_R[211][9];				r_cell_reg[423] = inform_R[723][9];				r_cell_reg[424] = inform_R[212][9];				r_cell_reg[425] = inform_R[724][9];				r_cell_reg[426] = inform_R[213][9];				r_cell_reg[427] = inform_R[725][9];				r_cell_reg[428] = inform_R[214][9];				r_cell_reg[429] = inform_R[726][9];				r_cell_reg[430] = inform_R[215][9];				r_cell_reg[431] = inform_R[727][9];				r_cell_reg[432] = inform_R[216][9];				r_cell_reg[433] = inform_R[728][9];				r_cell_reg[434] = inform_R[217][9];				r_cell_reg[435] = inform_R[729][9];				r_cell_reg[436] = inform_R[218][9];				r_cell_reg[437] = inform_R[730][9];				r_cell_reg[438] = inform_R[219][9];				r_cell_reg[439] = inform_R[731][9];				r_cell_reg[440] = inform_R[220][9];				r_cell_reg[441] = inform_R[732][9];				r_cell_reg[442] = inform_R[221][9];				r_cell_reg[443] = inform_R[733][9];				r_cell_reg[444] = inform_R[222][9];				r_cell_reg[445] = inform_R[734][9];				r_cell_reg[446] = inform_R[223][9];				r_cell_reg[447] = inform_R[735][9];				r_cell_reg[448] = inform_R[224][9];				r_cell_reg[449] = inform_R[736][9];				r_cell_reg[450] = inform_R[225][9];				r_cell_reg[451] = inform_R[737][9];				r_cell_reg[452] = inform_R[226][9];				r_cell_reg[453] = inform_R[738][9];				r_cell_reg[454] = inform_R[227][9];				r_cell_reg[455] = inform_R[739][9];				r_cell_reg[456] = inform_R[228][9];				r_cell_reg[457] = inform_R[740][9];				r_cell_reg[458] = inform_R[229][9];				r_cell_reg[459] = inform_R[741][9];				r_cell_reg[460] = inform_R[230][9];				r_cell_reg[461] = inform_R[742][9];				r_cell_reg[462] = inform_R[231][9];				r_cell_reg[463] = inform_R[743][9];				r_cell_reg[464] = inform_R[232][9];				r_cell_reg[465] = inform_R[744][9];				r_cell_reg[466] = inform_R[233][9];				r_cell_reg[467] = inform_R[745][9];				r_cell_reg[468] = inform_R[234][9];				r_cell_reg[469] = inform_R[746][9];				r_cell_reg[470] = inform_R[235][9];				r_cell_reg[471] = inform_R[747][9];				r_cell_reg[472] = inform_R[236][9];				r_cell_reg[473] = inform_R[748][9];				r_cell_reg[474] = inform_R[237][9];				r_cell_reg[475] = inform_R[749][9];				r_cell_reg[476] = inform_R[238][9];				r_cell_reg[477] = inform_R[750][9];				r_cell_reg[478] = inform_R[239][9];				r_cell_reg[479] = inform_R[751][9];				r_cell_reg[480] = inform_R[240][9];				r_cell_reg[481] = inform_R[752][9];				r_cell_reg[482] = inform_R[241][9];				r_cell_reg[483] = inform_R[753][9];				r_cell_reg[484] = inform_R[242][9];				r_cell_reg[485] = inform_R[754][9];				r_cell_reg[486] = inform_R[243][9];				r_cell_reg[487] = inform_R[755][9];				r_cell_reg[488] = inform_R[244][9];				r_cell_reg[489] = inform_R[756][9];				r_cell_reg[490] = inform_R[245][9];				r_cell_reg[491] = inform_R[757][9];				r_cell_reg[492] = inform_R[246][9];				r_cell_reg[493] = inform_R[758][9];				r_cell_reg[494] = inform_R[247][9];				r_cell_reg[495] = inform_R[759][9];				r_cell_reg[496] = inform_R[248][9];				r_cell_reg[497] = inform_R[760][9];				r_cell_reg[498] = inform_R[249][9];				r_cell_reg[499] = inform_R[761][9];				r_cell_reg[500] = inform_R[250][9];				r_cell_reg[501] = inform_R[762][9];				r_cell_reg[502] = inform_R[251][9];				r_cell_reg[503] = inform_R[763][9];				r_cell_reg[504] = inform_R[252][9];				r_cell_reg[505] = inform_R[764][9];				r_cell_reg[506] = inform_R[253][9];				r_cell_reg[507] = inform_R[765][9];				r_cell_reg[508] = inform_R[254][9];				r_cell_reg[509] = inform_R[766][9];				r_cell_reg[510] = inform_R[255][9];				r_cell_reg[511] = inform_R[767][9];				r_cell_reg[512] = inform_R[256][9];				r_cell_reg[513] = inform_R[768][9];				r_cell_reg[514] = inform_R[257][9];				r_cell_reg[515] = inform_R[769][9];				r_cell_reg[516] = inform_R[258][9];				r_cell_reg[517] = inform_R[770][9];				r_cell_reg[518] = inform_R[259][9];				r_cell_reg[519] = inform_R[771][9];				r_cell_reg[520] = inform_R[260][9];				r_cell_reg[521] = inform_R[772][9];				r_cell_reg[522] = inform_R[261][9];				r_cell_reg[523] = inform_R[773][9];				r_cell_reg[524] = inform_R[262][9];				r_cell_reg[525] = inform_R[774][9];				r_cell_reg[526] = inform_R[263][9];				r_cell_reg[527] = inform_R[775][9];				r_cell_reg[528] = inform_R[264][9];				r_cell_reg[529] = inform_R[776][9];				r_cell_reg[530] = inform_R[265][9];				r_cell_reg[531] = inform_R[777][9];				r_cell_reg[532] = inform_R[266][9];				r_cell_reg[533] = inform_R[778][9];				r_cell_reg[534] = inform_R[267][9];				r_cell_reg[535] = inform_R[779][9];				r_cell_reg[536] = inform_R[268][9];				r_cell_reg[537] = inform_R[780][9];				r_cell_reg[538] = inform_R[269][9];				r_cell_reg[539] = inform_R[781][9];				r_cell_reg[540] = inform_R[270][9];				r_cell_reg[541] = inform_R[782][9];				r_cell_reg[542] = inform_R[271][9];				r_cell_reg[543] = inform_R[783][9];				r_cell_reg[544] = inform_R[272][9];				r_cell_reg[545] = inform_R[784][9];				r_cell_reg[546] = inform_R[273][9];				r_cell_reg[547] = inform_R[785][9];				r_cell_reg[548] = inform_R[274][9];				r_cell_reg[549] = inform_R[786][9];				r_cell_reg[550] = inform_R[275][9];				r_cell_reg[551] = inform_R[787][9];				r_cell_reg[552] = inform_R[276][9];				r_cell_reg[553] = inform_R[788][9];				r_cell_reg[554] = inform_R[277][9];				r_cell_reg[555] = inform_R[789][9];				r_cell_reg[556] = inform_R[278][9];				r_cell_reg[557] = inform_R[790][9];				r_cell_reg[558] = inform_R[279][9];				r_cell_reg[559] = inform_R[791][9];				r_cell_reg[560] = inform_R[280][9];				r_cell_reg[561] = inform_R[792][9];				r_cell_reg[562] = inform_R[281][9];				r_cell_reg[563] = inform_R[793][9];				r_cell_reg[564] = inform_R[282][9];				r_cell_reg[565] = inform_R[794][9];				r_cell_reg[566] = inform_R[283][9];				r_cell_reg[567] = inform_R[795][9];				r_cell_reg[568] = inform_R[284][9];				r_cell_reg[569] = inform_R[796][9];				r_cell_reg[570] = inform_R[285][9];				r_cell_reg[571] = inform_R[797][9];				r_cell_reg[572] = inform_R[286][9];				r_cell_reg[573] = inform_R[798][9];				r_cell_reg[574] = inform_R[287][9];				r_cell_reg[575] = inform_R[799][9];				r_cell_reg[576] = inform_R[288][9];				r_cell_reg[577] = inform_R[800][9];				r_cell_reg[578] = inform_R[289][9];				r_cell_reg[579] = inform_R[801][9];				r_cell_reg[580] = inform_R[290][9];				r_cell_reg[581] = inform_R[802][9];				r_cell_reg[582] = inform_R[291][9];				r_cell_reg[583] = inform_R[803][9];				r_cell_reg[584] = inform_R[292][9];				r_cell_reg[585] = inform_R[804][9];				r_cell_reg[586] = inform_R[293][9];				r_cell_reg[587] = inform_R[805][9];				r_cell_reg[588] = inform_R[294][9];				r_cell_reg[589] = inform_R[806][9];				r_cell_reg[590] = inform_R[295][9];				r_cell_reg[591] = inform_R[807][9];				r_cell_reg[592] = inform_R[296][9];				r_cell_reg[593] = inform_R[808][9];				r_cell_reg[594] = inform_R[297][9];				r_cell_reg[595] = inform_R[809][9];				r_cell_reg[596] = inform_R[298][9];				r_cell_reg[597] = inform_R[810][9];				r_cell_reg[598] = inform_R[299][9];				r_cell_reg[599] = inform_R[811][9];				r_cell_reg[600] = inform_R[300][9];				r_cell_reg[601] = inform_R[812][9];				r_cell_reg[602] = inform_R[301][9];				r_cell_reg[603] = inform_R[813][9];				r_cell_reg[604] = inform_R[302][9];				r_cell_reg[605] = inform_R[814][9];				r_cell_reg[606] = inform_R[303][9];				r_cell_reg[607] = inform_R[815][9];				r_cell_reg[608] = inform_R[304][9];				r_cell_reg[609] = inform_R[816][9];				r_cell_reg[610] = inform_R[305][9];				r_cell_reg[611] = inform_R[817][9];				r_cell_reg[612] = inform_R[306][9];				r_cell_reg[613] = inform_R[818][9];				r_cell_reg[614] = inform_R[307][9];				r_cell_reg[615] = inform_R[819][9];				r_cell_reg[616] = inform_R[308][9];				r_cell_reg[617] = inform_R[820][9];				r_cell_reg[618] = inform_R[309][9];				r_cell_reg[619] = inform_R[821][9];				r_cell_reg[620] = inform_R[310][9];				r_cell_reg[621] = inform_R[822][9];				r_cell_reg[622] = inform_R[311][9];				r_cell_reg[623] = inform_R[823][9];				r_cell_reg[624] = inform_R[312][9];				r_cell_reg[625] = inform_R[824][9];				r_cell_reg[626] = inform_R[313][9];				r_cell_reg[627] = inform_R[825][9];				r_cell_reg[628] = inform_R[314][9];				r_cell_reg[629] = inform_R[826][9];				r_cell_reg[630] = inform_R[315][9];				r_cell_reg[631] = inform_R[827][9];				r_cell_reg[632] = inform_R[316][9];				r_cell_reg[633] = inform_R[828][9];				r_cell_reg[634] = inform_R[317][9];				r_cell_reg[635] = inform_R[829][9];				r_cell_reg[636] = inform_R[318][9];				r_cell_reg[637] = inform_R[830][9];				r_cell_reg[638] = inform_R[319][9];				r_cell_reg[639] = inform_R[831][9];				r_cell_reg[640] = inform_R[320][9];				r_cell_reg[641] = inform_R[832][9];				r_cell_reg[642] = inform_R[321][9];				r_cell_reg[643] = inform_R[833][9];				r_cell_reg[644] = inform_R[322][9];				r_cell_reg[645] = inform_R[834][9];				r_cell_reg[646] = inform_R[323][9];				r_cell_reg[647] = inform_R[835][9];				r_cell_reg[648] = inform_R[324][9];				r_cell_reg[649] = inform_R[836][9];				r_cell_reg[650] = inform_R[325][9];				r_cell_reg[651] = inform_R[837][9];				r_cell_reg[652] = inform_R[326][9];				r_cell_reg[653] = inform_R[838][9];				r_cell_reg[654] = inform_R[327][9];				r_cell_reg[655] = inform_R[839][9];				r_cell_reg[656] = inform_R[328][9];				r_cell_reg[657] = inform_R[840][9];				r_cell_reg[658] = inform_R[329][9];				r_cell_reg[659] = inform_R[841][9];				r_cell_reg[660] = inform_R[330][9];				r_cell_reg[661] = inform_R[842][9];				r_cell_reg[662] = inform_R[331][9];				r_cell_reg[663] = inform_R[843][9];				r_cell_reg[664] = inform_R[332][9];				r_cell_reg[665] = inform_R[844][9];				r_cell_reg[666] = inform_R[333][9];				r_cell_reg[667] = inform_R[845][9];				r_cell_reg[668] = inform_R[334][9];				r_cell_reg[669] = inform_R[846][9];				r_cell_reg[670] = inform_R[335][9];				r_cell_reg[671] = inform_R[847][9];				r_cell_reg[672] = inform_R[336][9];				r_cell_reg[673] = inform_R[848][9];				r_cell_reg[674] = inform_R[337][9];				r_cell_reg[675] = inform_R[849][9];				r_cell_reg[676] = inform_R[338][9];				r_cell_reg[677] = inform_R[850][9];				r_cell_reg[678] = inform_R[339][9];				r_cell_reg[679] = inform_R[851][9];				r_cell_reg[680] = inform_R[340][9];				r_cell_reg[681] = inform_R[852][9];				r_cell_reg[682] = inform_R[341][9];				r_cell_reg[683] = inform_R[853][9];				r_cell_reg[684] = inform_R[342][9];				r_cell_reg[685] = inform_R[854][9];				r_cell_reg[686] = inform_R[343][9];				r_cell_reg[687] = inform_R[855][9];				r_cell_reg[688] = inform_R[344][9];				r_cell_reg[689] = inform_R[856][9];				r_cell_reg[690] = inform_R[345][9];				r_cell_reg[691] = inform_R[857][9];				r_cell_reg[692] = inform_R[346][9];				r_cell_reg[693] = inform_R[858][9];				r_cell_reg[694] = inform_R[347][9];				r_cell_reg[695] = inform_R[859][9];				r_cell_reg[696] = inform_R[348][9];				r_cell_reg[697] = inform_R[860][9];				r_cell_reg[698] = inform_R[349][9];				r_cell_reg[699] = inform_R[861][9];				r_cell_reg[700] = inform_R[350][9];				r_cell_reg[701] = inform_R[862][9];				r_cell_reg[702] = inform_R[351][9];				r_cell_reg[703] = inform_R[863][9];				r_cell_reg[704] = inform_R[352][9];				r_cell_reg[705] = inform_R[864][9];				r_cell_reg[706] = inform_R[353][9];				r_cell_reg[707] = inform_R[865][9];				r_cell_reg[708] = inform_R[354][9];				r_cell_reg[709] = inform_R[866][9];				r_cell_reg[710] = inform_R[355][9];				r_cell_reg[711] = inform_R[867][9];				r_cell_reg[712] = inform_R[356][9];				r_cell_reg[713] = inform_R[868][9];				r_cell_reg[714] = inform_R[357][9];				r_cell_reg[715] = inform_R[869][9];				r_cell_reg[716] = inform_R[358][9];				r_cell_reg[717] = inform_R[870][9];				r_cell_reg[718] = inform_R[359][9];				r_cell_reg[719] = inform_R[871][9];				r_cell_reg[720] = inform_R[360][9];				r_cell_reg[721] = inform_R[872][9];				r_cell_reg[722] = inform_R[361][9];				r_cell_reg[723] = inform_R[873][9];				r_cell_reg[724] = inform_R[362][9];				r_cell_reg[725] = inform_R[874][9];				r_cell_reg[726] = inform_R[363][9];				r_cell_reg[727] = inform_R[875][9];				r_cell_reg[728] = inform_R[364][9];				r_cell_reg[729] = inform_R[876][9];				r_cell_reg[730] = inform_R[365][9];				r_cell_reg[731] = inform_R[877][9];				r_cell_reg[732] = inform_R[366][9];				r_cell_reg[733] = inform_R[878][9];				r_cell_reg[734] = inform_R[367][9];				r_cell_reg[735] = inform_R[879][9];				r_cell_reg[736] = inform_R[368][9];				r_cell_reg[737] = inform_R[880][9];				r_cell_reg[738] = inform_R[369][9];				r_cell_reg[739] = inform_R[881][9];				r_cell_reg[740] = inform_R[370][9];				r_cell_reg[741] = inform_R[882][9];				r_cell_reg[742] = inform_R[371][9];				r_cell_reg[743] = inform_R[883][9];				r_cell_reg[744] = inform_R[372][9];				r_cell_reg[745] = inform_R[884][9];				r_cell_reg[746] = inform_R[373][9];				r_cell_reg[747] = inform_R[885][9];				r_cell_reg[748] = inform_R[374][9];				r_cell_reg[749] = inform_R[886][9];				r_cell_reg[750] = inform_R[375][9];				r_cell_reg[751] = inform_R[887][9];				r_cell_reg[752] = inform_R[376][9];				r_cell_reg[753] = inform_R[888][9];				r_cell_reg[754] = inform_R[377][9];				r_cell_reg[755] = inform_R[889][9];				r_cell_reg[756] = inform_R[378][9];				r_cell_reg[757] = inform_R[890][9];				r_cell_reg[758] = inform_R[379][9];				r_cell_reg[759] = inform_R[891][9];				r_cell_reg[760] = inform_R[380][9];				r_cell_reg[761] = inform_R[892][9];				r_cell_reg[762] = inform_R[381][9];				r_cell_reg[763] = inform_R[893][9];				r_cell_reg[764] = inform_R[382][9];				r_cell_reg[765] = inform_R[894][9];				r_cell_reg[766] = inform_R[383][9];				r_cell_reg[767] = inform_R[895][9];				r_cell_reg[768] = inform_R[384][9];				r_cell_reg[769] = inform_R[896][9];				r_cell_reg[770] = inform_R[385][9];				r_cell_reg[771] = inform_R[897][9];				r_cell_reg[772] = inform_R[386][9];				r_cell_reg[773] = inform_R[898][9];				r_cell_reg[774] = inform_R[387][9];				r_cell_reg[775] = inform_R[899][9];				r_cell_reg[776] = inform_R[388][9];				r_cell_reg[777] = inform_R[900][9];				r_cell_reg[778] = inform_R[389][9];				r_cell_reg[779] = inform_R[901][9];				r_cell_reg[780] = inform_R[390][9];				r_cell_reg[781] = inform_R[902][9];				r_cell_reg[782] = inform_R[391][9];				r_cell_reg[783] = inform_R[903][9];				r_cell_reg[784] = inform_R[392][9];				r_cell_reg[785] = inform_R[904][9];				r_cell_reg[786] = inform_R[393][9];				r_cell_reg[787] = inform_R[905][9];				r_cell_reg[788] = inform_R[394][9];				r_cell_reg[789] = inform_R[906][9];				r_cell_reg[790] = inform_R[395][9];				r_cell_reg[791] = inform_R[907][9];				r_cell_reg[792] = inform_R[396][9];				r_cell_reg[793] = inform_R[908][9];				r_cell_reg[794] = inform_R[397][9];				r_cell_reg[795] = inform_R[909][9];				r_cell_reg[796] = inform_R[398][9];				r_cell_reg[797] = inform_R[910][9];				r_cell_reg[798] = inform_R[399][9];				r_cell_reg[799] = inform_R[911][9];				r_cell_reg[800] = inform_R[400][9];				r_cell_reg[801] = inform_R[912][9];				r_cell_reg[802] = inform_R[401][9];				r_cell_reg[803] = inform_R[913][9];				r_cell_reg[804] = inform_R[402][9];				r_cell_reg[805] = inform_R[914][9];				r_cell_reg[806] = inform_R[403][9];				r_cell_reg[807] = inform_R[915][9];				r_cell_reg[808] = inform_R[404][9];				r_cell_reg[809] = inform_R[916][9];				r_cell_reg[810] = inform_R[405][9];				r_cell_reg[811] = inform_R[917][9];				r_cell_reg[812] = inform_R[406][9];				r_cell_reg[813] = inform_R[918][9];				r_cell_reg[814] = inform_R[407][9];				r_cell_reg[815] = inform_R[919][9];				r_cell_reg[816] = inform_R[408][9];				r_cell_reg[817] = inform_R[920][9];				r_cell_reg[818] = inform_R[409][9];				r_cell_reg[819] = inform_R[921][9];				r_cell_reg[820] = inform_R[410][9];				r_cell_reg[821] = inform_R[922][9];				r_cell_reg[822] = inform_R[411][9];				r_cell_reg[823] = inform_R[923][9];				r_cell_reg[824] = inform_R[412][9];				r_cell_reg[825] = inform_R[924][9];				r_cell_reg[826] = inform_R[413][9];				r_cell_reg[827] = inform_R[925][9];				r_cell_reg[828] = inform_R[414][9];				r_cell_reg[829] = inform_R[926][9];				r_cell_reg[830] = inform_R[415][9];				r_cell_reg[831] = inform_R[927][9];				r_cell_reg[832] = inform_R[416][9];				r_cell_reg[833] = inform_R[928][9];				r_cell_reg[834] = inform_R[417][9];				r_cell_reg[835] = inform_R[929][9];				r_cell_reg[836] = inform_R[418][9];				r_cell_reg[837] = inform_R[930][9];				r_cell_reg[838] = inform_R[419][9];				r_cell_reg[839] = inform_R[931][9];				r_cell_reg[840] = inform_R[420][9];				r_cell_reg[841] = inform_R[932][9];				r_cell_reg[842] = inform_R[421][9];				r_cell_reg[843] = inform_R[933][9];				r_cell_reg[844] = inform_R[422][9];				r_cell_reg[845] = inform_R[934][9];				r_cell_reg[846] = inform_R[423][9];				r_cell_reg[847] = inform_R[935][9];				r_cell_reg[848] = inform_R[424][9];				r_cell_reg[849] = inform_R[936][9];				r_cell_reg[850] = inform_R[425][9];				r_cell_reg[851] = inform_R[937][9];				r_cell_reg[852] = inform_R[426][9];				r_cell_reg[853] = inform_R[938][9];				r_cell_reg[854] = inform_R[427][9];				r_cell_reg[855] = inform_R[939][9];				r_cell_reg[856] = inform_R[428][9];				r_cell_reg[857] = inform_R[940][9];				r_cell_reg[858] = inform_R[429][9];				r_cell_reg[859] = inform_R[941][9];				r_cell_reg[860] = inform_R[430][9];				r_cell_reg[861] = inform_R[942][9];				r_cell_reg[862] = inform_R[431][9];				r_cell_reg[863] = inform_R[943][9];				r_cell_reg[864] = inform_R[432][9];				r_cell_reg[865] = inform_R[944][9];				r_cell_reg[866] = inform_R[433][9];				r_cell_reg[867] = inform_R[945][9];				r_cell_reg[868] = inform_R[434][9];				r_cell_reg[869] = inform_R[946][9];				r_cell_reg[870] = inform_R[435][9];				r_cell_reg[871] = inform_R[947][9];				r_cell_reg[872] = inform_R[436][9];				r_cell_reg[873] = inform_R[948][9];				r_cell_reg[874] = inform_R[437][9];				r_cell_reg[875] = inform_R[949][9];				r_cell_reg[876] = inform_R[438][9];				r_cell_reg[877] = inform_R[950][9];				r_cell_reg[878] = inform_R[439][9];				r_cell_reg[879] = inform_R[951][9];				r_cell_reg[880] = inform_R[440][9];				r_cell_reg[881] = inform_R[952][9];				r_cell_reg[882] = inform_R[441][9];				r_cell_reg[883] = inform_R[953][9];				r_cell_reg[884] = inform_R[442][9];				r_cell_reg[885] = inform_R[954][9];				r_cell_reg[886] = inform_R[443][9];				r_cell_reg[887] = inform_R[955][9];				r_cell_reg[888] = inform_R[444][9];				r_cell_reg[889] = inform_R[956][9];				r_cell_reg[890] = inform_R[445][9];				r_cell_reg[891] = inform_R[957][9];				r_cell_reg[892] = inform_R[446][9];				r_cell_reg[893] = inform_R[958][9];				r_cell_reg[894] = inform_R[447][9];				r_cell_reg[895] = inform_R[959][9];				r_cell_reg[896] = inform_R[448][9];				r_cell_reg[897] = inform_R[960][9];				r_cell_reg[898] = inform_R[449][9];				r_cell_reg[899] = inform_R[961][9];				r_cell_reg[900] = inform_R[450][9];				r_cell_reg[901] = inform_R[962][9];				r_cell_reg[902] = inform_R[451][9];				r_cell_reg[903] = inform_R[963][9];				r_cell_reg[904] = inform_R[452][9];				r_cell_reg[905] = inform_R[964][9];				r_cell_reg[906] = inform_R[453][9];				r_cell_reg[907] = inform_R[965][9];				r_cell_reg[908] = inform_R[454][9];				r_cell_reg[909] = inform_R[966][9];				r_cell_reg[910] = inform_R[455][9];				r_cell_reg[911] = inform_R[967][9];				r_cell_reg[912] = inform_R[456][9];				r_cell_reg[913] = inform_R[968][9];				r_cell_reg[914] = inform_R[457][9];				r_cell_reg[915] = inform_R[969][9];				r_cell_reg[916] = inform_R[458][9];				r_cell_reg[917] = inform_R[970][9];				r_cell_reg[918] = inform_R[459][9];				r_cell_reg[919] = inform_R[971][9];				r_cell_reg[920] = inform_R[460][9];				r_cell_reg[921] = inform_R[972][9];				r_cell_reg[922] = inform_R[461][9];				r_cell_reg[923] = inform_R[973][9];				r_cell_reg[924] = inform_R[462][9];				r_cell_reg[925] = inform_R[974][9];				r_cell_reg[926] = inform_R[463][9];				r_cell_reg[927] = inform_R[975][9];				r_cell_reg[928] = inform_R[464][9];				r_cell_reg[929] = inform_R[976][9];				r_cell_reg[930] = inform_R[465][9];				r_cell_reg[931] = inform_R[977][9];				r_cell_reg[932] = inform_R[466][9];				r_cell_reg[933] = inform_R[978][9];				r_cell_reg[934] = inform_R[467][9];				r_cell_reg[935] = inform_R[979][9];				r_cell_reg[936] = inform_R[468][9];				r_cell_reg[937] = inform_R[980][9];				r_cell_reg[938] = inform_R[469][9];				r_cell_reg[939] = inform_R[981][9];				r_cell_reg[940] = inform_R[470][9];				r_cell_reg[941] = inform_R[982][9];				r_cell_reg[942] = inform_R[471][9];				r_cell_reg[943] = inform_R[983][9];				r_cell_reg[944] = inform_R[472][9];				r_cell_reg[945] = inform_R[984][9];				r_cell_reg[946] = inform_R[473][9];				r_cell_reg[947] = inform_R[985][9];				r_cell_reg[948] = inform_R[474][9];				r_cell_reg[949] = inform_R[986][9];				r_cell_reg[950] = inform_R[475][9];				r_cell_reg[951] = inform_R[987][9];				r_cell_reg[952] = inform_R[476][9];				r_cell_reg[953] = inform_R[988][9];				r_cell_reg[954] = inform_R[477][9];				r_cell_reg[955] = inform_R[989][9];				r_cell_reg[956] = inform_R[478][9];				r_cell_reg[957] = inform_R[990][9];				r_cell_reg[958] = inform_R[479][9];				r_cell_reg[959] = inform_R[991][9];				r_cell_reg[960] = inform_R[480][9];				r_cell_reg[961] = inform_R[992][9];				r_cell_reg[962] = inform_R[481][9];				r_cell_reg[963] = inform_R[993][9];				r_cell_reg[964] = inform_R[482][9];				r_cell_reg[965] = inform_R[994][9];				r_cell_reg[966] = inform_R[483][9];				r_cell_reg[967] = inform_R[995][9];				r_cell_reg[968] = inform_R[484][9];				r_cell_reg[969] = inform_R[996][9];				r_cell_reg[970] = inform_R[485][9];				r_cell_reg[971] = inform_R[997][9];				r_cell_reg[972] = inform_R[486][9];				r_cell_reg[973] = inform_R[998][9];				r_cell_reg[974] = inform_R[487][9];				r_cell_reg[975] = inform_R[999][9];				r_cell_reg[976] = inform_R[488][9];				r_cell_reg[977] = inform_R[1000][9];				r_cell_reg[978] = inform_R[489][9];				r_cell_reg[979] = inform_R[1001][9];				r_cell_reg[980] = inform_R[490][9];				r_cell_reg[981] = inform_R[1002][9];				r_cell_reg[982] = inform_R[491][9];				r_cell_reg[983] = inform_R[1003][9];				r_cell_reg[984] = inform_R[492][9];				r_cell_reg[985] = inform_R[1004][9];				r_cell_reg[986] = inform_R[493][9];				r_cell_reg[987] = inform_R[1005][9];				r_cell_reg[988] = inform_R[494][9];				r_cell_reg[989] = inform_R[1006][9];				r_cell_reg[990] = inform_R[495][9];				r_cell_reg[991] = inform_R[1007][9];				r_cell_reg[992] = inform_R[496][9];				r_cell_reg[993] = inform_R[1008][9];				r_cell_reg[994] = inform_R[497][9];				r_cell_reg[995] = inform_R[1009][9];				r_cell_reg[996] = inform_R[498][9];				r_cell_reg[997] = inform_R[1010][9];				r_cell_reg[998] = inform_R[499][9];				r_cell_reg[999] = inform_R[1011][9];				r_cell_reg[1000] = inform_R[500][9];				r_cell_reg[1001] = inform_R[1012][9];				r_cell_reg[1002] = inform_R[501][9];				r_cell_reg[1003] = inform_R[1013][9];				r_cell_reg[1004] = inform_R[502][9];				r_cell_reg[1005] = inform_R[1014][9];				r_cell_reg[1006] = inform_R[503][9];				r_cell_reg[1007] = inform_R[1015][9];				r_cell_reg[1008] = inform_R[504][9];				r_cell_reg[1009] = inform_R[1016][9];				r_cell_reg[1010] = inform_R[505][9];				r_cell_reg[1011] = inform_R[1017][9];				r_cell_reg[1012] = inform_R[506][9];				r_cell_reg[1013] = inform_R[1018][9];				r_cell_reg[1014] = inform_R[507][9];				r_cell_reg[1015] = inform_R[1019][9];				r_cell_reg[1016] = inform_R[508][9];				r_cell_reg[1017] = inform_R[1020][9];				r_cell_reg[1018] = inform_R[509][9];				r_cell_reg[1019] = inform_R[1021][9];				r_cell_reg[1020] = inform_R[510][9];				r_cell_reg[1021] = inform_R[1022][9];				r_cell_reg[1022] = inform_R[511][9];				r_cell_reg[1023] = inform_R[1023][9];				l_cell_reg[0] = inform_L[0][10];				l_cell_reg[1] = inform_L[512][10];				l_cell_reg[2] = inform_L[1][10];				l_cell_reg[3] = inform_L[513][10];				l_cell_reg[4] = inform_L[2][10];				l_cell_reg[5] = inform_L[514][10];				l_cell_reg[6] = inform_L[3][10];				l_cell_reg[7] = inform_L[515][10];				l_cell_reg[8] = inform_L[4][10];				l_cell_reg[9] = inform_L[516][10];				l_cell_reg[10] = inform_L[5][10];				l_cell_reg[11] = inform_L[517][10];				l_cell_reg[12] = inform_L[6][10];				l_cell_reg[13] = inform_L[518][10];				l_cell_reg[14] = inform_L[7][10];				l_cell_reg[15] = inform_L[519][10];				l_cell_reg[16] = inform_L[8][10];				l_cell_reg[17] = inform_L[520][10];				l_cell_reg[18] = inform_L[9][10];				l_cell_reg[19] = inform_L[521][10];				l_cell_reg[20] = inform_L[10][10];				l_cell_reg[21] = inform_L[522][10];				l_cell_reg[22] = inform_L[11][10];				l_cell_reg[23] = inform_L[523][10];				l_cell_reg[24] = inform_L[12][10];				l_cell_reg[25] = inform_L[524][10];				l_cell_reg[26] = inform_L[13][10];				l_cell_reg[27] = inform_L[525][10];				l_cell_reg[28] = inform_L[14][10];				l_cell_reg[29] = inform_L[526][10];				l_cell_reg[30] = inform_L[15][10];				l_cell_reg[31] = inform_L[527][10];				l_cell_reg[32] = inform_L[16][10];				l_cell_reg[33] = inform_L[528][10];				l_cell_reg[34] = inform_L[17][10];				l_cell_reg[35] = inform_L[529][10];				l_cell_reg[36] = inform_L[18][10];				l_cell_reg[37] = inform_L[530][10];				l_cell_reg[38] = inform_L[19][10];				l_cell_reg[39] = inform_L[531][10];				l_cell_reg[40] = inform_L[20][10];				l_cell_reg[41] = inform_L[532][10];				l_cell_reg[42] = inform_L[21][10];				l_cell_reg[43] = inform_L[533][10];				l_cell_reg[44] = inform_L[22][10];				l_cell_reg[45] = inform_L[534][10];				l_cell_reg[46] = inform_L[23][10];				l_cell_reg[47] = inform_L[535][10];				l_cell_reg[48] = inform_L[24][10];				l_cell_reg[49] = inform_L[536][10];				l_cell_reg[50] = inform_L[25][10];				l_cell_reg[51] = inform_L[537][10];				l_cell_reg[52] = inform_L[26][10];				l_cell_reg[53] = inform_L[538][10];				l_cell_reg[54] = inform_L[27][10];				l_cell_reg[55] = inform_L[539][10];				l_cell_reg[56] = inform_L[28][10];				l_cell_reg[57] = inform_L[540][10];				l_cell_reg[58] = inform_L[29][10];				l_cell_reg[59] = inform_L[541][10];				l_cell_reg[60] = inform_L[30][10];				l_cell_reg[61] = inform_L[542][10];				l_cell_reg[62] = inform_L[31][10];				l_cell_reg[63] = inform_L[543][10];				l_cell_reg[64] = inform_L[32][10];				l_cell_reg[65] = inform_L[544][10];				l_cell_reg[66] = inform_L[33][10];				l_cell_reg[67] = inform_L[545][10];				l_cell_reg[68] = inform_L[34][10];				l_cell_reg[69] = inform_L[546][10];				l_cell_reg[70] = inform_L[35][10];				l_cell_reg[71] = inform_L[547][10];				l_cell_reg[72] = inform_L[36][10];				l_cell_reg[73] = inform_L[548][10];				l_cell_reg[74] = inform_L[37][10];				l_cell_reg[75] = inform_L[549][10];				l_cell_reg[76] = inform_L[38][10];				l_cell_reg[77] = inform_L[550][10];				l_cell_reg[78] = inform_L[39][10];				l_cell_reg[79] = inform_L[551][10];				l_cell_reg[80] = inform_L[40][10];				l_cell_reg[81] = inform_L[552][10];				l_cell_reg[82] = inform_L[41][10];				l_cell_reg[83] = inform_L[553][10];				l_cell_reg[84] = inform_L[42][10];				l_cell_reg[85] = inform_L[554][10];				l_cell_reg[86] = inform_L[43][10];				l_cell_reg[87] = inform_L[555][10];				l_cell_reg[88] = inform_L[44][10];				l_cell_reg[89] = inform_L[556][10];				l_cell_reg[90] = inform_L[45][10];				l_cell_reg[91] = inform_L[557][10];				l_cell_reg[92] = inform_L[46][10];				l_cell_reg[93] = inform_L[558][10];				l_cell_reg[94] = inform_L[47][10];				l_cell_reg[95] = inform_L[559][10];				l_cell_reg[96] = inform_L[48][10];				l_cell_reg[97] = inform_L[560][10];				l_cell_reg[98] = inform_L[49][10];				l_cell_reg[99] = inform_L[561][10];				l_cell_reg[100] = inform_L[50][10];				l_cell_reg[101] = inform_L[562][10];				l_cell_reg[102] = inform_L[51][10];				l_cell_reg[103] = inform_L[563][10];				l_cell_reg[104] = inform_L[52][10];				l_cell_reg[105] = inform_L[564][10];				l_cell_reg[106] = inform_L[53][10];				l_cell_reg[107] = inform_L[565][10];				l_cell_reg[108] = inform_L[54][10];				l_cell_reg[109] = inform_L[566][10];				l_cell_reg[110] = inform_L[55][10];				l_cell_reg[111] = inform_L[567][10];				l_cell_reg[112] = inform_L[56][10];				l_cell_reg[113] = inform_L[568][10];				l_cell_reg[114] = inform_L[57][10];				l_cell_reg[115] = inform_L[569][10];				l_cell_reg[116] = inform_L[58][10];				l_cell_reg[117] = inform_L[570][10];				l_cell_reg[118] = inform_L[59][10];				l_cell_reg[119] = inform_L[571][10];				l_cell_reg[120] = inform_L[60][10];				l_cell_reg[121] = inform_L[572][10];				l_cell_reg[122] = inform_L[61][10];				l_cell_reg[123] = inform_L[573][10];				l_cell_reg[124] = inform_L[62][10];				l_cell_reg[125] = inform_L[574][10];				l_cell_reg[126] = inform_L[63][10];				l_cell_reg[127] = inform_L[575][10];				l_cell_reg[128] = inform_L[64][10];				l_cell_reg[129] = inform_L[576][10];				l_cell_reg[130] = inform_L[65][10];				l_cell_reg[131] = inform_L[577][10];				l_cell_reg[132] = inform_L[66][10];				l_cell_reg[133] = inform_L[578][10];				l_cell_reg[134] = inform_L[67][10];				l_cell_reg[135] = inform_L[579][10];				l_cell_reg[136] = inform_L[68][10];				l_cell_reg[137] = inform_L[580][10];				l_cell_reg[138] = inform_L[69][10];				l_cell_reg[139] = inform_L[581][10];				l_cell_reg[140] = inform_L[70][10];				l_cell_reg[141] = inform_L[582][10];				l_cell_reg[142] = inform_L[71][10];				l_cell_reg[143] = inform_L[583][10];				l_cell_reg[144] = inform_L[72][10];				l_cell_reg[145] = inform_L[584][10];				l_cell_reg[146] = inform_L[73][10];				l_cell_reg[147] = inform_L[585][10];				l_cell_reg[148] = inform_L[74][10];				l_cell_reg[149] = inform_L[586][10];				l_cell_reg[150] = inform_L[75][10];				l_cell_reg[151] = inform_L[587][10];				l_cell_reg[152] = inform_L[76][10];				l_cell_reg[153] = inform_L[588][10];				l_cell_reg[154] = inform_L[77][10];				l_cell_reg[155] = inform_L[589][10];				l_cell_reg[156] = inform_L[78][10];				l_cell_reg[157] = inform_L[590][10];				l_cell_reg[158] = inform_L[79][10];				l_cell_reg[159] = inform_L[591][10];				l_cell_reg[160] = inform_L[80][10];				l_cell_reg[161] = inform_L[592][10];				l_cell_reg[162] = inform_L[81][10];				l_cell_reg[163] = inform_L[593][10];				l_cell_reg[164] = inform_L[82][10];				l_cell_reg[165] = inform_L[594][10];				l_cell_reg[166] = inform_L[83][10];				l_cell_reg[167] = inform_L[595][10];				l_cell_reg[168] = inform_L[84][10];				l_cell_reg[169] = inform_L[596][10];				l_cell_reg[170] = inform_L[85][10];				l_cell_reg[171] = inform_L[597][10];				l_cell_reg[172] = inform_L[86][10];				l_cell_reg[173] = inform_L[598][10];				l_cell_reg[174] = inform_L[87][10];				l_cell_reg[175] = inform_L[599][10];				l_cell_reg[176] = inform_L[88][10];				l_cell_reg[177] = inform_L[600][10];				l_cell_reg[178] = inform_L[89][10];				l_cell_reg[179] = inform_L[601][10];				l_cell_reg[180] = inform_L[90][10];				l_cell_reg[181] = inform_L[602][10];				l_cell_reg[182] = inform_L[91][10];				l_cell_reg[183] = inform_L[603][10];				l_cell_reg[184] = inform_L[92][10];				l_cell_reg[185] = inform_L[604][10];				l_cell_reg[186] = inform_L[93][10];				l_cell_reg[187] = inform_L[605][10];				l_cell_reg[188] = inform_L[94][10];				l_cell_reg[189] = inform_L[606][10];				l_cell_reg[190] = inform_L[95][10];				l_cell_reg[191] = inform_L[607][10];				l_cell_reg[192] = inform_L[96][10];				l_cell_reg[193] = inform_L[608][10];				l_cell_reg[194] = inform_L[97][10];				l_cell_reg[195] = inform_L[609][10];				l_cell_reg[196] = inform_L[98][10];				l_cell_reg[197] = inform_L[610][10];				l_cell_reg[198] = inform_L[99][10];				l_cell_reg[199] = inform_L[611][10];				l_cell_reg[200] = inform_L[100][10];				l_cell_reg[201] = inform_L[612][10];				l_cell_reg[202] = inform_L[101][10];				l_cell_reg[203] = inform_L[613][10];				l_cell_reg[204] = inform_L[102][10];				l_cell_reg[205] = inform_L[614][10];				l_cell_reg[206] = inform_L[103][10];				l_cell_reg[207] = inform_L[615][10];				l_cell_reg[208] = inform_L[104][10];				l_cell_reg[209] = inform_L[616][10];				l_cell_reg[210] = inform_L[105][10];				l_cell_reg[211] = inform_L[617][10];				l_cell_reg[212] = inform_L[106][10];				l_cell_reg[213] = inform_L[618][10];				l_cell_reg[214] = inform_L[107][10];				l_cell_reg[215] = inform_L[619][10];				l_cell_reg[216] = inform_L[108][10];				l_cell_reg[217] = inform_L[620][10];				l_cell_reg[218] = inform_L[109][10];				l_cell_reg[219] = inform_L[621][10];				l_cell_reg[220] = inform_L[110][10];				l_cell_reg[221] = inform_L[622][10];				l_cell_reg[222] = inform_L[111][10];				l_cell_reg[223] = inform_L[623][10];				l_cell_reg[224] = inform_L[112][10];				l_cell_reg[225] = inform_L[624][10];				l_cell_reg[226] = inform_L[113][10];				l_cell_reg[227] = inform_L[625][10];				l_cell_reg[228] = inform_L[114][10];				l_cell_reg[229] = inform_L[626][10];				l_cell_reg[230] = inform_L[115][10];				l_cell_reg[231] = inform_L[627][10];				l_cell_reg[232] = inform_L[116][10];				l_cell_reg[233] = inform_L[628][10];				l_cell_reg[234] = inform_L[117][10];				l_cell_reg[235] = inform_L[629][10];				l_cell_reg[236] = inform_L[118][10];				l_cell_reg[237] = inform_L[630][10];				l_cell_reg[238] = inform_L[119][10];				l_cell_reg[239] = inform_L[631][10];				l_cell_reg[240] = inform_L[120][10];				l_cell_reg[241] = inform_L[632][10];				l_cell_reg[242] = inform_L[121][10];				l_cell_reg[243] = inform_L[633][10];				l_cell_reg[244] = inform_L[122][10];				l_cell_reg[245] = inform_L[634][10];				l_cell_reg[246] = inform_L[123][10];				l_cell_reg[247] = inform_L[635][10];				l_cell_reg[248] = inform_L[124][10];				l_cell_reg[249] = inform_L[636][10];				l_cell_reg[250] = inform_L[125][10];				l_cell_reg[251] = inform_L[637][10];				l_cell_reg[252] = inform_L[126][10];				l_cell_reg[253] = inform_L[638][10];				l_cell_reg[254] = inform_L[127][10];				l_cell_reg[255] = inform_L[639][10];				l_cell_reg[256] = inform_L[128][10];				l_cell_reg[257] = inform_L[640][10];				l_cell_reg[258] = inform_L[129][10];				l_cell_reg[259] = inform_L[641][10];				l_cell_reg[260] = inform_L[130][10];				l_cell_reg[261] = inform_L[642][10];				l_cell_reg[262] = inform_L[131][10];				l_cell_reg[263] = inform_L[643][10];				l_cell_reg[264] = inform_L[132][10];				l_cell_reg[265] = inform_L[644][10];				l_cell_reg[266] = inform_L[133][10];				l_cell_reg[267] = inform_L[645][10];				l_cell_reg[268] = inform_L[134][10];				l_cell_reg[269] = inform_L[646][10];				l_cell_reg[270] = inform_L[135][10];				l_cell_reg[271] = inform_L[647][10];				l_cell_reg[272] = inform_L[136][10];				l_cell_reg[273] = inform_L[648][10];				l_cell_reg[274] = inform_L[137][10];				l_cell_reg[275] = inform_L[649][10];				l_cell_reg[276] = inform_L[138][10];				l_cell_reg[277] = inform_L[650][10];				l_cell_reg[278] = inform_L[139][10];				l_cell_reg[279] = inform_L[651][10];				l_cell_reg[280] = inform_L[140][10];				l_cell_reg[281] = inform_L[652][10];				l_cell_reg[282] = inform_L[141][10];				l_cell_reg[283] = inform_L[653][10];				l_cell_reg[284] = inform_L[142][10];				l_cell_reg[285] = inform_L[654][10];				l_cell_reg[286] = inform_L[143][10];				l_cell_reg[287] = inform_L[655][10];				l_cell_reg[288] = inform_L[144][10];				l_cell_reg[289] = inform_L[656][10];				l_cell_reg[290] = inform_L[145][10];				l_cell_reg[291] = inform_L[657][10];				l_cell_reg[292] = inform_L[146][10];				l_cell_reg[293] = inform_L[658][10];				l_cell_reg[294] = inform_L[147][10];				l_cell_reg[295] = inform_L[659][10];				l_cell_reg[296] = inform_L[148][10];				l_cell_reg[297] = inform_L[660][10];				l_cell_reg[298] = inform_L[149][10];				l_cell_reg[299] = inform_L[661][10];				l_cell_reg[300] = inform_L[150][10];				l_cell_reg[301] = inform_L[662][10];				l_cell_reg[302] = inform_L[151][10];				l_cell_reg[303] = inform_L[663][10];				l_cell_reg[304] = inform_L[152][10];				l_cell_reg[305] = inform_L[664][10];				l_cell_reg[306] = inform_L[153][10];				l_cell_reg[307] = inform_L[665][10];				l_cell_reg[308] = inform_L[154][10];				l_cell_reg[309] = inform_L[666][10];				l_cell_reg[310] = inform_L[155][10];				l_cell_reg[311] = inform_L[667][10];				l_cell_reg[312] = inform_L[156][10];				l_cell_reg[313] = inform_L[668][10];				l_cell_reg[314] = inform_L[157][10];				l_cell_reg[315] = inform_L[669][10];				l_cell_reg[316] = inform_L[158][10];				l_cell_reg[317] = inform_L[670][10];				l_cell_reg[318] = inform_L[159][10];				l_cell_reg[319] = inform_L[671][10];				l_cell_reg[320] = inform_L[160][10];				l_cell_reg[321] = inform_L[672][10];				l_cell_reg[322] = inform_L[161][10];				l_cell_reg[323] = inform_L[673][10];				l_cell_reg[324] = inform_L[162][10];				l_cell_reg[325] = inform_L[674][10];				l_cell_reg[326] = inform_L[163][10];				l_cell_reg[327] = inform_L[675][10];				l_cell_reg[328] = inform_L[164][10];				l_cell_reg[329] = inform_L[676][10];				l_cell_reg[330] = inform_L[165][10];				l_cell_reg[331] = inform_L[677][10];				l_cell_reg[332] = inform_L[166][10];				l_cell_reg[333] = inform_L[678][10];				l_cell_reg[334] = inform_L[167][10];				l_cell_reg[335] = inform_L[679][10];				l_cell_reg[336] = inform_L[168][10];				l_cell_reg[337] = inform_L[680][10];				l_cell_reg[338] = inform_L[169][10];				l_cell_reg[339] = inform_L[681][10];				l_cell_reg[340] = inform_L[170][10];				l_cell_reg[341] = inform_L[682][10];				l_cell_reg[342] = inform_L[171][10];				l_cell_reg[343] = inform_L[683][10];				l_cell_reg[344] = inform_L[172][10];				l_cell_reg[345] = inform_L[684][10];				l_cell_reg[346] = inform_L[173][10];				l_cell_reg[347] = inform_L[685][10];				l_cell_reg[348] = inform_L[174][10];				l_cell_reg[349] = inform_L[686][10];				l_cell_reg[350] = inform_L[175][10];				l_cell_reg[351] = inform_L[687][10];				l_cell_reg[352] = inform_L[176][10];				l_cell_reg[353] = inform_L[688][10];				l_cell_reg[354] = inform_L[177][10];				l_cell_reg[355] = inform_L[689][10];				l_cell_reg[356] = inform_L[178][10];				l_cell_reg[357] = inform_L[690][10];				l_cell_reg[358] = inform_L[179][10];				l_cell_reg[359] = inform_L[691][10];				l_cell_reg[360] = inform_L[180][10];				l_cell_reg[361] = inform_L[692][10];				l_cell_reg[362] = inform_L[181][10];				l_cell_reg[363] = inform_L[693][10];				l_cell_reg[364] = inform_L[182][10];				l_cell_reg[365] = inform_L[694][10];				l_cell_reg[366] = inform_L[183][10];				l_cell_reg[367] = inform_L[695][10];				l_cell_reg[368] = inform_L[184][10];				l_cell_reg[369] = inform_L[696][10];				l_cell_reg[370] = inform_L[185][10];				l_cell_reg[371] = inform_L[697][10];				l_cell_reg[372] = inform_L[186][10];				l_cell_reg[373] = inform_L[698][10];				l_cell_reg[374] = inform_L[187][10];				l_cell_reg[375] = inform_L[699][10];				l_cell_reg[376] = inform_L[188][10];				l_cell_reg[377] = inform_L[700][10];				l_cell_reg[378] = inform_L[189][10];				l_cell_reg[379] = inform_L[701][10];				l_cell_reg[380] = inform_L[190][10];				l_cell_reg[381] = inform_L[702][10];				l_cell_reg[382] = inform_L[191][10];				l_cell_reg[383] = inform_L[703][10];				l_cell_reg[384] = inform_L[192][10];				l_cell_reg[385] = inform_L[704][10];				l_cell_reg[386] = inform_L[193][10];				l_cell_reg[387] = inform_L[705][10];				l_cell_reg[388] = inform_L[194][10];				l_cell_reg[389] = inform_L[706][10];				l_cell_reg[390] = inform_L[195][10];				l_cell_reg[391] = inform_L[707][10];				l_cell_reg[392] = inform_L[196][10];				l_cell_reg[393] = inform_L[708][10];				l_cell_reg[394] = inform_L[197][10];				l_cell_reg[395] = inform_L[709][10];				l_cell_reg[396] = inform_L[198][10];				l_cell_reg[397] = inform_L[710][10];				l_cell_reg[398] = inform_L[199][10];				l_cell_reg[399] = inform_L[711][10];				l_cell_reg[400] = inform_L[200][10];				l_cell_reg[401] = inform_L[712][10];				l_cell_reg[402] = inform_L[201][10];				l_cell_reg[403] = inform_L[713][10];				l_cell_reg[404] = inform_L[202][10];				l_cell_reg[405] = inform_L[714][10];				l_cell_reg[406] = inform_L[203][10];				l_cell_reg[407] = inform_L[715][10];				l_cell_reg[408] = inform_L[204][10];				l_cell_reg[409] = inform_L[716][10];				l_cell_reg[410] = inform_L[205][10];				l_cell_reg[411] = inform_L[717][10];				l_cell_reg[412] = inform_L[206][10];				l_cell_reg[413] = inform_L[718][10];				l_cell_reg[414] = inform_L[207][10];				l_cell_reg[415] = inform_L[719][10];				l_cell_reg[416] = inform_L[208][10];				l_cell_reg[417] = inform_L[720][10];				l_cell_reg[418] = inform_L[209][10];				l_cell_reg[419] = inform_L[721][10];				l_cell_reg[420] = inform_L[210][10];				l_cell_reg[421] = inform_L[722][10];				l_cell_reg[422] = inform_L[211][10];				l_cell_reg[423] = inform_L[723][10];				l_cell_reg[424] = inform_L[212][10];				l_cell_reg[425] = inform_L[724][10];				l_cell_reg[426] = inform_L[213][10];				l_cell_reg[427] = inform_L[725][10];				l_cell_reg[428] = inform_L[214][10];				l_cell_reg[429] = inform_L[726][10];				l_cell_reg[430] = inform_L[215][10];				l_cell_reg[431] = inform_L[727][10];				l_cell_reg[432] = inform_L[216][10];				l_cell_reg[433] = inform_L[728][10];				l_cell_reg[434] = inform_L[217][10];				l_cell_reg[435] = inform_L[729][10];				l_cell_reg[436] = inform_L[218][10];				l_cell_reg[437] = inform_L[730][10];				l_cell_reg[438] = inform_L[219][10];				l_cell_reg[439] = inform_L[731][10];				l_cell_reg[440] = inform_L[220][10];				l_cell_reg[441] = inform_L[732][10];				l_cell_reg[442] = inform_L[221][10];				l_cell_reg[443] = inform_L[733][10];				l_cell_reg[444] = inform_L[222][10];				l_cell_reg[445] = inform_L[734][10];				l_cell_reg[446] = inform_L[223][10];				l_cell_reg[447] = inform_L[735][10];				l_cell_reg[448] = inform_L[224][10];				l_cell_reg[449] = inform_L[736][10];				l_cell_reg[450] = inform_L[225][10];				l_cell_reg[451] = inform_L[737][10];				l_cell_reg[452] = inform_L[226][10];				l_cell_reg[453] = inform_L[738][10];				l_cell_reg[454] = inform_L[227][10];				l_cell_reg[455] = inform_L[739][10];				l_cell_reg[456] = inform_L[228][10];				l_cell_reg[457] = inform_L[740][10];				l_cell_reg[458] = inform_L[229][10];				l_cell_reg[459] = inform_L[741][10];				l_cell_reg[460] = inform_L[230][10];				l_cell_reg[461] = inform_L[742][10];				l_cell_reg[462] = inform_L[231][10];				l_cell_reg[463] = inform_L[743][10];				l_cell_reg[464] = inform_L[232][10];				l_cell_reg[465] = inform_L[744][10];				l_cell_reg[466] = inform_L[233][10];				l_cell_reg[467] = inform_L[745][10];				l_cell_reg[468] = inform_L[234][10];				l_cell_reg[469] = inform_L[746][10];				l_cell_reg[470] = inform_L[235][10];				l_cell_reg[471] = inform_L[747][10];				l_cell_reg[472] = inform_L[236][10];				l_cell_reg[473] = inform_L[748][10];				l_cell_reg[474] = inform_L[237][10];				l_cell_reg[475] = inform_L[749][10];				l_cell_reg[476] = inform_L[238][10];				l_cell_reg[477] = inform_L[750][10];				l_cell_reg[478] = inform_L[239][10];				l_cell_reg[479] = inform_L[751][10];				l_cell_reg[480] = inform_L[240][10];				l_cell_reg[481] = inform_L[752][10];				l_cell_reg[482] = inform_L[241][10];				l_cell_reg[483] = inform_L[753][10];				l_cell_reg[484] = inform_L[242][10];				l_cell_reg[485] = inform_L[754][10];				l_cell_reg[486] = inform_L[243][10];				l_cell_reg[487] = inform_L[755][10];				l_cell_reg[488] = inform_L[244][10];				l_cell_reg[489] = inform_L[756][10];				l_cell_reg[490] = inform_L[245][10];				l_cell_reg[491] = inform_L[757][10];				l_cell_reg[492] = inform_L[246][10];				l_cell_reg[493] = inform_L[758][10];				l_cell_reg[494] = inform_L[247][10];				l_cell_reg[495] = inform_L[759][10];				l_cell_reg[496] = inform_L[248][10];				l_cell_reg[497] = inform_L[760][10];				l_cell_reg[498] = inform_L[249][10];				l_cell_reg[499] = inform_L[761][10];				l_cell_reg[500] = inform_L[250][10];				l_cell_reg[501] = inform_L[762][10];				l_cell_reg[502] = inform_L[251][10];				l_cell_reg[503] = inform_L[763][10];				l_cell_reg[504] = inform_L[252][10];				l_cell_reg[505] = inform_L[764][10];				l_cell_reg[506] = inform_L[253][10];				l_cell_reg[507] = inform_L[765][10];				l_cell_reg[508] = inform_L[254][10];				l_cell_reg[509] = inform_L[766][10];				l_cell_reg[510] = inform_L[255][10];				l_cell_reg[511] = inform_L[767][10];				l_cell_reg[512] = inform_L[256][10];				l_cell_reg[513] = inform_L[768][10];				l_cell_reg[514] = inform_L[257][10];				l_cell_reg[515] = inform_L[769][10];				l_cell_reg[516] = inform_L[258][10];				l_cell_reg[517] = inform_L[770][10];				l_cell_reg[518] = inform_L[259][10];				l_cell_reg[519] = inform_L[771][10];				l_cell_reg[520] = inform_L[260][10];				l_cell_reg[521] = inform_L[772][10];				l_cell_reg[522] = inform_L[261][10];				l_cell_reg[523] = inform_L[773][10];				l_cell_reg[524] = inform_L[262][10];				l_cell_reg[525] = inform_L[774][10];				l_cell_reg[526] = inform_L[263][10];				l_cell_reg[527] = inform_L[775][10];				l_cell_reg[528] = inform_L[264][10];				l_cell_reg[529] = inform_L[776][10];				l_cell_reg[530] = inform_L[265][10];				l_cell_reg[531] = inform_L[777][10];				l_cell_reg[532] = inform_L[266][10];				l_cell_reg[533] = inform_L[778][10];				l_cell_reg[534] = inform_L[267][10];				l_cell_reg[535] = inform_L[779][10];				l_cell_reg[536] = inform_L[268][10];				l_cell_reg[537] = inform_L[780][10];				l_cell_reg[538] = inform_L[269][10];				l_cell_reg[539] = inform_L[781][10];				l_cell_reg[540] = inform_L[270][10];				l_cell_reg[541] = inform_L[782][10];				l_cell_reg[542] = inform_L[271][10];				l_cell_reg[543] = inform_L[783][10];				l_cell_reg[544] = inform_L[272][10];				l_cell_reg[545] = inform_L[784][10];				l_cell_reg[546] = inform_L[273][10];				l_cell_reg[547] = inform_L[785][10];				l_cell_reg[548] = inform_L[274][10];				l_cell_reg[549] = inform_L[786][10];				l_cell_reg[550] = inform_L[275][10];				l_cell_reg[551] = inform_L[787][10];				l_cell_reg[552] = inform_L[276][10];				l_cell_reg[553] = inform_L[788][10];				l_cell_reg[554] = inform_L[277][10];				l_cell_reg[555] = inform_L[789][10];				l_cell_reg[556] = inform_L[278][10];				l_cell_reg[557] = inform_L[790][10];				l_cell_reg[558] = inform_L[279][10];				l_cell_reg[559] = inform_L[791][10];				l_cell_reg[560] = inform_L[280][10];				l_cell_reg[561] = inform_L[792][10];				l_cell_reg[562] = inform_L[281][10];				l_cell_reg[563] = inform_L[793][10];				l_cell_reg[564] = inform_L[282][10];				l_cell_reg[565] = inform_L[794][10];				l_cell_reg[566] = inform_L[283][10];				l_cell_reg[567] = inform_L[795][10];				l_cell_reg[568] = inform_L[284][10];				l_cell_reg[569] = inform_L[796][10];				l_cell_reg[570] = inform_L[285][10];				l_cell_reg[571] = inform_L[797][10];				l_cell_reg[572] = inform_L[286][10];				l_cell_reg[573] = inform_L[798][10];				l_cell_reg[574] = inform_L[287][10];				l_cell_reg[575] = inform_L[799][10];				l_cell_reg[576] = inform_L[288][10];				l_cell_reg[577] = inform_L[800][10];				l_cell_reg[578] = inform_L[289][10];				l_cell_reg[579] = inform_L[801][10];				l_cell_reg[580] = inform_L[290][10];				l_cell_reg[581] = inform_L[802][10];				l_cell_reg[582] = inform_L[291][10];				l_cell_reg[583] = inform_L[803][10];				l_cell_reg[584] = inform_L[292][10];				l_cell_reg[585] = inform_L[804][10];				l_cell_reg[586] = inform_L[293][10];				l_cell_reg[587] = inform_L[805][10];				l_cell_reg[588] = inform_L[294][10];				l_cell_reg[589] = inform_L[806][10];				l_cell_reg[590] = inform_L[295][10];				l_cell_reg[591] = inform_L[807][10];				l_cell_reg[592] = inform_L[296][10];				l_cell_reg[593] = inform_L[808][10];				l_cell_reg[594] = inform_L[297][10];				l_cell_reg[595] = inform_L[809][10];				l_cell_reg[596] = inform_L[298][10];				l_cell_reg[597] = inform_L[810][10];				l_cell_reg[598] = inform_L[299][10];				l_cell_reg[599] = inform_L[811][10];				l_cell_reg[600] = inform_L[300][10];				l_cell_reg[601] = inform_L[812][10];				l_cell_reg[602] = inform_L[301][10];				l_cell_reg[603] = inform_L[813][10];				l_cell_reg[604] = inform_L[302][10];				l_cell_reg[605] = inform_L[814][10];				l_cell_reg[606] = inform_L[303][10];				l_cell_reg[607] = inform_L[815][10];				l_cell_reg[608] = inform_L[304][10];				l_cell_reg[609] = inform_L[816][10];				l_cell_reg[610] = inform_L[305][10];				l_cell_reg[611] = inform_L[817][10];				l_cell_reg[612] = inform_L[306][10];				l_cell_reg[613] = inform_L[818][10];				l_cell_reg[614] = inform_L[307][10];				l_cell_reg[615] = inform_L[819][10];				l_cell_reg[616] = inform_L[308][10];				l_cell_reg[617] = inform_L[820][10];				l_cell_reg[618] = inform_L[309][10];				l_cell_reg[619] = inform_L[821][10];				l_cell_reg[620] = inform_L[310][10];				l_cell_reg[621] = inform_L[822][10];				l_cell_reg[622] = inform_L[311][10];				l_cell_reg[623] = inform_L[823][10];				l_cell_reg[624] = inform_L[312][10];				l_cell_reg[625] = inform_L[824][10];				l_cell_reg[626] = inform_L[313][10];				l_cell_reg[627] = inform_L[825][10];				l_cell_reg[628] = inform_L[314][10];				l_cell_reg[629] = inform_L[826][10];				l_cell_reg[630] = inform_L[315][10];				l_cell_reg[631] = inform_L[827][10];				l_cell_reg[632] = inform_L[316][10];				l_cell_reg[633] = inform_L[828][10];				l_cell_reg[634] = inform_L[317][10];				l_cell_reg[635] = inform_L[829][10];				l_cell_reg[636] = inform_L[318][10];				l_cell_reg[637] = inform_L[830][10];				l_cell_reg[638] = inform_L[319][10];				l_cell_reg[639] = inform_L[831][10];				l_cell_reg[640] = inform_L[320][10];				l_cell_reg[641] = inform_L[832][10];				l_cell_reg[642] = inform_L[321][10];				l_cell_reg[643] = inform_L[833][10];				l_cell_reg[644] = inform_L[322][10];				l_cell_reg[645] = inform_L[834][10];				l_cell_reg[646] = inform_L[323][10];				l_cell_reg[647] = inform_L[835][10];				l_cell_reg[648] = inform_L[324][10];				l_cell_reg[649] = inform_L[836][10];				l_cell_reg[650] = inform_L[325][10];				l_cell_reg[651] = inform_L[837][10];				l_cell_reg[652] = inform_L[326][10];				l_cell_reg[653] = inform_L[838][10];				l_cell_reg[654] = inform_L[327][10];				l_cell_reg[655] = inform_L[839][10];				l_cell_reg[656] = inform_L[328][10];				l_cell_reg[657] = inform_L[840][10];				l_cell_reg[658] = inform_L[329][10];				l_cell_reg[659] = inform_L[841][10];				l_cell_reg[660] = inform_L[330][10];				l_cell_reg[661] = inform_L[842][10];				l_cell_reg[662] = inform_L[331][10];				l_cell_reg[663] = inform_L[843][10];				l_cell_reg[664] = inform_L[332][10];				l_cell_reg[665] = inform_L[844][10];				l_cell_reg[666] = inform_L[333][10];				l_cell_reg[667] = inform_L[845][10];				l_cell_reg[668] = inform_L[334][10];				l_cell_reg[669] = inform_L[846][10];				l_cell_reg[670] = inform_L[335][10];				l_cell_reg[671] = inform_L[847][10];				l_cell_reg[672] = inform_L[336][10];				l_cell_reg[673] = inform_L[848][10];				l_cell_reg[674] = inform_L[337][10];				l_cell_reg[675] = inform_L[849][10];				l_cell_reg[676] = inform_L[338][10];				l_cell_reg[677] = inform_L[850][10];				l_cell_reg[678] = inform_L[339][10];				l_cell_reg[679] = inform_L[851][10];				l_cell_reg[680] = inform_L[340][10];				l_cell_reg[681] = inform_L[852][10];				l_cell_reg[682] = inform_L[341][10];				l_cell_reg[683] = inform_L[853][10];				l_cell_reg[684] = inform_L[342][10];				l_cell_reg[685] = inform_L[854][10];				l_cell_reg[686] = inform_L[343][10];				l_cell_reg[687] = inform_L[855][10];				l_cell_reg[688] = inform_L[344][10];				l_cell_reg[689] = inform_L[856][10];				l_cell_reg[690] = inform_L[345][10];				l_cell_reg[691] = inform_L[857][10];				l_cell_reg[692] = inform_L[346][10];				l_cell_reg[693] = inform_L[858][10];				l_cell_reg[694] = inform_L[347][10];				l_cell_reg[695] = inform_L[859][10];				l_cell_reg[696] = inform_L[348][10];				l_cell_reg[697] = inform_L[860][10];				l_cell_reg[698] = inform_L[349][10];				l_cell_reg[699] = inform_L[861][10];				l_cell_reg[700] = inform_L[350][10];				l_cell_reg[701] = inform_L[862][10];				l_cell_reg[702] = inform_L[351][10];				l_cell_reg[703] = inform_L[863][10];				l_cell_reg[704] = inform_L[352][10];				l_cell_reg[705] = inform_L[864][10];				l_cell_reg[706] = inform_L[353][10];				l_cell_reg[707] = inform_L[865][10];				l_cell_reg[708] = inform_L[354][10];				l_cell_reg[709] = inform_L[866][10];				l_cell_reg[710] = inform_L[355][10];				l_cell_reg[711] = inform_L[867][10];				l_cell_reg[712] = inform_L[356][10];				l_cell_reg[713] = inform_L[868][10];				l_cell_reg[714] = inform_L[357][10];				l_cell_reg[715] = inform_L[869][10];				l_cell_reg[716] = inform_L[358][10];				l_cell_reg[717] = inform_L[870][10];				l_cell_reg[718] = inform_L[359][10];				l_cell_reg[719] = inform_L[871][10];				l_cell_reg[720] = inform_L[360][10];				l_cell_reg[721] = inform_L[872][10];				l_cell_reg[722] = inform_L[361][10];				l_cell_reg[723] = inform_L[873][10];				l_cell_reg[724] = inform_L[362][10];				l_cell_reg[725] = inform_L[874][10];				l_cell_reg[726] = inform_L[363][10];				l_cell_reg[727] = inform_L[875][10];				l_cell_reg[728] = inform_L[364][10];				l_cell_reg[729] = inform_L[876][10];				l_cell_reg[730] = inform_L[365][10];				l_cell_reg[731] = inform_L[877][10];				l_cell_reg[732] = inform_L[366][10];				l_cell_reg[733] = inform_L[878][10];				l_cell_reg[734] = inform_L[367][10];				l_cell_reg[735] = inform_L[879][10];				l_cell_reg[736] = inform_L[368][10];				l_cell_reg[737] = inform_L[880][10];				l_cell_reg[738] = inform_L[369][10];				l_cell_reg[739] = inform_L[881][10];				l_cell_reg[740] = inform_L[370][10];				l_cell_reg[741] = inform_L[882][10];				l_cell_reg[742] = inform_L[371][10];				l_cell_reg[743] = inform_L[883][10];				l_cell_reg[744] = inform_L[372][10];				l_cell_reg[745] = inform_L[884][10];				l_cell_reg[746] = inform_L[373][10];				l_cell_reg[747] = inform_L[885][10];				l_cell_reg[748] = inform_L[374][10];				l_cell_reg[749] = inform_L[886][10];				l_cell_reg[750] = inform_L[375][10];				l_cell_reg[751] = inform_L[887][10];				l_cell_reg[752] = inform_L[376][10];				l_cell_reg[753] = inform_L[888][10];				l_cell_reg[754] = inform_L[377][10];				l_cell_reg[755] = inform_L[889][10];				l_cell_reg[756] = inform_L[378][10];				l_cell_reg[757] = inform_L[890][10];				l_cell_reg[758] = inform_L[379][10];				l_cell_reg[759] = inform_L[891][10];				l_cell_reg[760] = inform_L[380][10];				l_cell_reg[761] = inform_L[892][10];				l_cell_reg[762] = inform_L[381][10];				l_cell_reg[763] = inform_L[893][10];				l_cell_reg[764] = inform_L[382][10];				l_cell_reg[765] = inform_L[894][10];				l_cell_reg[766] = inform_L[383][10];				l_cell_reg[767] = inform_L[895][10];				l_cell_reg[768] = inform_L[384][10];				l_cell_reg[769] = inform_L[896][10];				l_cell_reg[770] = inform_L[385][10];				l_cell_reg[771] = inform_L[897][10];				l_cell_reg[772] = inform_L[386][10];				l_cell_reg[773] = inform_L[898][10];				l_cell_reg[774] = inform_L[387][10];				l_cell_reg[775] = inform_L[899][10];				l_cell_reg[776] = inform_L[388][10];				l_cell_reg[777] = inform_L[900][10];				l_cell_reg[778] = inform_L[389][10];				l_cell_reg[779] = inform_L[901][10];				l_cell_reg[780] = inform_L[390][10];				l_cell_reg[781] = inform_L[902][10];				l_cell_reg[782] = inform_L[391][10];				l_cell_reg[783] = inform_L[903][10];				l_cell_reg[784] = inform_L[392][10];				l_cell_reg[785] = inform_L[904][10];				l_cell_reg[786] = inform_L[393][10];				l_cell_reg[787] = inform_L[905][10];				l_cell_reg[788] = inform_L[394][10];				l_cell_reg[789] = inform_L[906][10];				l_cell_reg[790] = inform_L[395][10];				l_cell_reg[791] = inform_L[907][10];				l_cell_reg[792] = inform_L[396][10];				l_cell_reg[793] = inform_L[908][10];				l_cell_reg[794] = inform_L[397][10];				l_cell_reg[795] = inform_L[909][10];				l_cell_reg[796] = inform_L[398][10];				l_cell_reg[797] = inform_L[910][10];				l_cell_reg[798] = inform_L[399][10];				l_cell_reg[799] = inform_L[911][10];				l_cell_reg[800] = inform_L[400][10];				l_cell_reg[801] = inform_L[912][10];				l_cell_reg[802] = inform_L[401][10];				l_cell_reg[803] = inform_L[913][10];				l_cell_reg[804] = inform_L[402][10];				l_cell_reg[805] = inform_L[914][10];				l_cell_reg[806] = inform_L[403][10];				l_cell_reg[807] = inform_L[915][10];				l_cell_reg[808] = inform_L[404][10];				l_cell_reg[809] = inform_L[916][10];				l_cell_reg[810] = inform_L[405][10];				l_cell_reg[811] = inform_L[917][10];				l_cell_reg[812] = inform_L[406][10];				l_cell_reg[813] = inform_L[918][10];				l_cell_reg[814] = inform_L[407][10];				l_cell_reg[815] = inform_L[919][10];				l_cell_reg[816] = inform_L[408][10];				l_cell_reg[817] = inform_L[920][10];				l_cell_reg[818] = inform_L[409][10];				l_cell_reg[819] = inform_L[921][10];				l_cell_reg[820] = inform_L[410][10];				l_cell_reg[821] = inform_L[922][10];				l_cell_reg[822] = inform_L[411][10];				l_cell_reg[823] = inform_L[923][10];				l_cell_reg[824] = inform_L[412][10];				l_cell_reg[825] = inform_L[924][10];				l_cell_reg[826] = inform_L[413][10];				l_cell_reg[827] = inform_L[925][10];				l_cell_reg[828] = inform_L[414][10];				l_cell_reg[829] = inform_L[926][10];				l_cell_reg[830] = inform_L[415][10];				l_cell_reg[831] = inform_L[927][10];				l_cell_reg[832] = inform_L[416][10];				l_cell_reg[833] = inform_L[928][10];				l_cell_reg[834] = inform_L[417][10];				l_cell_reg[835] = inform_L[929][10];				l_cell_reg[836] = inform_L[418][10];				l_cell_reg[837] = inform_L[930][10];				l_cell_reg[838] = inform_L[419][10];				l_cell_reg[839] = inform_L[931][10];				l_cell_reg[840] = inform_L[420][10];				l_cell_reg[841] = inform_L[932][10];				l_cell_reg[842] = inform_L[421][10];				l_cell_reg[843] = inform_L[933][10];				l_cell_reg[844] = inform_L[422][10];				l_cell_reg[845] = inform_L[934][10];				l_cell_reg[846] = inform_L[423][10];				l_cell_reg[847] = inform_L[935][10];				l_cell_reg[848] = inform_L[424][10];				l_cell_reg[849] = inform_L[936][10];				l_cell_reg[850] = inform_L[425][10];				l_cell_reg[851] = inform_L[937][10];				l_cell_reg[852] = inform_L[426][10];				l_cell_reg[853] = inform_L[938][10];				l_cell_reg[854] = inform_L[427][10];				l_cell_reg[855] = inform_L[939][10];				l_cell_reg[856] = inform_L[428][10];				l_cell_reg[857] = inform_L[940][10];				l_cell_reg[858] = inform_L[429][10];				l_cell_reg[859] = inform_L[941][10];				l_cell_reg[860] = inform_L[430][10];				l_cell_reg[861] = inform_L[942][10];				l_cell_reg[862] = inform_L[431][10];				l_cell_reg[863] = inform_L[943][10];				l_cell_reg[864] = inform_L[432][10];				l_cell_reg[865] = inform_L[944][10];				l_cell_reg[866] = inform_L[433][10];				l_cell_reg[867] = inform_L[945][10];				l_cell_reg[868] = inform_L[434][10];				l_cell_reg[869] = inform_L[946][10];				l_cell_reg[870] = inform_L[435][10];				l_cell_reg[871] = inform_L[947][10];				l_cell_reg[872] = inform_L[436][10];				l_cell_reg[873] = inform_L[948][10];				l_cell_reg[874] = inform_L[437][10];				l_cell_reg[875] = inform_L[949][10];				l_cell_reg[876] = inform_L[438][10];				l_cell_reg[877] = inform_L[950][10];				l_cell_reg[878] = inform_L[439][10];				l_cell_reg[879] = inform_L[951][10];				l_cell_reg[880] = inform_L[440][10];				l_cell_reg[881] = inform_L[952][10];				l_cell_reg[882] = inform_L[441][10];				l_cell_reg[883] = inform_L[953][10];				l_cell_reg[884] = inform_L[442][10];				l_cell_reg[885] = inform_L[954][10];				l_cell_reg[886] = inform_L[443][10];				l_cell_reg[887] = inform_L[955][10];				l_cell_reg[888] = inform_L[444][10];				l_cell_reg[889] = inform_L[956][10];				l_cell_reg[890] = inform_L[445][10];				l_cell_reg[891] = inform_L[957][10];				l_cell_reg[892] = inform_L[446][10];				l_cell_reg[893] = inform_L[958][10];				l_cell_reg[894] = inform_L[447][10];				l_cell_reg[895] = inform_L[959][10];				l_cell_reg[896] = inform_L[448][10];				l_cell_reg[897] = inform_L[960][10];				l_cell_reg[898] = inform_L[449][10];				l_cell_reg[899] = inform_L[961][10];				l_cell_reg[900] = inform_L[450][10];				l_cell_reg[901] = inform_L[962][10];				l_cell_reg[902] = inform_L[451][10];				l_cell_reg[903] = inform_L[963][10];				l_cell_reg[904] = inform_L[452][10];				l_cell_reg[905] = inform_L[964][10];				l_cell_reg[906] = inform_L[453][10];				l_cell_reg[907] = inform_L[965][10];				l_cell_reg[908] = inform_L[454][10];				l_cell_reg[909] = inform_L[966][10];				l_cell_reg[910] = inform_L[455][10];				l_cell_reg[911] = inform_L[967][10];				l_cell_reg[912] = inform_L[456][10];				l_cell_reg[913] = inform_L[968][10];				l_cell_reg[914] = inform_L[457][10];				l_cell_reg[915] = inform_L[969][10];				l_cell_reg[916] = inform_L[458][10];				l_cell_reg[917] = inform_L[970][10];				l_cell_reg[918] = inform_L[459][10];				l_cell_reg[919] = inform_L[971][10];				l_cell_reg[920] = inform_L[460][10];				l_cell_reg[921] = inform_L[972][10];				l_cell_reg[922] = inform_L[461][10];				l_cell_reg[923] = inform_L[973][10];				l_cell_reg[924] = inform_L[462][10];				l_cell_reg[925] = inform_L[974][10];				l_cell_reg[926] = inform_L[463][10];				l_cell_reg[927] = inform_L[975][10];				l_cell_reg[928] = inform_L[464][10];				l_cell_reg[929] = inform_L[976][10];				l_cell_reg[930] = inform_L[465][10];				l_cell_reg[931] = inform_L[977][10];				l_cell_reg[932] = inform_L[466][10];				l_cell_reg[933] = inform_L[978][10];				l_cell_reg[934] = inform_L[467][10];				l_cell_reg[935] = inform_L[979][10];				l_cell_reg[936] = inform_L[468][10];				l_cell_reg[937] = inform_L[980][10];				l_cell_reg[938] = inform_L[469][10];				l_cell_reg[939] = inform_L[981][10];				l_cell_reg[940] = inform_L[470][10];				l_cell_reg[941] = inform_L[982][10];				l_cell_reg[942] = inform_L[471][10];				l_cell_reg[943] = inform_L[983][10];				l_cell_reg[944] = inform_L[472][10];				l_cell_reg[945] = inform_L[984][10];				l_cell_reg[946] = inform_L[473][10];				l_cell_reg[947] = inform_L[985][10];				l_cell_reg[948] = inform_L[474][10];				l_cell_reg[949] = inform_L[986][10];				l_cell_reg[950] = inform_L[475][10];				l_cell_reg[951] = inform_L[987][10];				l_cell_reg[952] = inform_L[476][10];				l_cell_reg[953] = inform_L[988][10];				l_cell_reg[954] = inform_L[477][10];				l_cell_reg[955] = inform_L[989][10];				l_cell_reg[956] = inform_L[478][10];				l_cell_reg[957] = inform_L[990][10];				l_cell_reg[958] = inform_L[479][10];				l_cell_reg[959] = inform_L[991][10];				l_cell_reg[960] = inform_L[480][10];				l_cell_reg[961] = inform_L[992][10];				l_cell_reg[962] = inform_L[481][10];				l_cell_reg[963] = inform_L[993][10];				l_cell_reg[964] = inform_L[482][10];				l_cell_reg[965] = inform_L[994][10];				l_cell_reg[966] = inform_L[483][10];				l_cell_reg[967] = inform_L[995][10];				l_cell_reg[968] = inform_L[484][10];				l_cell_reg[969] = inform_L[996][10];				l_cell_reg[970] = inform_L[485][10];				l_cell_reg[971] = inform_L[997][10];				l_cell_reg[972] = inform_L[486][10];				l_cell_reg[973] = inform_L[998][10];				l_cell_reg[974] = inform_L[487][10];				l_cell_reg[975] = inform_L[999][10];				l_cell_reg[976] = inform_L[488][10];				l_cell_reg[977] = inform_L[1000][10];				l_cell_reg[978] = inform_L[489][10];				l_cell_reg[979] = inform_L[1001][10];				l_cell_reg[980] = inform_L[490][10];				l_cell_reg[981] = inform_L[1002][10];				l_cell_reg[982] = inform_L[491][10];				l_cell_reg[983] = inform_L[1003][10];				l_cell_reg[984] = inform_L[492][10];				l_cell_reg[985] = inform_L[1004][10];				l_cell_reg[986] = inform_L[493][10];				l_cell_reg[987] = inform_L[1005][10];				l_cell_reg[988] = inform_L[494][10];				l_cell_reg[989] = inform_L[1006][10];				l_cell_reg[990] = inform_L[495][10];				l_cell_reg[991] = inform_L[1007][10];				l_cell_reg[992] = inform_L[496][10];				l_cell_reg[993] = inform_L[1008][10];				l_cell_reg[994] = inform_L[497][10];				l_cell_reg[995] = inform_L[1009][10];				l_cell_reg[996] = inform_L[498][10];				l_cell_reg[997] = inform_L[1010][10];				l_cell_reg[998] = inform_L[499][10];				l_cell_reg[999] = inform_L[1011][10];				l_cell_reg[1000] = inform_L[500][10];				l_cell_reg[1001] = inform_L[1012][10];				l_cell_reg[1002] = inform_L[501][10];				l_cell_reg[1003] = inform_L[1013][10];				l_cell_reg[1004] = inform_L[502][10];				l_cell_reg[1005] = inform_L[1014][10];				l_cell_reg[1006] = inform_L[503][10];				l_cell_reg[1007] = inform_L[1015][10];				l_cell_reg[1008] = inform_L[504][10];				l_cell_reg[1009] = inform_L[1016][10];				l_cell_reg[1010] = inform_L[505][10];				l_cell_reg[1011] = inform_L[1017][10];				l_cell_reg[1012] = inform_L[506][10];				l_cell_reg[1013] = inform_L[1018][10];				l_cell_reg[1014] = inform_L[507][10];				l_cell_reg[1015] = inform_L[1019][10];				l_cell_reg[1016] = inform_L[508][10];				l_cell_reg[1017] = inform_L[1020][10];				l_cell_reg[1018] = inform_L[509][10];				l_cell_reg[1019] = inform_L[1021][10];				l_cell_reg[1020] = inform_L[510][10];				l_cell_reg[1021] = inform_L[1022][10];				l_cell_reg[1022] = inform_L[511][10];				l_cell_reg[1023] = inform_L[1023][10];			end
			default:			begin					r_cell_reg[0] <= 0;					r_cell_reg[1] <= 0;					r_cell_reg[2] <= 0;					r_cell_reg[3] <= 0;					r_cell_reg[4] <= 0;					r_cell_reg[5] <= 0;					r_cell_reg[6] <= 0;					r_cell_reg[7] <= 0;					r_cell_reg[8] <= 0;					r_cell_reg[9] <= 0;					r_cell_reg[10] <= 0;					r_cell_reg[11] <= 0;					r_cell_reg[12] <= 0;					r_cell_reg[13] <= 0;					r_cell_reg[14] <= 0;					r_cell_reg[15] <= 0;					r_cell_reg[16] <= 0;					r_cell_reg[17] <= 0;					r_cell_reg[18] <= 0;					r_cell_reg[19] <= 0;					r_cell_reg[20] <= 0;					r_cell_reg[21] <= 0;					r_cell_reg[22] <= 0;					r_cell_reg[23] <= 0;					r_cell_reg[24] <= 0;					r_cell_reg[25] <= 0;					r_cell_reg[26] <= 0;					r_cell_reg[27] <= 0;					r_cell_reg[28] <= 0;					r_cell_reg[29] <= 0;					r_cell_reg[30] <= 0;					r_cell_reg[31] <= 0;					r_cell_reg[32] <= 0;					r_cell_reg[33] <= 0;					r_cell_reg[34] <= 0;					r_cell_reg[35] <= 0;					r_cell_reg[36] <= 0;					r_cell_reg[37] <= 0;					r_cell_reg[38] <= 0;					r_cell_reg[39] <= 0;					r_cell_reg[40] <= 0;					r_cell_reg[41] <= 0;					r_cell_reg[42] <= 0;					r_cell_reg[43] <= 0;					r_cell_reg[44] <= 0;					r_cell_reg[45] <= 0;					r_cell_reg[46] <= 0;					r_cell_reg[47] <= 0;					r_cell_reg[48] <= 0;					r_cell_reg[49] <= 0;					r_cell_reg[50] <= 0;					r_cell_reg[51] <= 0;					r_cell_reg[52] <= 0;					r_cell_reg[53] <= 0;					r_cell_reg[54] <= 0;					r_cell_reg[55] <= 0;					r_cell_reg[56] <= 0;					r_cell_reg[57] <= 0;					r_cell_reg[58] <= 0;					r_cell_reg[59] <= 0;					r_cell_reg[60] <= 0;					r_cell_reg[61] <= 0;					r_cell_reg[62] <= 0;					r_cell_reg[63] <= 0;					r_cell_reg[64] <= 0;					r_cell_reg[65] <= 0;					r_cell_reg[66] <= 0;					r_cell_reg[67] <= 0;					r_cell_reg[68] <= 0;					r_cell_reg[69] <= 0;					r_cell_reg[70] <= 0;					r_cell_reg[71] <= 0;					r_cell_reg[72] <= 0;					r_cell_reg[73] <= 0;					r_cell_reg[74] <= 0;					r_cell_reg[75] <= 0;					r_cell_reg[76] <= 0;					r_cell_reg[77] <= 0;					r_cell_reg[78] <= 0;					r_cell_reg[79] <= 0;					r_cell_reg[80] <= 0;					r_cell_reg[81] <= 0;					r_cell_reg[82] <= 0;					r_cell_reg[83] <= 0;					r_cell_reg[84] <= 0;					r_cell_reg[85] <= 0;					r_cell_reg[86] <= 0;					r_cell_reg[87] <= 0;					r_cell_reg[88] <= 0;					r_cell_reg[89] <= 0;					r_cell_reg[90] <= 0;					r_cell_reg[91] <= 0;					r_cell_reg[92] <= 0;					r_cell_reg[93] <= 0;					r_cell_reg[94] <= 0;					r_cell_reg[95] <= 0;					r_cell_reg[96] <= 0;					r_cell_reg[97] <= 0;					r_cell_reg[98] <= 0;					r_cell_reg[99] <= 0;					r_cell_reg[100] <= 0;					r_cell_reg[101] <= 0;					r_cell_reg[102] <= 0;					r_cell_reg[103] <= 0;					r_cell_reg[104] <= 0;					r_cell_reg[105] <= 0;					r_cell_reg[106] <= 0;					r_cell_reg[107] <= 0;					r_cell_reg[108] <= 0;					r_cell_reg[109] <= 0;					r_cell_reg[110] <= 0;					r_cell_reg[111] <= 0;					r_cell_reg[112] <= 0;					r_cell_reg[113] <= 0;					r_cell_reg[114] <= 0;					r_cell_reg[115] <= 0;					r_cell_reg[116] <= 0;					r_cell_reg[117] <= 0;					r_cell_reg[118] <= 0;					r_cell_reg[119] <= 0;					r_cell_reg[120] <= 0;					r_cell_reg[121] <= 0;					r_cell_reg[122] <= 0;					r_cell_reg[123] <= 0;					r_cell_reg[124] <= 0;					r_cell_reg[125] <= 0;					r_cell_reg[126] <= 0;					r_cell_reg[127] <= 0;					r_cell_reg[128] <= 0;					r_cell_reg[129] <= 0;					r_cell_reg[130] <= 0;					r_cell_reg[131] <= 0;					r_cell_reg[132] <= 0;					r_cell_reg[133] <= 0;					r_cell_reg[134] <= 0;					r_cell_reg[135] <= 0;					r_cell_reg[136] <= 0;					r_cell_reg[137] <= 0;					r_cell_reg[138] <= 0;					r_cell_reg[139] <= 0;					r_cell_reg[140] <= 0;					r_cell_reg[141] <= 0;					r_cell_reg[142] <= 0;					r_cell_reg[143] <= 0;					r_cell_reg[144] <= 0;					r_cell_reg[145] <= 0;					r_cell_reg[146] <= 0;					r_cell_reg[147] <= 0;					r_cell_reg[148] <= 0;					r_cell_reg[149] <= 0;					r_cell_reg[150] <= 0;					r_cell_reg[151] <= 0;					r_cell_reg[152] <= 0;					r_cell_reg[153] <= 0;					r_cell_reg[154] <= 0;					r_cell_reg[155] <= 0;					r_cell_reg[156] <= 0;					r_cell_reg[157] <= 0;					r_cell_reg[158] <= 0;					r_cell_reg[159] <= 0;					r_cell_reg[160] <= 0;					r_cell_reg[161] <= 0;					r_cell_reg[162] <= 0;					r_cell_reg[163] <= 0;					r_cell_reg[164] <= 0;					r_cell_reg[165] <= 0;					r_cell_reg[166] <= 0;					r_cell_reg[167] <= 0;					r_cell_reg[168] <= 0;					r_cell_reg[169] <= 0;					r_cell_reg[170] <= 0;					r_cell_reg[171] <= 0;					r_cell_reg[172] <= 0;					r_cell_reg[173] <= 0;					r_cell_reg[174] <= 0;					r_cell_reg[175] <= 0;					r_cell_reg[176] <= 0;					r_cell_reg[177] <= 0;					r_cell_reg[178] <= 0;					r_cell_reg[179] <= 0;					r_cell_reg[180] <= 0;					r_cell_reg[181] <= 0;					r_cell_reg[182] <= 0;					r_cell_reg[183] <= 0;					r_cell_reg[184] <= 0;					r_cell_reg[185] <= 0;					r_cell_reg[186] <= 0;					r_cell_reg[187] <= 0;					r_cell_reg[188] <= 0;					r_cell_reg[189] <= 0;					r_cell_reg[190] <= 0;					r_cell_reg[191] <= 0;					r_cell_reg[192] <= 0;					r_cell_reg[193] <= 0;					r_cell_reg[194] <= 0;					r_cell_reg[195] <= 0;					r_cell_reg[196] <= 0;					r_cell_reg[197] <= 0;					r_cell_reg[198] <= 0;					r_cell_reg[199] <= 0;					r_cell_reg[200] <= 0;					r_cell_reg[201] <= 0;					r_cell_reg[202] <= 0;					r_cell_reg[203] <= 0;					r_cell_reg[204] <= 0;					r_cell_reg[205] <= 0;					r_cell_reg[206] <= 0;					r_cell_reg[207] <= 0;					r_cell_reg[208] <= 0;					r_cell_reg[209] <= 0;					r_cell_reg[210] <= 0;					r_cell_reg[211] <= 0;					r_cell_reg[212] <= 0;					r_cell_reg[213] <= 0;					r_cell_reg[214] <= 0;					r_cell_reg[215] <= 0;					r_cell_reg[216] <= 0;					r_cell_reg[217] <= 0;					r_cell_reg[218] <= 0;					r_cell_reg[219] <= 0;					r_cell_reg[220] <= 0;					r_cell_reg[221] <= 0;					r_cell_reg[222] <= 0;					r_cell_reg[223] <= 0;					r_cell_reg[224] <= 0;					r_cell_reg[225] <= 0;					r_cell_reg[226] <= 0;					r_cell_reg[227] <= 0;					r_cell_reg[228] <= 0;					r_cell_reg[229] <= 0;					r_cell_reg[230] <= 0;					r_cell_reg[231] <= 0;					r_cell_reg[232] <= 0;					r_cell_reg[233] <= 0;					r_cell_reg[234] <= 0;					r_cell_reg[235] <= 0;					r_cell_reg[236] <= 0;					r_cell_reg[237] <= 0;					r_cell_reg[238] <= 0;					r_cell_reg[239] <= 0;					r_cell_reg[240] <= 0;					r_cell_reg[241] <= 0;					r_cell_reg[242] <= 0;					r_cell_reg[243] <= 0;					r_cell_reg[244] <= 0;					r_cell_reg[245] <= 0;					r_cell_reg[246] <= 0;					r_cell_reg[247] <= 0;					r_cell_reg[248] <= 0;					r_cell_reg[249] <= 0;					r_cell_reg[250] <= 0;					r_cell_reg[251] <= 0;					r_cell_reg[252] <= 0;					r_cell_reg[253] <= 0;					r_cell_reg[254] <= 0;					r_cell_reg[255] <= 0;					r_cell_reg[256] <= 0;					r_cell_reg[257] <= 0;					r_cell_reg[258] <= 0;					r_cell_reg[259] <= 0;					r_cell_reg[260] <= 0;					r_cell_reg[261] <= 0;					r_cell_reg[262] <= 0;					r_cell_reg[263] <= 0;					r_cell_reg[264] <= 0;					r_cell_reg[265] <= 0;					r_cell_reg[266] <= 0;					r_cell_reg[267] <= 0;					r_cell_reg[268] <= 0;					r_cell_reg[269] <= 0;					r_cell_reg[270] <= 0;					r_cell_reg[271] <= 0;					r_cell_reg[272] <= 0;					r_cell_reg[273] <= 0;					r_cell_reg[274] <= 0;					r_cell_reg[275] <= 0;					r_cell_reg[276] <= 0;					r_cell_reg[277] <= 0;					r_cell_reg[278] <= 0;					r_cell_reg[279] <= 0;					r_cell_reg[280] <= 0;					r_cell_reg[281] <= 0;					r_cell_reg[282] <= 0;					r_cell_reg[283] <= 0;					r_cell_reg[284] <= 0;					r_cell_reg[285] <= 0;					r_cell_reg[286] <= 0;					r_cell_reg[287] <= 0;					r_cell_reg[288] <= 0;					r_cell_reg[289] <= 0;					r_cell_reg[290] <= 0;					r_cell_reg[291] <= 0;					r_cell_reg[292] <= 0;					r_cell_reg[293] <= 0;					r_cell_reg[294] <= 0;					r_cell_reg[295] <= 0;					r_cell_reg[296] <= 0;					r_cell_reg[297] <= 0;					r_cell_reg[298] <= 0;					r_cell_reg[299] <= 0;					r_cell_reg[300] <= 0;					r_cell_reg[301] <= 0;					r_cell_reg[302] <= 0;					r_cell_reg[303] <= 0;					r_cell_reg[304] <= 0;					r_cell_reg[305] <= 0;					r_cell_reg[306] <= 0;					r_cell_reg[307] <= 0;					r_cell_reg[308] <= 0;					r_cell_reg[309] <= 0;					r_cell_reg[310] <= 0;					r_cell_reg[311] <= 0;					r_cell_reg[312] <= 0;					r_cell_reg[313] <= 0;					r_cell_reg[314] <= 0;					r_cell_reg[315] <= 0;					r_cell_reg[316] <= 0;					r_cell_reg[317] <= 0;					r_cell_reg[318] <= 0;					r_cell_reg[319] <= 0;					r_cell_reg[320] <= 0;					r_cell_reg[321] <= 0;					r_cell_reg[322] <= 0;					r_cell_reg[323] <= 0;					r_cell_reg[324] <= 0;					r_cell_reg[325] <= 0;					r_cell_reg[326] <= 0;					r_cell_reg[327] <= 0;					r_cell_reg[328] <= 0;					r_cell_reg[329] <= 0;					r_cell_reg[330] <= 0;					r_cell_reg[331] <= 0;					r_cell_reg[332] <= 0;					r_cell_reg[333] <= 0;					r_cell_reg[334] <= 0;					r_cell_reg[335] <= 0;					r_cell_reg[336] <= 0;					r_cell_reg[337] <= 0;					r_cell_reg[338] <= 0;					r_cell_reg[339] <= 0;					r_cell_reg[340] <= 0;					r_cell_reg[341] <= 0;					r_cell_reg[342] <= 0;					r_cell_reg[343] <= 0;					r_cell_reg[344] <= 0;					r_cell_reg[345] <= 0;					r_cell_reg[346] <= 0;					r_cell_reg[347] <= 0;					r_cell_reg[348] <= 0;					r_cell_reg[349] <= 0;					r_cell_reg[350] <= 0;					r_cell_reg[351] <= 0;					r_cell_reg[352] <= 0;					r_cell_reg[353] <= 0;					r_cell_reg[354] <= 0;					r_cell_reg[355] <= 0;					r_cell_reg[356] <= 0;					r_cell_reg[357] <= 0;					r_cell_reg[358] <= 0;					r_cell_reg[359] <= 0;					r_cell_reg[360] <= 0;					r_cell_reg[361] <= 0;					r_cell_reg[362] <= 0;					r_cell_reg[363] <= 0;					r_cell_reg[364] <= 0;					r_cell_reg[365] <= 0;					r_cell_reg[366] <= 0;					r_cell_reg[367] <= 0;					r_cell_reg[368] <= 0;					r_cell_reg[369] <= 0;					r_cell_reg[370] <= 0;					r_cell_reg[371] <= 0;					r_cell_reg[372] <= 0;					r_cell_reg[373] <= 0;					r_cell_reg[374] <= 0;					r_cell_reg[375] <= 0;					r_cell_reg[376] <= 0;					r_cell_reg[377] <= 0;					r_cell_reg[378] <= 0;					r_cell_reg[379] <= 0;					r_cell_reg[380] <= 0;					r_cell_reg[381] <= 0;					r_cell_reg[382] <= 0;					r_cell_reg[383] <= 0;					r_cell_reg[384] <= 0;					r_cell_reg[385] <= 0;					r_cell_reg[386] <= 0;					r_cell_reg[387] <= 0;					r_cell_reg[388] <= 0;					r_cell_reg[389] <= 0;					r_cell_reg[390] <= 0;					r_cell_reg[391] <= 0;					r_cell_reg[392] <= 0;					r_cell_reg[393] <= 0;					r_cell_reg[394] <= 0;					r_cell_reg[395] <= 0;					r_cell_reg[396] <= 0;					r_cell_reg[397] <= 0;					r_cell_reg[398] <= 0;					r_cell_reg[399] <= 0;					r_cell_reg[400] <= 0;					r_cell_reg[401] <= 0;					r_cell_reg[402] <= 0;					r_cell_reg[403] <= 0;					r_cell_reg[404] <= 0;					r_cell_reg[405] <= 0;					r_cell_reg[406] <= 0;					r_cell_reg[407] <= 0;					r_cell_reg[408] <= 0;					r_cell_reg[409] <= 0;					r_cell_reg[410] <= 0;					r_cell_reg[411] <= 0;					r_cell_reg[412] <= 0;					r_cell_reg[413] <= 0;					r_cell_reg[414] <= 0;					r_cell_reg[415] <= 0;					r_cell_reg[416] <= 0;					r_cell_reg[417] <= 0;					r_cell_reg[418] <= 0;					r_cell_reg[419] <= 0;					r_cell_reg[420] <= 0;					r_cell_reg[421] <= 0;					r_cell_reg[422] <= 0;					r_cell_reg[423] <= 0;					r_cell_reg[424] <= 0;					r_cell_reg[425] <= 0;					r_cell_reg[426] <= 0;					r_cell_reg[427] <= 0;					r_cell_reg[428] <= 0;					r_cell_reg[429] <= 0;					r_cell_reg[430] <= 0;					r_cell_reg[431] <= 0;					r_cell_reg[432] <= 0;					r_cell_reg[433] <= 0;					r_cell_reg[434] <= 0;					r_cell_reg[435] <= 0;					r_cell_reg[436] <= 0;					r_cell_reg[437] <= 0;					r_cell_reg[438] <= 0;					r_cell_reg[439] <= 0;					r_cell_reg[440] <= 0;					r_cell_reg[441] <= 0;					r_cell_reg[442] <= 0;					r_cell_reg[443] <= 0;					r_cell_reg[444] <= 0;					r_cell_reg[445] <= 0;					r_cell_reg[446] <= 0;					r_cell_reg[447] <= 0;					r_cell_reg[448] <= 0;					r_cell_reg[449] <= 0;					r_cell_reg[450] <= 0;					r_cell_reg[451] <= 0;					r_cell_reg[452] <= 0;					r_cell_reg[453] <= 0;					r_cell_reg[454] <= 0;					r_cell_reg[455] <= 0;					r_cell_reg[456] <= 0;					r_cell_reg[457] <= 0;					r_cell_reg[458] <= 0;					r_cell_reg[459] <= 0;					r_cell_reg[460] <= 0;					r_cell_reg[461] <= 0;					r_cell_reg[462] <= 0;					r_cell_reg[463] <= 0;					r_cell_reg[464] <= 0;					r_cell_reg[465] <= 0;					r_cell_reg[466] <= 0;					r_cell_reg[467] <= 0;					r_cell_reg[468] <= 0;					r_cell_reg[469] <= 0;					r_cell_reg[470] <= 0;					r_cell_reg[471] <= 0;					r_cell_reg[472] <= 0;					r_cell_reg[473] <= 0;					r_cell_reg[474] <= 0;					r_cell_reg[475] <= 0;					r_cell_reg[476] <= 0;					r_cell_reg[477] <= 0;					r_cell_reg[478] <= 0;					r_cell_reg[479] <= 0;					r_cell_reg[480] <= 0;					r_cell_reg[481] <= 0;					r_cell_reg[482] <= 0;					r_cell_reg[483] <= 0;					r_cell_reg[484] <= 0;					r_cell_reg[485] <= 0;					r_cell_reg[486] <= 0;					r_cell_reg[487] <= 0;					r_cell_reg[488] <= 0;					r_cell_reg[489] <= 0;					r_cell_reg[490] <= 0;					r_cell_reg[491] <= 0;					r_cell_reg[492] <= 0;					r_cell_reg[493] <= 0;					r_cell_reg[494] <= 0;					r_cell_reg[495] <= 0;					r_cell_reg[496] <= 0;					r_cell_reg[497] <= 0;					r_cell_reg[498] <= 0;					r_cell_reg[499] <= 0;					r_cell_reg[500] <= 0;					r_cell_reg[501] <= 0;					r_cell_reg[502] <= 0;					r_cell_reg[503] <= 0;					r_cell_reg[504] <= 0;					r_cell_reg[505] <= 0;					r_cell_reg[506] <= 0;					r_cell_reg[507] <= 0;					r_cell_reg[508] <= 0;					r_cell_reg[509] <= 0;					r_cell_reg[510] <= 0;					r_cell_reg[511] <= 0;					r_cell_reg[512] <= 0;					r_cell_reg[513] <= 0;					r_cell_reg[514] <= 0;					r_cell_reg[515] <= 0;					r_cell_reg[516] <= 0;					r_cell_reg[517] <= 0;					r_cell_reg[518] <= 0;					r_cell_reg[519] <= 0;					r_cell_reg[520] <= 0;					r_cell_reg[521] <= 0;					r_cell_reg[522] <= 0;					r_cell_reg[523] <= 0;					r_cell_reg[524] <= 0;					r_cell_reg[525] <= 0;					r_cell_reg[526] <= 0;					r_cell_reg[527] <= 0;					r_cell_reg[528] <= 0;					r_cell_reg[529] <= 0;					r_cell_reg[530] <= 0;					r_cell_reg[531] <= 0;					r_cell_reg[532] <= 0;					r_cell_reg[533] <= 0;					r_cell_reg[534] <= 0;					r_cell_reg[535] <= 0;					r_cell_reg[536] <= 0;					r_cell_reg[537] <= 0;					r_cell_reg[538] <= 0;					r_cell_reg[539] <= 0;					r_cell_reg[540] <= 0;					r_cell_reg[541] <= 0;					r_cell_reg[542] <= 0;					r_cell_reg[543] <= 0;					r_cell_reg[544] <= 0;					r_cell_reg[545] <= 0;					r_cell_reg[546] <= 0;					r_cell_reg[547] <= 0;					r_cell_reg[548] <= 0;					r_cell_reg[549] <= 0;					r_cell_reg[550] <= 0;					r_cell_reg[551] <= 0;					r_cell_reg[552] <= 0;					r_cell_reg[553] <= 0;					r_cell_reg[554] <= 0;					r_cell_reg[555] <= 0;					r_cell_reg[556] <= 0;					r_cell_reg[557] <= 0;					r_cell_reg[558] <= 0;					r_cell_reg[559] <= 0;					r_cell_reg[560] <= 0;					r_cell_reg[561] <= 0;					r_cell_reg[562] <= 0;					r_cell_reg[563] <= 0;					r_cell_reg[564] <= 0;					r_cell_reg[565] <= 0;					r_cell_reg[566] <= 0;					r_cell_reg[567] <= 0;					r_cell_reg[568] <= 0;					r_cell_reg[569] <= 0;					r_cell_reg[570] <= 0;					r_cell_reg[571] <= 0;					r_cell_reg[572] <= 0;					r_cell_reg[573] <= 0;					r_cell_reg[574] <= 0;					r_cell_reg[575] <= 0;					r_cell_reg[576] <= 0;					r_cell_reg[577] <= 0;					r_cell_reg[578] <= 0;					r_cell_reg[579] <= 0;					r_cell_reg[580] <= 0;					r_cell_reg[581] <= 0;					r_cell_reg[582] <= 0;					r_cell_reg[583] <= 0;					r_cell_reg[584] <= 0;					r_cell_reg[585] <= 0;					r_cell_reg[586] <= 0;					r_cell_reg[587] <= 0;					r_cell_reg[588] <= 0;					r_cell_reg[589] <= 0;					r_cell_reg[590] <= 0;					r_cell_reg[591] <= 0;					r_cell_reg[592] <= 0;					r_cell_reg[593] <= 0;					r_cell_reg[594] <= 0;					r_cell_reg[595] <= 0;					r_cell_reg[596] <= 0;					r_cell_reg[597] <= 0;					r_cell_reg[598] <= 0;					r_cell_reg[599] <= 0;					r_cell_reg[600] <= 0;					r_cell_reg[601] <= 0;					r_cell_reg[602] <= 0;					r_cell_reg[603] <= 0;					r_cell_reg[604] <= 0;					r_cell_reg[605] <= 0;					r_cell_reg[606] <= 0;					r_cell_reg[607] <= 0;					r_cell_reg[608] <= 0;					r_cell_reg[609] <= 0;					r_cell_reg[610] <= 0;					r_cell_reg[611] <= 0;					r_cell_reg[612] <= 0;					r_cell_reg[613] <= 0;					r_cell_reg[614] <= 0;					r_cell_reg[615] <= 0;					r_cell_reg[616] <= 0;					r_cell_reg[617] <= 0;					r_cell_reg[618] <= 0;					r_cell_reg[619] <= 0;					r_cell_reg[620] <= 0;					r_cell_reg[621] <= 0;					r_cell_reg[622] <= 0;					r_cell_reg[623] <= 0;					r_cell_reg[624] <= 0;					r_cell_reg[625] <= 0;					r_cell_reg[626] <= 0;					r_cell_reg[627] <= 0;					r_cell_reg[628] <= 0;					r_cell_reg[629] <= 0;					r_cell_reg[630] <= 0;					r_cell_reg[631] <= 0;					r_cell_reg[632] <= 0;					r_cell_reg[633] <= 0;					r_cell_reg[634] <= 0;					r_cell_reg[635] <= 0;					r_cell_reg[636] <= 0;					r_cell_reg[637] <= 0;					r_cell_reg[638] <= 0;					r_cell_reg[639] <= 0;					r_cell_reg[640] <= 0;					r_cell_reg[641] <= 0;					r_cell_reg[642] <= 0;					r_cell_reg[643] <= 0;					r_cell_reg[644] <= 0;					r_cell_reg[645] <= 0;					r_cell_reg[646] <= 0;					r_cell_reg[647] <= 0;					r_cell_reg[648] <= 0;					r_cell_reg[649] <= 0;					r_cell_reg[650] <= 0;					r_cell_reg[651] <= 0;					r_cell_reg[652] <= 0;					r_cell_reg[653] <= 0;					r_cell_reg[654] <= 0;					r_cell_reg[655] <= 0;					r_cell_reg[656] <= 0;					r_cell_reg[657] <= 0;					r_cell_reg[658] <= 0;					r_cell_reg[659] <= 0;					r_cell_reg[660] <= 0;					r_cell_reg[661] <= 0;					r_cell_reg[662] <= 0;					r_cell_reg[663] <= 0;					r_cell_reg[664] <= 0;					r_cell_reg[665] <= 0;					r_cell_reg[666] <= 0;					r_cell_reg[667] <= 0;					r_cell_reg[668] <= 0;					r_cell_reg[669] <= 0;					r_cell_reg[670] <= 0;					r_cell_reg[671] <= 0;					r_cell_reg[672] <= 0;					r_cell_reg[673] <= 0;					r_cell_reg[674] <= 0;					r_cell_reg[675] <= 0;					r_cell_reg[676] <= 0;					r_cell_reg[677] <= 0;					r_cell_reg[678] <= 0;					r_cell_reg[679] <= 0;					r_cell_reg[680] <= 0;					r_cell_reg[681] <= 0;					r_cell_reg[682] <= 0;					r_cell_reg[683] <= 0;					r_cell_reg[684] <= 0;					r_cell_reg[685] <= 0;					r_cell_reg[686] <= 0;					r_cell_reg[687] <= 0;					r_cell_reg[688] <= 0;					r_cell_reg[689] <= 0;					r_cell_reg[690] <= 0;					r_cell_reg[691] <= 0;					r_cell_reg[692] <= 0;					r_cell_reg[693] <= 0;					r_cell_reg[694] <= 0;					r_cell_reg[695] <= 0;					r_cell_reg[696] <= 0;					r_cell_reg[697] <= 0;					r_cell_reg[698] <= 0;					r_cell_reg[699] <= 0;					r_cell_reg[700] <= 0;					r_cell_reg[701] <= 0;					r_cell_reg[702] <= 0;					r_cell_reg[703] <= 0;					r_cell_reg[704] <= 0;					r_cell_reg[705] <= 0;					r_cell_reg[706] <= 0;					r_cell_reg[707] <= 0;					r_cell_reg[708] <= 0;					r_cell_reg[709] <= 0;					r_cell_reg[710] <= 0;					r_cell_reg[711] <= 0;					r_cell_reg[712] <= 0;					r_cell_reg[713] <= 0;					r_cell_reg[714] <= 0;					r_cell_reg[715] <= 0;					r_cell_reg[716] <= 0;					r_cell_reg[717] <= 0;					r_cell_reg[718] <= 0;					r_cell_reg[719] <= 0;					r_cell_reg[720] <= 0;					r_cell_reg[721] <= 0;					r_cell_reg[722] <= 0;					r_cell_reg[723] <= 0;					r_cell_reg[724] <= 0;					r_cell_reg[725] <= 0;					r_cell_reg[726] <= 0;					r_cell_reg[727] <= 0;					r_cell_reg[728] <= 0;					r_cell_reg[729] <= 0;					r_cell_reg[730] <= 0;					r_cell_reg[731] <= 0;					r_cell_reg[732] <= 0;					r_cell_reg[733] <= 0;					r_cell_reg[734] <= 0;					r_cell_reg[735] <= 0;					r_cell_reg[736] <= 0;					r_cell_reg[737] <= 0;					r_cell_reg[738] <= 0;					r_cell_reg[739] <= 0;					r_cell_reg[740] <= 0;					r_cell_reg[741] <= 0;					r_cell_reg[742] <= 0;					r_cell_reg[743] <= 0;					r_cell_reg[744] <= 0;					r_cell_reg[745] <= 0;					r_cell_reg[746] <= 0;					r_cell_reg[747] <= 0;					r_cell_reg[748] <= 0;					r_cell_reg[749] <= 0;					r_cell_reg[750] <= 0;					r_cell_reg[751] <= 0;					r_cell_reg[752] <= 0;					r_cell_reg[753] <= 0;					r_cell_reg[754] <= 0;					r_cell_reg[755] <= 0;					r_cell_reg[756] <= 0;					r_cell_reg[757] <= 0;					r_cell_reg[758] <= 0;					r_cell_reg[759] <= 0;					r_cell_reg[760] <= 0;					r_cell_reg[761] <= 0;					r_cell_reg[762] <= 0;					r_cell_reg[763] <= 0;					r_cell_reg[764] <= 0;					r_cell_reg[765] <= 0;					r_cell_reg[766] <= 0;					r_cell_reg[767] <= 0;					r_cell_reg[768] <= 0;					r_cell_reg[769] <= 0;					r_cell_reg[770] <= 0;					r_cell_reg[771] <= 0;					r_cell_reg[772] <= 0;					r_cell_reg[773] <= 0;					r_cell_reg[774] <= 0;					r_cell_reg[775] <= 0;					r_cell_reg[776] <= 0;					r_cell_reg[777] <= 0;					r_cell_reg[778] <= 0;					r_cell_reg[779] <= 0;					r_cell_reg[780] <= 0;					r_cell_reg[781] <= 0;					r_cell_reg[782] <= 0;					r_cell_reg[783] <= 0;					r_cell_reg[784] <= 0;					r_cell_reg[785] <= 0;					r_cell_reg[786] <= 0;					r_cell_reg[787] <= 0;					r_cell_reg[788] <= 0;					r_cell_reg[789] <= 0;					r_cell_reg[790] <= 0;					r_cell_reg[791] <= 0;					r_cell_reg[792] <= 0;					r_cell_reg[793] <= 0;					r_cell_reg[794] <= 0;					r_cell_reg[795] <= 0;					r_cell_reg[796] <= 0;					r_cell_reg[797] <= 0;					r_cell_reg[798] <= 0;					r_cell_reg[799] <= 0;					r_cell_reg[800] <= 0;					r_cell_reg[801] <= 0;					r_cell_reg[802] <= 0;					r_cell_reg[803] <= 0;					r_cell_reg[804] <= 0;					r_cell_reg[805] <= 0;					r_cell_reg[806] <= 0;					r_cell_reg[807] <= 0;					r_cell_reg[808] <= 0;					r_cell_reg[809] <= 0;					r_cell_reg[810] <= 0;					r_cell_reg[811] <= 0;					r_cell_reg[812] <= 0;					r_cell_reg[813] <= 0;					r_cell_reg[814] <= 0;					r_cell_reg[815] <= 0;					r_cell_reg[816] <= 0;					r_cell_reg[817] <= 0;					r_cell_reg[818] <= 0;					r_cell_reg[819] <= 0;					r_cell_reg[820] <= 0;					r_cell_reg[821] <= 0;					r_cell_reg[822] <= 0;					r_cell_reg[823] <= 0;					r_cell_reg[824] <= 0;					r_cell_reg[825] <= 0;					r_cell_reg[826] <= 0;					r_cell_reg[827] <= 0;					r_cell_reg[828] <= 0;					r_cell_reg[829] <= 0;					r_cell_reg[830] <= 0;					r_cell_reg[831] <= 0;					r_cell_reg[832] <= 0;					r_cell_reg[833] <= 0;					r_cell_reg[834] <= 0;					r_cell_reg[835] <= 0;					r_cell_reg[836] <= 0;					r_cell_reg[837] <= 0;					r_cell_reg[838] <= 0;					r_cell_reg[839] <= 0;					r_cell_reg[840] <= 0;					r_cell_reg[841] <= 0;					r_cell_reg[842] <= 0;					r_cell_reg[843] <= 0;					r_cell_reg[844] <= 0;					r_cell_reg[845] <= 0;					r_cell_reg[846] <= 0;					r_cell_reg[847] <= 0;					r_cell_reg[848] <= 0;					r_cell_reg[849] <= 0;					r_cell_reg[850] <= 0;					r_cell_reg[851] <= 0;					r_cell_reg[852] <= 0;					r_cell_reg[853] <= 0;					r_cell_reg[854] <= 0;					r_cell_reg[855] <= 0;					r_cell_reg[856] <= 0;					r_cell_reg[857] <= 0;					r_cell_reg[858] <= 0;					r_cell_reg[859] <= 0;					r_cell_reg[860] <= 0;					r_cell_reg[861] <= 0;					r_cell_reg[862] <= 0;					r_cell_reg[863] <= 0;					r_cell_reg[864] <= 0;					r_cell_reg[865] <= 0;					r_cell_reg[866] <= 0;					r_cell_reg[867] <= 0;					r_cell_reg[868] <= 0;					r_cell_reg[869] <= 0;					r_cell_reg[870] <= 0;					r_cell_reg[871] <= 0;					r_cell_reg[872] <= 0;					r_cell_reg[873] <= 0;					r_cell_reg[874] <= 0;					r_cell_reg[875] <= 0;					r_cell_reg[876] <= 0;					r_cell_reg[877] <= 0;					r_cell_reg[878] <= 0;					r_cell_reg[879] <= 0;					r_cell_reg[880] <= 0;					r_cell_reg[881] <= 0;					r_cell_reg[882] <= 0;					r_cell_reg[883] <= 0;					r_cell_reg[884] <= 0;					r_cell_reg[885] <= 0;					r_cell_reg[886] <= 0;					r_cell_reg[887] <= 0;					r_cell_reg[888] <= 0;					r_cell_reg[889] <= 0;					r_cell_reg[890] <= 0;					r_cell_reg[891] <= 0;					r_cell_reg[892] <= 0;					r_cell_reg[893] <= 0;					r_cell_reg[894] <= 0;					r_cell_reg[895] <= 0;					r_cell_reg[896] <= 0;					r_cell_reg[897] <= 0;					r_cell_reg[898] <= 0;					r_cell_reg[899] <= 0;					r_cell_reg[900] <= 0;					r_cell_reg[901] <= 0;					r_cell_reg[902] <= 0;					r_cell_reg[903] <= 0;					r_cell_reg[904] <= 0;					r_cell_reg[905] <= 0;					r_cell_reg[906] <= 0;					r_cell_reg[907] <= 0;					r_cell_reg[908] <= 0;					r_cell_reg[909] <= 0;					r_cell_reg[910] <= 0;					r_cell_reg[911] <= 0;					r_cell_reg[912] <= 0;					r_cell_reg[913] <= 0;					r_cell_reg[914] <= 0;					r_cell_reg[915] <= 0;					r_cell_reg[916] <= 0;					r_cell_reg[917] <= 0;					r_cell_reg[918] <= 0;					r_cell_reg[919] <= 0;					r_cell_reg[920] <= 0;					r_cell_reg[921] <= 0;					r_cell_reg[922] <= 0;					r_cell_reg[923] <= 0;					r_cell_reg[924] <= 0;					r_cell_reg[925] <= 0;					r_cell_reg[926] <= 0;					r_cell_reg[927] <= 0;					r_cell_reg[928] <= 0;					r_cell_reg[929] <= 0;					r_cell_reg[930] <= 0;					r_cell_reg[931] <= 0;					r_cell_reg[932] <= 0;					r_cell_reg[933] <= 0;					r_cell_reg[934] <= 0;					r_cell_reg[935] <= 0;					r_cell_reg[936] <= 0;					r_cell_reg[937] <= 0;					r_cell_reg[938] <= 0;					r_cell_reg[939] <= 0;					r_cell_reg[940] <= 0;					r_cell_reg[941] <= 0;					r_cell_reg[942] <= 0;					r_cell_reg[943] <= 0;					r_cell_reg[944] <= 0;					r_cell_reg[945] <= 0;					r_cell_reg[946] <= 0;					r_cell_reg[947] <= 0;					r_cell_reg[948] <= 0;					r_cell_reg[949] <= 0;					r_cell_reg[950] <= 0;					r_cell_reg[951] <= 0;					r_cell_reg[952] <= 0;					r_cell_reg[953] <= 0;					r_cell_reg[954] <= 0;					r_cell_reg[955] <= 0;					r_cell_reg[956] <= 0;					r_cell_reg[957] <= 0;					r_cell_reg[958] <= 0;					r_cell_reg[959] <= 0;					r_cell_reg[960] <= 0;					r_cell_reg[961] <= 0;					r_cell_reg[962] <= 0;					r_cell_reg[963] <= 0;					r_cell_reg[964] <= 0;					r_cell_reg[965] <= 0;					r_cell_reg[966] <= 0;					r_cell_reg[967] <= 0;					r_cell_reg[968] <= 0;					r_cell_reg[969] <= 0;					r_cell_reg[970] <= 0;					r_cell_reg[971] <= 0;					r_cell_reg[972] <= 0;					r_cell_reg[973] <= 0;					r_cell_reg[974] <= 0;					r_cell_reg[975] <= 0;					r_cell_reg[976] <= 0;					r_cell_reg[977] <= 0;					r_cell_reg[978] <= 0;					r_cell_reg[979] <= 0;					r_cell_reg[980] <= 0;					r_cell_reg[981] <= 0;					r_cell_reg[982] <= 0;					r_cell_reg[983] <= 0;					r_cell_reg[984] <= 0;					r_cell_reg[985] <= 0;					r_cell_reg[986] <= 0;					r_cell_reg[987] <= 0;					r_cell_reg[988] <= 0;					r_cell_reg[989] <= 0;					r_cell_reg[990] <= 0;					r_cell_reg[991] <= 0;					r_cell_reg[992] <= 0;					r_cell_reg[993] <= 0;					r_cell_reg[994] <= 0;					r_cell_reg[995] <= 0;					r_cell_reg[996] <= 0;					r_cell_reg[997] <= 0;					r_cell_reg[998] <= 0;					r_cell_reg[999] <= 0;					r_cell_reg[1000] <= 0;					r_cell_reg[1001] <= 0;					r_cell_reg[1002] <= 0;					r_cell_reg[1003] <= 0;					r_cell_reg[1004] <= 0;					r_cell_reg[1005] <= 0;					r_cell_reg[1006] <= 0;					r_cell_reg[1007] <= 0;					r_cell_reg[1008] <= 0;					r_cell_reg[1009] <= 0;					r_cell_reg[1010] <= 0;					r_cell_reg[1011] <= 0;					r_cell_reg[1012] <= 0;					r_cell_reg[1013] <= 0;					r_cell_reg[1014] <= 0;					r_cell_reg[1015] <= 0;					r_cell_reg[1016] <= 0;					r_cell_reg[1017] <= 0;					r_cell_reg[1018] <= 0;					r_cell_reg[1019] <= 0;					r_cell_reg[1020] <= 0;					r_cell_reg[1021] <= 0;					r_cell_reg[1022] <= 0;					r_cell_reg[1023] <= 0;					l_cell_reg[0] <= 0;					l_cell_reg[1] <= 0;					l_cell_reg[2] <= 0;					l_cell_reg[3] <= 0;					l_cell_reg[4] <= 0;					l_cell_reg[5] <= 0;					l_cell_reg[6] <= 0;					l_cell_reg[7] <= 0;					l_cell_reg[8] <= 0;					l_cell_reg[9] <= 0;					l_cell_reg[10] <= 0;					l_cell_reg[11] <= 0;					l_cell_reg[12] <= 0;					l_cell_reg[13] <= 0;					l_cell_reg[14] <= 0;					l_cell_reg[15] <= 0;					l_cell_reg[16] <= 0;					l_cell_reg[17] <= 0;					l_cell_reg[18] <= 0;					l_cell_reg[19] <= 0;					l_cell_reg[20] <= 0;					l_cell_reg[21] <= 0;					l_cell_reg[22] <= 0;					l_cell_reg[23] <= 0;					l_cell_reg[24] <= 0;					l_cell_reg[25] <= 0;					l_cell_reg[26] <= 0;					l_cell_reg[27] <= 0;					l_cell_reg[28] <= 0;					l_cell_reg[29] <= 0;					l_cell_reg[30] <= 0;					l_cell_reg[31] <= 0;					l_cell_reg[32] <= 0;					l_cell_reg[33] <= 0;					l_cell_reg[34] <= 0;					l_cell_reg[35] <= 0;					l_cell_reg[36] <= 0;					l_cell_reg[37] <= 0;					l_cell_reg[38] <= 0;					l_cell_reg[39] <= 0;					l_cell_reg[40] <= 0;					l_cell_reg[41] <= 0;					l_cell_reg[42] <= 0;					l_cell_reg[43] <= 0;					l_cell_reg[44] <= 0;					l_cell_reg[45] <= 0;					l_cell_reg[46] <= 0;					l_cell_reg[47] <= 0;					l_cell_reg[48] <= 0;					l_cell_reg[49] <= 0;					l_cell_reg[50] <= 0;					l_cell_reg[51] <= 0;					l_cell_reg[52] <= 0;					l_cell_reg[53] <= 0;					l_cell_reg[54] <= 0;					l_cell_reg[55] <= 0;					l_cell_reg[56] <= 0;					l_cell_reg[57] <= 0;					l_cell_reg[58] <= 0;					l_cell_reg[59] <= 0;					l_cell_reg[60] <= 0;					l_cell_reg[61] <= 0;					l_cell_reg[62] <= 0;					l_cell_reg[63] <= 0;					l_cell_reg[64] <= 0;					l_cell_reg[65] <= 0;					l_cell_reg[66] <= 0;					l_cell_reg[67] <= 0;					l_cell_reg[68] <= 0;					l_cell_reg[69] <= 0;					l_cell_reg[70] <= 0;					l_cell_reg[71] <= 0;					l_cell_reg[72] <= 0;					l_cell_reg[73] <= 0;					l_cell_reg[74] <= 0;					l_cell_reg[75] <= 0;					l_cell_reg[76] <= 0;					l_cell_reg[77] <= 0;					l_cell_reg[78] <= 0;					l_cell_reg[79] <= 0;					l_cell_reg[80] <= 0;					l_cell_reg[81] <= 0;					l_cell_reg[82] <= 0;					l_cell_reg[83] <= 0;					l_cell_reg[84] <= 0;					l_cell_reg[85] <= 0;					l_cell_reg[86] <= 0;					l_cell_reg[87] <= 0;					l_cell_reg[88] <= 0;					l_cell_reg[89] <= 0;					l_cell_reg[90] <= 0;					l_cell_reg[91] <= 0;					l_cell_reg[92] <= 0;					l_cell_reg[93] <= 0;					l_cell_reg[94] <= 0;					l_cell_reg[95] <= 0;					l_cell_reg[96] <= 0;					l_cell_reg[97] <= 0;					l_cell_reg[98] <= 0;					l_cell_reg[99] <= 0;					l_cell_reg[100] <= 0;					l_cell_reg[101] <= 0;					l_cell_reg[102] <= 0;					l_cell_reg[103] <= 0;					l_cell_reg[104] <= 0;					l_cell_reg[105] <= 0;					l_cell_reg[106] <= 0;					l_cell_reg[107] <= 0;					l_cell_reg[108] <= 0;					l_cell_reg[109] <= 0;					l_cell_reg[110] <= 0;					l_cell_reg[111] <= 0;					l_cell_reg[112] <= 0;					l_cell_reg[113] <= 0;					l_cell_reg[114] <= 0;					l_cell_reg[115] <= 0;					l_cell_reg[116] <= 0;					l_cell_reg[117] <= 0;					l_cell_reg[118] <= 0;					l_cell_reg[119] <= 0;					l_cell_reg[120] <= 0;					l_cell_reg[121] <= 0;					l_cell_reg[122] <= 0;					l_cell_reg[123] <= 0;					l_cell_reg[124] <= 0;					l_cell_reg[125] <= 0;					l_cell_reg[126] <= 0;					l_cell_reg[127] <= 0;					l_cell_reg[128] <= 0;					l_cell_reg[129] <= 0;					l_cell_reg[130] <= 0;					l_cell_reg[131] <= 0;					l_cell_reg[132] <= 0;					l_cell_reg[133] <= 0;					l_cell_reg[134] <= 0;					l_cell_reg[135] <= 0;					l_cell_reg[136] <= 0;					l_cell_reg[137] <= 0;					l_cell_reg[138] <= 0;					l_cell_reg[139] <= 0;					l_cell_reg[140] <= 0;					l_cell_reg[141] <= 0;					l_cell_reg[142] <= 0;					l_cell_reg[143] <= 0;					l_cell_reg[144] <= 0;					l_cell_reg[145] <= 0;					l_cell_reg[146] <= 0;					l_cell_reg[147] <= 0;					l_cell_reg[148] <= 0;					l_cell_reg[149] <= 0;					l_cell_reg[150] <= 0;					l_cell_reg[151] <= 0;					l_cell_reg[152] <= 0;					l_cell_reg[153] <= 0;					l_cell_reg[154] <= 0;					l_cell_reg[155] <= 0;					l_cell_reg[156] <= 0;					l_cell_reg[157] <= 0;					l_cell_reg[158] <= 0;					l_cell_reg[159] <= 0;					l_cell_reg[160] <= 0;					l_cell_reg[161] <= 0;					l_cell_reg[162] <= 0;					l_cell_reg[163] <= 0;					l_cell_reg[164] <= 0;					l_cell_reg[165] <= 0;					l_cell_reg[166] <= 0;					l_cell_reg[167] <= 0;					l_cell_reg[168] <= 0;					l_cell_reg[169] <= 0;					l_cell_reg[170] <= 0;					l_cell_reg[171] <= 0;					l_cell_reg[172] <= 0;					l_cell_reg[173] <= 0;					l_cell_reg[174] <= 0;					l_cell_reg[175] <= 0;					l_cell_reg[176] <= 0;					l_cell_reg[177] <= 0;					l_cell_reg[178] <= 0;					l_cell_reg[179] <= 0;					l_cell_reg[180] <= 0;					l_cell_reg[181] <= 0;					l_cell_reg[182] <= 0;					l_cell_reg[183] <= 0;					l_cell_reg[184] <= 0;					l_cell_reg[185] <= 0;					l_cell_reg[186] <= 0;					l_cell_reg[187] <= 0;					l_cell_reg[188] <= 0;					l_cell_reg[189] <= 0;					l_cell_reg[190] <= 0;					l_cell_reg[191] <= 0;					l_cell_reg[192] <= 0;					l_cell_reg[193] <= 0;					l_cell_reg[194] <= 0;					l_cell_reg[195] <= 0;					l_cell_reg[196] <= 0;					l_cell_reg[197] <= 0;					l_cell_reg[198] <= 0;					l_cell_reg[199] <= 0;					l_cell_reg[200] <= 0;					l_cell_reg[201] <= 0;					l_cell_reg[202] <= 0;					l_cell_reg[203] <= 0;					l_cell_reg[204] <= 0;					l_cell_reg[205] <= 0;					l_cell_reg[206] <= 0;					l_cell_reg[207] <= 0;					l_cell_reg[208] <= 0;					l_cell_reg[209] <= 0;					l_cell_reg[210] <= 0;					l_cell_reg[211] <= 0;					l_cell_reg[212] <= 0;					l_cell_reg[213] <= 0;					l_cell_reg[214] <= 0;					l_cell_reg[215] <= 0;					l_cell_reg[216] <= 0;					l_cell_reg[217] <= 0;					l_cell_reg[218] <= 0;					l_cell_reg[219] <= 0;					l_cell_reg[220] <= 0;					l_cell_reg[221] <= 0;					l_cell_reg[222] <= 0;					l_cell_reg[223] <= 0;					l_cell_reg[224] <= 0;					l_cell_reg[225] <= 0;					l_cell_reg[226] <= 0;					l_cell_reg[227] <= 0;					l_cell_reg[228] <= 0;					l_cell_reg[229] <= 0;					l_cell_reg[230] <= 0;					l_cell_reg[231] <= 0;					l_cell_reg[232] <= 0;					l_cell_reg[233] <= 0;					l_cell_reg[234] <= 0;					l_cell_reg[235] <= 0;					l_cell_reg[236] <= 0;					l_cell_reg[237] <= 0;					l_cell_reg[238] <= 0;					l_cell_reg[239] <= 0;					l_cell_reg[240] <= 0;					l_cell_reg[241] <= 0;					l_cell_reg[242] <= 0;					l_cell_reg[243] <= 0;					l_cell_reg[244] <= 0;					l_cell_reg[245] <= 0;					l_cell_reg[246] <= 0;					l_cell_reg[247] <= 0;					l_cell_reg[248] <= 0;					l_cell_reg[249] <= 0;					l_cell_reg[250] <= 0;					l_cell_reg[251] <= 0;					l_cell_reg[252] <= 0;					l_cell_reg[253] <= 0;					l_cell_reg[254] <= 0;					l_cell_reg[255] <= 0;					l_cell_reg[256] <= 0;					l_cell_reg[257] <= 0;					l_cell_reg[258] <= 0;					l_cell_reg[259] <= 0;					l_cell_reg[260] <= 0;					l_cell_reg[261] <= 0;					l_cell_reg[262] <= 0;					l_cell_reg[263] <= 0;					l_cell_reg[264] <= 0;					l_cell_reg[265] <= 0;					l_cell_reg[266] <= 0;					l_cell_reg[267] <= 0;					l_cell_reg[268] <= 0;					l_cell_reg[269] <= 0;					l_cell_reg[270] <= 0;					l_cell_reg[271] <= 0;					l_cell_reg[272] <= 0;					l_cell_reg[273] <= 0;					l_cell_reg[274] <= 0;					l_cell_reg[275] <= 0;					l_cell_reg[276] <= 0;					l_cell_reg[277] <= 0;					l_cell_reg[278] <= 0;					l_cell_reg[279] <= 0;					l_cell_reg[280] <= 0;					l_cell_reg[281] <= 0;					l_cell_reg[282] <= 0;					l_cell_reg[283] <= 0;					l_cell_reg[284] <= 0;					l_cell_reg[285] <= 0;					l_cell_reg[286] <= 0;					l_cell_reg[287] <= 0;					l_cell_reg[288] <= 0;					l_cell_reg[289] <= 0;					l_cell_reg[290] <= 0;					l_cell_reg[291] <= 0;					l_cell_reg[292] <= 0;					l_cell_reg[293] <= 0;					l_cell_reg[294] <= 0;					l_cell_reg[295] <= 0;					l_cell_reg[296] <= 0;					l_cell_reg[297] <= 0;					l_cell_reg[298] <= 0;					l_cell_reg[299] <= 0;					l_cell_reg[300] <= 0;					l_cell_reg[301] <= 0;					l_cell_reg[302] <= 0;					l_cell_reg[303] <= 0;					l_cell_reg[304] <= 0;					l_cell_reg[305] <= 0;					l_cell_reg[306] <= 0;					l_cell_reg[307] <= 0;					l_cell_reg[308] <= 0;					l_cell_reg[309] <= 0;					l_cell_reg[310] <= 0;					l_cell_reg[311] <= 0;					l_cell_reg[312] <= 0;					l_cell_reg[313] <= 0;					l_cell_reg[314] <= 0;					l_cell_reg[315] <= 0;					l_cell_reg[316] <= 0;					l_cell_reg[317] <= 0;					l_cell_reg[318] <= 0;					l_cell_reg[319] <= 0;					l_cell_reg[320] <= 0;					l_cell_reg[321] <= 0;					l_cell_reg[322] <= 0;					l_cell_reg[323] <= 0;					l_cell_reg[324] <= 0;					l_cell_reg[325] <= 0;					l_cell_reg[326] <= 0;					l_cell_reg[327] <= 0;					l_cell_reg[328] <= 0;					l_cell_reg[329] <= 0;					l_cell_reg[330] <= 0;					l_cell_reg[331] <= 0;					l_cell_reg[332] <= 0;					l_cell_reg[333] <= 0;					l_cell_reg[334] <= 0;					l_cell_reg[335] <= 0;					l_cell_reg[336] <= 0;					l_cell_reg[337] <= 0;					l_cell_reg[338] <= 0;					l_cell_reg[339] <= 0;					l_cell_reg[340] <= 0;					l_cell_reg[341] <= 0;					l_cell_reg[342] <= 0;					l_cell_reg[343] <= 0;					l_cell_reg[344] <= 0;					l_cell_reg[345] <= 0;					l_cell_reg[346] <= 0;					l_cell_reg[347] <= 0;					l_cell_reg[348] <= 0;					l_cell_reg[349] <= 0;					l_cell_reg[350] <= 0;					l_cell_reg[351] <= 0;					l_cell_reg[352] <= 0;					l_cell_reg[353] <= 0;					l_cell_reg[354] <= 0;					l_cell_reg[355] <= 0;					l_cell_reg[356] <= 0;					l_cell_reg[357] <= 0;					l_cell_reg[358] <= 0;					l_cell_reg[359] <= 0;					l_cell_reg[360] <= 0;					l_cell_reg[361] <= 0;					l_cell_reg[362] <= 0;					l_cell_reg[363] <= 0;					l_cell_reg[364] <= 0;					l_cell_reg[365] <= 0;					l_cell_reg[366] <= 0;					l_cell_reg[367] <= 0;					l_cell_reg[368] <= 0;					l_cell_reg[369] <= 0;					l_cell_reg[370] <= 0;					l_cell_reg[371] <= 0;					l_cell_reg[372] <= 0;					l_cell_reg[373] <= 0;					l_cell_reg[374] <= 0;					l_cell_reg[375] <= 0;					l_cell_reg[376] <= 0;					l_cell_reg[377] <= 0;					l_cell_reg[378] <= 0;					l_cell_reg[379] <= 0;					l_cell_reg[380] <= 0;					l_cell_reg[381] <= 0;					l_cell_reg[382] <= 0;					l_cell_reg[383] <= 0;					l_cell_reg[384] <= 0;					l_cell_reg[385] <= 0;					l_cell_reg[386] <= 0;					l_cell_reg[387] <= 0;					l_cell_reg[388] <= 0;					l_cell_reg[389] <= 0;					l_cell_reg[390] <= 0;					l_cell_reg[391] <= 0;					l_cell_reg[392] <= 0;					l_cell_reg[393] <= 0;					l_cell_reg[394] <= 0;					l_cell_reg[395] <= 0;					l_cell_reg[396] <= 0;					l_cell_reg[397] <= 0;					l_cell_reg[398] <= 0;					l_cell_reg[399] <= 0;					l_cell_reg[400] <= 0;					l_cell_reg[401] <= 0;					l_cell_reg[402] <= 0;					l_cell_reg[403] <= 0;					l_cell_reg[404] <= 0;					l_cell_reg[405] <= 0;					l_cell_reg[406] <= 0;					l_cell_reg[407] <= 0;					l_cell_reg[408] <= 0;					l_cell_reg[409] <= 0;					l_cell_reg[410] <= 0;					l_cell_reg[411] <= 0;					l_cell_reg[412] <= 0;					l_cell_reg[413] <= 0;					l_cell_reg[414] <= 0;					l_cell_reg[415] <= 0;					l_cell_reg[416] <= 0;					l_cell_reg[417] <= 0;					l_cell_reg[418] <= 0;					l_cell_reg[419] <= 0;					l_cell_reg[420] <= 0;					l_cell_reg[421] <= 0;					l_cell_reg[422] <= 0;					l_cell_reg[423] <= 0;					l_cell_reg[424] <= 0;					l_cell_reg[425] <= 0;					l_cell_reg[426] <= 0;					l_cell_reg[427] <= 0;					l_cell_reg[428] <= 0;					l_cell_reg[429] <= 0;					l_cell_reg[430] <= 0;					l_cell_reg[431] <= 0;					l_cell_reg[432] <= 0;					l_cell_reg[433] <= 0;					l_cell_reg[434] <= 0;					l_cell_reg[435] <= 0;					l_cell_reg[436] <= 0;					l_cell_reg[437] <= 0;					l_cell_reg[438] <= 0;					l_cell_reg[439] <= 0;					l_cell_reg[440] <= 0;					l_cell_reg[441] <= 0;					l_cell_reg[442] <= 0;					l_cell_reg[443] <= 0;					l_cell_reg[444] <= 0;					l_cell_reg[445] <= 0;					l_cell_reg[446] <= 0;					l_cell_reg[447] <= 0;					l_cell_reg[448] <= 0;					l_cell_reg[449] <= 0;					l_cell_reg[450] <= 0;					l_cell_reg[451] <= 0;					l_cell_reg[452] <= 0;					l_cell_reg[453] <= 0;					l_cell_reg[454] <= 0;					l_cell_reg[455] <= 0;					l_cell_reg[456] <= 0;					l_cell_reg[457] <= 0;					l_cell_reg[458] <= 0;					l_cell_reg[459] <= 0;					l_cell_reg[460] <= 0;					l_cell_reg[461] <= 0;					l_cell_reg[462] <= 0;					l_cell_reg[463] <= 0;					l_cell_reg[464] <= 0;					l_cell_reg[465] <= 0;					l_cell_reg[466] <= 0;					l_cell_reg[467] <= 0;					l_cell_reg[468] <= 0;					l_cell_reg[469] <= 0;					l_cell_reg[470] <= 0;					l_cell_reg[471] <= 0;					l_cell_reg[472] <= 0;					l_cell_reg[473] <= 0;					l_cell_reg[474] <= 0;					l_cell_reg[475] <= 0;					l_cell_reg[476] <= 0;					l_cell_reg[477] <= 0;					l_cell_reg[478] <= 0;					l_cell_reg[479] <= 0;					l_cell_reg[480] <= 0;					l_cell_reg[481] <= 0;					l_cell_reg[482] <= 0;					l_cell_reg[483] <= 0;					l_cell_reg[484] <= 0;					l_cell_reg[485] <= 0;					l_cell_reg[486] <= 0;					l_cell_reg[487] <= 0;					l_cell_reg[488] <= 0;					l_cell_reg[489] <= 0;					l_cell_reg[490] <= 0;					l_cell_reg[491] <= 0;					l_cell_reg[492] <= 0;					l_cell_reg[493] <= 0;					l_cell_reg[494] <= 0;					l_cell_reg[495] <= 0;					l_cell_reg[496] <= 0;					l_cell_reg[497] <= 0;					l_cell_reg[498] <= 0;					l_cell_reg[499] <= 0;					l_cell_reg[500] <= 0;					l_cell_reg[501] <= 0;					l_cell_reg[502] <= 0;					l_cell_reg[503] <= 0;					l_cell_reg[504] <= 0;					l_cell_reg[505] <= 0;					l_cell_reg[506] <= 0;					l_cell_reg[507] <= 0;					l_cell_reg[508] <= 0;					l_cell_reg[509] <= 0;					l_cell_reg[510] <= 0;					l_cell_reg[511] <= 0;					l_cell_reg[512] <= 0;					l_cell_reg[513] <= 0;					l_cell_reg[514] <= 0;					l_cell_reg[515] <= 0;					l_cell_reg[516] <= 0;					l_cell_reg[517] <= 0;					l_cell_reg[518] <= 0;					l_cell_reg[519] <= 0;					l_cell_reg[520] <= 0;					l_cell_reg[521] <= 0;					l_cell_reg[522] <= 0;					l_cell_reg[523] <= 0;					l_cell_reg[524] <= 0;					l_cell_reg[525] <= 0;					l_cell_reg[526] <= 0;					l_cell_reg[527] <= 0;					l_cell_reg[528] <= 0;					l_cell_reg[529] <= 0;					l_cell_reg[530] <= 0;					l_cell_reg[531] <= 0;					l_cell_reg[532] <= 0;					l_cell_reg[533] <= 0;					l_cell_reg[534] <= 0;					l_cell_reg[535] <= 0;					l_cell_reg[536] <= 0;					l_cell_reg[537] <= 0;					l_cell_reg[538] <= 0;					l_cell_reg[539] <= 0;					l_cell_reg[540] <= 0;					l_cell_reg[541] <= 0;					l_cell_reg[542] <= 0;					l_cell_reg[543] <= 0;					l_cell_reg[544] <= 0;					l_cell_reg[545] <= 0;					l_cell_reg[546] <= 0;					l_cell_reg[547] <= 0;					l_cell_reg[548] <= 0;					l_cell_reg[549] <= 0;					l_cell_reg[550] <= 0;					l_cell_reg[551] <= 0;					l_cell_reg[552] <= 0;					l_cell_reg[553] <= 0;					l_cell_reg[554] <= 0;					l_cell_reg[555] <= 0;					l_cell_reg[556] <= 0;					l_cell_reg[557] <= 0;					l_cell_reg[558] <= 0;					l_cell_reg[559] <= 0;					l_cell_reg[560] <= 0;					l_cell_reg[561] <= 0;					l_cell_reg[562] <= 0;					l_cell_reg[563] <= 0;					l_cell_reg[564] <= 0;					l_cell_reg[565] <= 0;					l_cell_reg[566] <= 0;					l_cell_reg[567] <= 0;					l_cell_reg[568] <= 0;					l_cell_reg[569] <= 0;					l_cell_reg[570] <= 0;					l_cell_reg[571] <= 0;					l_cell_reg[572] <= 0;					l_cell_reg[573] <= 0;					l_cell_reg[574] <= 0;					l_cell_reg[575] <= 0;					l_cell_reg[576] <= 0;					l_cell_reg[577] <= 0;					l_cell_reg[578] <= 0;					l_cell_reg[579] <= 0;					l_cell_reg[580] <= 0;					l_cell_reg[581] <= 0;					l_cell_reg[582] <= 0;					l_cell_reg[583] <= 0;					l_cell_reg[584] <= 0;					l_cell_reg[585] <= 0;					l_cell_reg[586] <= 0;					l_cell_reg[587] <= 0;					l_cell_reg[588] <= 0;					l_cell_reg[589] <= 0;					l_cell_reg[590] <= 0;					l_cell_reg[591] <= 0;					l_cell_reg[592] <= 0;					l_cell_reg[593] <= 0;					l_cell_reg[594] <= 0;					l_cell_reg[595] <= 0;					l_cell_reg[596] <= 0;					l_cell_reg[597] <= 0;					l_cell_reg[598] <= 0;					l_cell_reg[599] <= 0;					l_cell_reg[600] <= 0;					l_cell_reg[601] <= 0;					l_cell_reg[602] <= 0;					l_cell_reg[603] <= 0;					l_cell_reg[604] <= 0;					l_cell_reg[605] <= 0;					l_cell_reg[606] <= 0;					l_cell_reg[607] <= 0;					l_cell_reg[608] <= 0;					l_cell_reg[609] <= 0;					l_cell_reg[610] <= 0;					l_cell_reg[611] <= 0;					l_cell_reg[612] <= 0;					l_cell_reg[613] <= 0;					l_cell_reg[614] <= 0;					l_cell_reg[615] <= 0;					l_cell_reg[616] <= 0;					l_cell_reg[617] <= 0;					l_cell_reg[618] <= 0;					l_cell_reg[619] <= 0;					l_cell_reg[620] <= 0;					l_cell_reg[621] <= 0;					l_cell_reg[622] <= 0;					l_cell_reg[623] <= 0;					l_cell_reg[624] <= 0;					l_cell_reg[625] <= 0;					l_cell_reg[626] <= 0;					l_cell_reg[627] <= 0;					l_cell_reg[628] <= 0;					l_cell_reg[629] <= 0;					l_cell_reg[630] <= 0;					l_cell_reg[631] <= 0;					l_cell_reg[632] <= 0;					l_cell_reg[633] <= 0;					l_cell_reg[634] <= 0;					l_cell_reg[635] <= 0;					l_cell_reg[636] <= 0;					l_cell_reg[637] <= 0;					l_cell_reg[638] <= 0;					l_cell_reg[639] <= 0;					l_cell_reg[640] <= 0;					l_cell_reg[641] <= 0;					l_cell_reg[642] <= 0;					l_cell_reg[643] <= 0;					l_cell_reg[644] <= 0;					l_cell_reg[645] <= 0;					l_cell_reg[646] <= 0;					l_cell_reg[647] <= 0;					l_cell_reg[648] <= 0;					l_cell_reg[649] <= 0;					l_cell_reg[650] <= 0;					l_cell_reg[651] <= 0;					l_cell_reg[652] <= 0;					l_cell_reg[653] <= 0;					l_cell_reg[654] <= 0;					l_cell_reg[655] <= 0;					l_cell_reg[656] <= 0;					l_cell_reg[657] <= 0;					l_cell_reg[658] <= 0;					l_cell_reg[659] <= 0;					l_cell_reg[660] <= 0;					l_cell_reg[661] <= 0;					l_cell_reg[662] <= 0;					l_cell_reg[663] <= 0;					l_cell_reg[664] <= 0;					l_cell_reg[665] <= 0;					l_cell_reg[666] <= 0;					l_cell_reg[667] <= 0;					l_cell_reg[668] <= 0;					l_cell_reg[669] <= 0;					l_cell_reg[670] <= 0;					l_cell_reg[671] <= 0;					l_cell_reg[672] <= 0;					l_cell_reg[673] <= 0;					l_cell_reg[674] <= 0;					l_cell_reg[675] <= 0;					l_cell_reg[676] <= 0;					l_cell_reg[677] <= 0;					l_cell_reg[678] <= 0;					l_cell_reg[679] <= 0;					l_cell_reg[680] <= 0;					l_cell_reg[681] <= 0;					l_cell_reg[682] <= 0;					l_cell_reg[683] <= 0;					l_cell_reg[684] <= 0;					l_cell_reg[685] <= 0;					l_cell_reg[686] <= 0;					l_cell_reg[687] <= 0;					l_cell_reg[688] <= 0;					l_cell_reg[689] <= 0;					l_cell_reg[690] <= 0;					l_cell_reg[691] <= 0;					l_cell_reg[692] <= 0;					l_cell_reg[693] <= 0;					l_cell_reg[694] <= 0;					l_cell_reg[695] <= 0;					l_cell_reg[696] <= 0;					l_cell_reg[697] <= 0;					l_cell_reg[698] <= 0;					l_cell_reg[699] <= 0;					l_cell_reg[700] <= 0;					l_cell_reg[701] <= 0;					l_cell_reg[702] <= 0;					l_cell_reg[703] <= 0;					l_cell_reg[704] <= 0;					l_cell_reg[705] <= 0;					l_cell_reg[706] <= 0;					l_cell_reg[707] <= 0;					l_cell_reg[708] <= 0;					l_cell_reg[709] <= 0;					l_cell_reg[710] <= 0;					l_cell_reg[711] <= 0;					l_cell_reg[712] <= 0;					l_cell_reg[713] <= 0;					l_cell_reg[714] <= 0;					l_cell_reg[715] <= 0;					l_cell_reg[716] <= 0;					l_cell_reg[717] <= 0;					l_cell_reg[718] <= 0;					l_cell_reg[719] <= 0;					l_cell_reg[720] <= 0;					l_cell_reg[721] <= 0;					l_cell_reg[722] <= 0;					l_cell_reg[723] <= 0;					l_cell_reg[724] <= 0;					l_cell_reg[725] <= 0;					l_cell_reg[726] <= 0;					l_cell_reg[727] <= 0;					l_cell_reg[728] <= 0;					l_cell_reg[729] <= 0;					l_cell_reg[730] <= 0;					l_cell_reg[731] <= 0;					l_cell_reg[732] <= 0;					l_cell_reg[733] <= 0;					l_cell_reg[734] <= 0;					l_cell_reg[735] <= 0;					l_cell_reg[736] <= 0;					l_cell_reg[737] <= 0;					l_cell_reg[738] <= 0;					l_cell_reg[739] <= 0;					l_cell_reg[740] <= 0;					l_cell_reg[741] <= 0;					l_cell_reg[742] <= 0;					l_cell_reg[743] <= 0;					l_cell_reg[744] <= 0;					l_cell_reg[745] <= 0;					l_cell_reg[746] <= 0;					l_cell_reg[747] <= 0;					l_cell_reg[748] <= 0;					l_cell_reg[749] <= 0;					l_cell_reg[750] <= 0;					l_cell_reg[751] <= 0;					l_cell_reg[752] <= 0;					l_cell_reg[753] <= 0;					l_cell_reg[754] <= 0;					l_cell_reg[755] <= 0;					l_cell_reg[756] <= 0;					l_cell_reg[757] <= 0;					l_cell_reg[758] <= 0;					l_cell_reg[759] <= 0;					l_cell_reg[760] <= 0;					l_cell_reg[761] <= 0;					l_cell_reg[762] <= 0;					l_cell_reg[763] <= 0;					l_cell_reg[764] <= 0;					l_cell_reg[765] <= 0;					l_cell_reg[766] <= 0;					l_cell_reg[767] <= 0;					l_cell_reg[768] <= 0;					l_cell_reg[769] <= 0;					l_cell_reg[770] <= 0;					l_cell_reg[771] <= 0;					l_cell_reg[772] <= 0;					l_cell_reg[773] <= 0;					l_cell_reg[774] <= 0;					l_cell_reg[775] <= 0;					l_cell_reg[776] <= 0;					l_cell_reg[777] <= 0;					l_cell_reg[778] <= 0;					l_cell_reg[779] <= 0;					l_cell_reg[780] <= 0;					l_cell_reg[781] <= 0;					l_cell_reg[782] <= 0;					l_cell_reg[783] <= 0;					l_cell_reg[784] <= 0;					l_cell_reg[785] <= 0;					l_cell_reg[786] <= 0;					l_cell_reg[787] <= 0;					l_cell_reg[788] <= 0;					l_cell_reg[789] <= 0;					l_cell_reg[790] <= 0;					l_cell_reg[791] <= 0;					l_cell_reg[792] <= 0;					l_cell_reg[793] <= 0;					l_cell_reg[794] <= 0;					l_cell_reg[795] <= 0;					l_cell_reg[796] <= 0;					l_cell_reg[797] <= 0;					l_cell_reg[798] <= 0;					l_cell_reg[799] <= 0;					l_cell_reg[800] <= 0;					l_cell_reg[801] <= 0;					l_cell_reg[802] <= 0;					l_cell_reg[803] <= 0;					l_cell_reg[804] <= 0;					l_cell_reg[805] <= 0;					l_cell_reg[806] <= 0;					l_cell_reg[807] <= 0;					l_cell_reg[808] <= 0;					l_cell_reg[809] <= 0;					l_cell_reg[810] <= 0;					l_cell_reg[811] <= 0;					l_cell_reg[812] <= 0;					l_cell_reg[813] <= 0;					l_cell_reg[814] <= 0;					l_cell_reg[815] <= 0;					l_cell_reg[816] <= 0;					l_cell_reg[817] <= 0;					l_cell_reg[818] <= 0;					l_cell_reg[819] <= 0;					l_cell_reg[820] <= 0;					l_cell_reg[821] <= 0;					l_cell_reg[822] <= 0;					l_cell_reg[823] <= 0;					l_cell_reg[824] <= 0;					l_cell_reg[825] <= 0;					l_cell_reg[826] <= 0;					l_cell_reg[827] <= 0;					l_cell_reg[828] <= 0;					l_cell_reg[829] <= 0;					l_cell_reg[830] <= 0;					l_cell_reg[831] <= 0;					l_cell_reg[832] <= 0;					l_cell_reg[833] <= 0;					l_cell_reg[834] <= 0;					l_cell_reg[835] <= 0;					l_cell_reg[836] <= 0;					l_cell_reg[837] <= 0;					l_cell_reg[838] <= 0;					l_cell_reg[839] <= 0;					l_cell_reg[840] <= 0;					l_cell_reg[841] <= 0;					l_cell_reg[842] <= 0;					l_cell_reg[843] <= 0;					l_cell_reg[844] <= 0;					l_cell_reg[845] <= 0;					l_cell_reg[846] <= 0;					l_cell_reg[847] <= 0;					l_cell_reg[848] <= 0;					l_cell_reg[849] <= 0;					l_cell_reg[850] <= 0;					l_cell_reg[851] <= 0;					l_cell_reg[852] <= 0;					l_cell_reg[853] <= 0;					l_cell_reg[854] <= 0;					l_cell_reg[855] <= 0;					l_cell_reg[856] <= 0;					l_cell_reg[857] <= 0;					l_cell_reg[858] <= 0;					l_cell_reg[859] <= 0;					l_cell_reg[860] <= 0;					l_cell_reg[861] <= 0;					l_cell_reg[862] <= 0;					l_cell_reg[863] <= 0;					l_cell_reg[864] <= 0;					l_cell_reg[865] <= 0;					l_cell_reg[866] <= 0;					l_cell_reg[867] <= 0;					l_cell_reg[868] <= 0;					l_cell_reg[869] <= 0;					l_cell_reg[870] <= 0;					l_cell_reg[871] <= 0;					l_cell_reg[872] <= 0;					l_cell_reg[873] <= 0;					l_cell_reg[874] <= 0;					l_cell_reg[875] <= 0;					l_cell_reg[876] <= 0;					l_cell_reg[877] <= 0;					l_cell_reg[878] <= 0;					l_cell_reg[879] <= 0;					l_cell_reg[880] <= 0;					l_cell_reg[881] <= 0;					l_cell_reg[882] <= 0;					l_cell_reg[883] <= 0;					l_cell_reg[884] <= 0;					l_cell_reg[885] <= 0;					l_cell_reg[886] <= 0;					l_cell_reg[887] <= 0;					l_cell_reg[888] <= 0;					l_cell_reg[889] <= 0;					l_cell_reg[890] <= 0;					l_cell_reg[891] <= 0;					l_cell_reg[892] <= 0;					l_cell_reg[893] <= 0;					l_cell_reg[894] <= 0;					l_cell_reg[895] <= 0;					l_cell_reg[896] <= 0;					l_cell_reg[897] <= 0;					l_cell_reg[898] <= 0;					l_cell_reg[899] <= 0;					l_cell_reg[900] <= 0;					l_cell_reg[901] <= 0;					l_cell_reg[902] <= 0;					l_cell_reg[903] <= 0;					l_cell_reg[904] <= 0;					l_cell_reg[905] <= 0;					l_cell_reg[906] <= 0;					l_cell_reg[907] <= 0;					l_cell_reg[908] <= 0;					l_cell_reg[909] <= 0;					l_cell_reg[910] <= 0;					l_cell_reg[911] <= 0;					l_cell_reg[912] <= 0;					l_cell_reg[913] <= 0;					l_cell_reg[914] <= 0;					l_cell_reg[915] <= 0;					l_cell_reg[916] <= 0;					l_cell_reg[917] <= 0;					l_cell_reg[918] <= 0;					l_cell_reg[919] <= 0;					l_cell_reg[920] <= 0;					l_cell_reg[921] <= 0;					l_cell_reg[922] <= 0;					l_cell_reg[923] <= 0;					l_cell_reg[924] <= 0;					l_cell_reg[925] <= 0;					l_cell_reg[926] <= 0;					l_cell_reg[927] <= 0;					l_cell_reg[928] <= 0;					l_cell_reg[929] <= 0;					l_cell_reg[930] <= 0;					l_cell_reg[931] <= 0;					l_cell_reg[932] <= 0;					l_cell_reg[933] <= 0;					l_cell_reg[934] <= 0;					l_cell_reg[935] <= 0;					l_cell_reg[936] <= 0;					l_cell_reg[937] <= 0;					l_cell_reg[938] <= 0;					l_cell_reg[939] <= 0;					l_cell_reg[940] <= 0;					l_cell_reg[941] <= 0;					l_cell_reg[942] <= 0;					l_cell_reg[943] <= 0;					l_cell_reg[944] <= 0;					l_cell_reg[945] <= 0;					l_cell_reg[946] <= 0;					l_cell_reg[947] <= 0;					l_cell_reg[948] <= 0;					l_cell_reg[949] <= 0;					l_cell_reg[950] <= 0;					l_cell_reg[951] <= 0;					l_cell_reg[952] <= 0;					l_cell_reg[953] <= 0;					l_cell_reg[954] <= 0;					l_cell_reg[955] <= 0;					l_cell_reg[956] <= 0;					l_cell_reg[957] <= 0;					l_cell_reg[958] <= 0;					l_cell_reg[959] <= 0;					l_cell_reg[960] <= 0;					l_cell_reg[961] <= 0;					l_cell_reg[962] <= 0;					l_cell_reg[963] <= 0;					l_cell_reg[964] <= 0;					l_cell_reg[965] <= 0;					l_cell_reg[966] <= 0;					l_cell_reg[967] <= 0;					l_cell_reg[968] <= 0;					l_cell_reg[969] <= 0;					l_cell_reg[970] <= 0;					l_cell_reg[971] <= 0;					l_cell_reg[972] <= 0;					l_cell_reg[973] <= 0;					l_cell_reg[974] <= 0;					l_cell_reg[975] <= 0;					l_cell_reg[976] <= 0;					l_cell_reg[977] <= 0;					l_cell_reg[978] <= 0;					l_cell_reg[979] <= 0;					l_cell_reg[980] <= 0;					l_cell_reg[981] <= 0;					l_cell_reg[982] <= 0;					l_cell_reg[983] <= 0;					l_cell_reg[984] <= 0;					l_cell_reg[985] <= 0;					l_cell_reg[986] <= 0;					l_cell_reg[987] <= 0;					l_cell_reg[988] <= 0;					l_cell_reg[989] <= 0;					l_cell_reg[990] <= 0;					l_cell_reg[991] <= 0;					l_cell_reg[992] <= 0;					l_cell_reg[993] <= 0;					l_cell_reg[994] <= 0;					l_cell_reg[995] <= 0;					l_cell_reg[996] <= 0;					l_cell_reg[997] <= 0;					l_cell_reg[998] <= 0;					l_cell_reg[999] <= 0;					l_cell_reg[1000] <= 0;					l_cell_reg[1001] <= 0;					l_cell_reg[1002] <= 0;					l_cell_reg[1003] <= 0;					l_cell_reg[1004] <= 0;					l_cell_reg[1005] <= 0;					l_cell_reg[1006] <= 0;					l_cell_reg[1007] <= 0;					l_cell_reg[1008] <= 0;					l_cell_reg[1009] <= 0;					l_cell_reg[1010] <= 0;					l_cell_reg[1011] <= 0;					l_cell_reg[1012] <= 0;					l_cell_reg[1013] <= 0;					l_cell_reg[1014] <= 0;					l_cell_reg[1015] <= 0;					l_cell_reg[1016] <= 0;					l_cell_reg[1017] <= 0;					l_cell_reg[1018] <= 0;					l_cell_reg[1019] <= 0;					l_cell_reg[1020] <= 0;					l_cell_reg[1021] <= 0;					l_cell_reg[1022] <= 0;					l_cell_reg[1023] <= 0;			end
		endcase	end
	genvar i;	generate		for (i = 0; i < 1024 ; i = i+2)			begin :bp_2				bp_2_cell fun(					.clk(clk),					.en(1),					.R_IN1(r_cell_reg[i]),					.R_IN2(r_cell_reg[i+1]),					.L_IN1(l_cell_reg[i]),					.L_IN2(l_cell_reg[i+1]),					.R_OUT1(r_cell_wire[i]),					.R_OUT2(r_cell_wire[i+1]),					.L_OUT1(l_cell_wire[i]),					.L_OUT2(l_cell_wire[i+1])				);			end	endgenerate
	always @(posedge clk) begin		if (bp_over_flag) begin			OUT_1 <= inform_L [0][0] ;			OUT_2 <= inform_L [1][0] ;			OUT_3 <= inform_L [2][0] ;			OUT_4 <= inform_L [3][0] ;			OUT_5 <= inform_L [4][0] ;			OUT_6 <= inform_L [5][0] ;			OUT_7 <= inform_L [6][0] ;			OUT_8 <= inform_L [7][0] ;			OUT_9 <= inform_L [8][0] ;			OUT_10 <= inform_L [9][0] ;			OUT_11 <= inform_L [10][0] ;			OUT_12 <= inform_L [11][0] ;			OUT_13 <= inform_L [12][0] ;			OUT_14 <= inform_L [13][0] ;			OUT_15 <= inform_L [14][0] ;			OUT_16 <= inform_L [15][0] ;			OUT_17 <= inform_L [16][0] ;			OUT_18 <= inform_L [17][0] ;			OUT_19 <= inform_L [18][0] ;			OUT_20 <= inform_L [19][0] ;			OUT_21 <= inform_L [20][0] ;			OUT_22 <= inform_L [21][0] ;			OUT_23 <= inform_L [22][0] ;			OUT_24 <= inform_L [23][0] ;			OUT_25 <= inform_L [24][0] ;			OUT_26 <= inform_L [25][0] ;			OUT_27 <= inform_L [26][0] ;			OUT_28 <= inform_L [27][0] ;			OUT_29 <= inform_L [28][0] ;			OUT_30 <= inform_L [29][0] ;			OUT_31 <= inform_L [30][0] ;			OUT_32 <= inform_L [31][0] ;			OUT_33 <= inform_L [32][0] ;			OUT_34 <= inform_L [33][0] ;			OUT_35 <= inform_L [34][0] ;			OUT_36 <= inform_L [35][0] ;			OUT_37 <= inform_L [36][0] ;			OUT_38 <= inform_L [37][0] ;			OUT_39 <= inform_L [38][0] ;			OUT_40 <= inform_L [39][0] ;			OUT_41 <= inform_L [40][0] ;			OUT_42 <= inform_L [41][0] ;			OUT_43 <= inform_L [42][0] ;			OUT_44 <= inform_L [43][0] ;			OUT_45 <= inform_L [44][0] ;			OUT_46 <= inform_L [45][0] ;			OUT_47 <= inform_L [46][0] ;			OUT_48 <= inform_L [47][0] ;			OUT_49 <= inform_L [48][0] ;			OUT_50 <= inform_L [49][0] ;			OUT_51 <= inform_L [50][0] ;			OUT_52 <= inform_L [51][0] ;			OUT_53 <= inform_L [52][0] ;			OUT_54 <= inform_L [53][0] ;			OUT_55 <= inform_L [54][0] ;			OUT_56 <= inform_L [55][0] ;			OUT_57 <= inform_L [56][0] ;			OUT_58 <= inform_L [57][0] ;			OUT_59 <= inform_L [58][0] ;			OUT_60 <= inform_L [59][0] ;			OUT_61 <= inform_L [60][0] ;			OUT_62 <= inform_L [61][0] ;			OUT_63 <= inform_L [62][0] ;			OUT_64 <= inform_L [63][0] ;			OUT_65 <= inform_L [64][0] ;			OUT_66 <= inform_L [65][0] ;			OUT_67 <= inform_L [66][0] ;			OUT_68 <= inform_L [67][0] ;			OUT_69 <= inform_L [68][0] ;			OUT_70 <= inform_L [69][0] ;			OUT_71 <= inform_L [70][0] ;			OUT_72 <= inform_L [71][0] ;			OUT_73 <= inform_L [72][0] ;			OUT_74 <= inform_L [73][0] ;			OUT_75 <= inform_L [74][0] ;			OUT_76 <= inform_L [75][0] ;			OUT_77 <= inform_L [76][0] ;			OUT_78 <= inform_L [77][0] ;			OUT_79 <= inform_L [78][0] ;			OUT_80 <= inform_L [79][0] ;			OUT_81 <= inform_L [80][0] ;			OUT_82 <= inform_L [81][0] ;			OUT_83 <= inform_L [82][0] ;			OUT_84 <= inform_L [83][0] ;			OUT_85 <= inform_L [84][0] ;			OUT_86 <= inform_L [85][0] ;			OUT_87 <= inform_L [86][0] ;			OUT_88 <= inform_L [87][0] ;			OUT_89 <= inform_L [88][0] ;			OUT_90 <= inform_L [89][0] ;			OUT_91 <= inform_L [90][0] ;			OUT_92 <= inform_L [91][0] ;			OUT_93 <= inform_L [92][0] ;			OUT_94 <= inform_L [93][0] ;			OUT_95 <= inform_L [94][0] ;			OUT_96 <= inform_L [95][0] ;			OUT_97 <= inform_L [96][0] ;			OUT_98 <= inform_L [97][0] ;			OUT_99 <= inform_L [98][0] ;			OUT_100 <= inform_L [99][0] ;			OUT_101 <= inform_L [100][0] ;			OUT_102 <= inform_L [101][0] ;			OUT_103 <= inform_L [102][0] ;			OUT_104 <= inform_L [103][0] ;			OUT_105 <= inform_L [104][0] ;			OUT_106 <= inform_L [105][0] ;			OUT_107 <= inform_L [106][0] ;			OUT_108 <= inform_L [107][0] ;			OUT_109 <= inform_L [108][0] ;			OUT_110 <= inform_L [109][0] ;			OUT_111 <= inform_L [110][0] ;			OUT_112 <= inform_L [111][0] ;			OUT_113 <= inform_L [112][0] ;			OUT_114 <= inform_L [113][0] ;			OUT_115 <= inform_L [114][0] ;			OUT_116 <= inform_L [115][0] ;			OUT_117 <= inform_L [116][0] ;			OUT_118 <= inform_L [117][0] ;			OUT_119 <= inform_L [118][0] ;			OUT_120 <= inform_L [119][0] ;			OUT_121 <= inform_L [120][0] ;			OUT_122 <= inform_L [121][0] ;			OUT_123 <= inform_L [122][0] ;			OUT_124 <= inform_L [123][0] ;			OUT_125 <= inform_L [124][0] ;			OUT_126 <= inform_L [125][0] ;			OUT_127 <= inform_L [126][0] ;			OUT_128 <= inform_L [127][0] ;			OUT_129 <= inform_L [128][0] ;			OUT_130 <= inform_L [129][0] ;			OUT_131 <= inform_L [130][0] ;			OUT_132 <= inform_L [131][0] ;			OUT_133 <= inform_L [132][0] ;			OUT_134 <= inform_L [133][0] ;			OUT_135 <= inform_L [134][0] ;			OUT_136 <= inform_L [135][0] ;			OUT_137 <= inform_L [136][0] ;			OUT_138 <= inform_L [137][0] ;			OUT_139 <= inform_L [138][0] ;			OUT_140 <= inform_L [139][0] ;			OUT_141 <= inform_L [140][0] ;			OUT_142 <= inform_L [141][0] ;			OUT_143 <= inform_L [142][0] ;			OUT_144 <= inform_L [143][0] ;			OUT_145 <= inform_L [144][0] ;			OUT_146 <= inform_L [145][0] ;			OUT_147 <= inform_L [146][0] ;			OUT_148 <= inform_L [147][0] ;			OUT_149 <= inform_L [148][0] ;			OUT_150 <= inform_L [149][0] ;			OUT_151 <= inform_L [150][0] ;			OUT_152 <= inform_L [151][0] ;			OUT_153 <= inform_L [152][0] ;			OUT_154 <= inform_L [153][0] ;			OUT_155 <= inform_L [154][0] ;			OUT_156 <= inform_L [155][0] ;			OUT_157 <= inform_L [156][0] ;			OUT_158 <= inform_L [157][0] ;			OUT_159 <= inform_L [158][0] ;			OUT_160 <= inform_L [159][0] ;			OUT_161 <= inform_L [160][0] ;			OUT_162 <= inform_L [161][0] ;			OUT_163 <= inform_L [162][0] ;			OUT_164 <= inform_L [163][0] ;			OUT_165 <= inform_L [164][0] ;			OUT_166 <= inform_L [165][0] ;			OUT_167 <= inform_L [166][0] ;			OUT_168 <= inform_L [167][0] ;			OUT_169 <= inform_L [168][0] ;			OUT_170 <= inform_L [169][0] ;			OUT_171 <= inform_L [170][0] ;			OUT_172 <= inform_L [171][0] ;			OUT_173 <= inform_L [172][0] ;			OUT_174 <= inform_L [173][0] ;			OUT_175 <= inform_L [174][0] ;			OUT_176 <= inform_L [175][0] ;			OUT_177 <= inform_L [176][0] ;			OUT_178 <= inform_L [177][0] ;			OUT_179 <= inform_L [178][0] ;			OUT_180 <= inform_L [179][0] ;			OUT_181 <= inform_L [180][0] ;			OUT_182 <= inform_L [181][0] ;			OUT_183 <= inform_L [182][0] ;			OUT_184 <= inform_L [183][0] ;			OUT_185 <= inform_L [184][0] ;			OUT_186 <= inform_L [185][0] ;			OUT_187 <= inform_L [186][0] ;			OUT_188 <= inform_L [187][0] ;			OUT_189 <= inform_L [188][0] ;			OUT_190 <= inform_L [189][0] ;			OUT_191 <= inform_L [190][0] ;			OUT_192 <= inform_L [191][0] ;			OUT_193 <= inform_L [192][0] ;			OUT_194 <= inform_L [193][0] ;			OUT_195 <= inform_L [194][0] ;			OUT_196 <= inform_L [195][0] ;			OUT_197 <= inform_L [196][0] ;			OUT_198 <= inform_L [197][0] ;			OUT_199 <= inform_L [198][0] ;			OUT_200 <= inform_L [199][0] ;			OUT_201 <= inform_L [200][0] ;			OUT_202 <= inform_L [201][0] ;			OUT_203 <= inform_L [202][0] ;			OUT_204 <= inform_L [203][0] ;			OUT_205 <= inform_L [204][0] ;			OUT_206 <= inform_L [205][0] ;			OUT_207 <= inform_L [206][0] ;			OUT_208 <= inform_L [207][0] ;			OUT_209 <= inform_L [208][0] ;			OUT_210 <= inform_L [209][0] ;			OUT_211 <= inform_L [210][0] ;			OUT_212 <= inform_L [211][0] ;			OUT_213 <= inform_L [212][0] ;			OUT_214 <= inform_L [213][0] ;			OUT_215 <= inform_L [214][0] ;			OUT_216 <= inform_L [215][0] ;			OUT_217 <= inform_L [216][0] ;			OUT_218 <= inform_L [217][0] ;			OUT_219 <= inform_L [218][0] ;			OUT_220 <= inform_L [219][0] ;			OUT_221 <= inform_L [220][0] ;			OUT_222 <= inform_L [221][0] ;			OUT_223 <= inform_L [222][0] ;			OUT_224 <= inform_L [223][0] ;			OUT_225 <= inform_L [224][0] ;			OUT_226 <= inform_L [225][0] ;			OUT_227 <= inform_L [226][0] ;			OUT_228 <= inform_L [227][0] ;			OUT_229 <= inform_L [228][0] ;			OUT_230 <= inform_L [229][0] ;			OUT_231 <= inform_L [230][0] ;			OUT_232 <= inform_L [231][0] ;			OUT_233 <= inform_L [232][0] ;			OUT_234 <= inform_L [233][0] ;			OUT_235 <= inform_L [234][0] ;			OUT_236 <= inform_L [235][0] ;			OUT_237 <= inform_L [236][0] ;			OUT_238 <= inform_L [237][0] ;			OUT_239 <= inform_L [238][0] ;			OUT_240 <= inform_L [239][0] ;			OUT_241 <= inform_L [240][0] ;			OUT_242 <= inform_L [241][0] ;			OUT_243 <= inform_L [242][0] ;			OUT_244 <= inform_L [243][0] ;			OUT_245 <= inform_L [244][0] ;			OUT_246 <= inform_L [245][0] ;			OUT_247 <= inform_L [246][0] ;			OUT_248 <= inform_L [247][0] ;			OUT_249 <= inform_L [248][0] ;			OUT_250 <= inform_L [249][0] ;			OUT_251 <= inform_L [250][0] ;			OUT_252 <= inform_L [251][0] ;			OUT_253 <= inform_L [252][0] ;			OUT_254 <= inform_L [253][0] ;			OUT_255 <= inform_L [254][0] ;			OUT_256 <= inform_L [255][0] ;			OUT_257 <= inform_L [256][0] ;			OUT_258 <= inform_L [257][0] ;			OUT_259 <= inform_L [258][0] ;			OUT_260 <= inform_L [259][0] ;			OUT_261 <= inform_L [260][0] ;			OUT_262 <= inform_L [261][0] ;			OUT_263 <= inform_L [262][0] ;			OUT_264 <= inform_L [263][0] ;			OUT_265 <= inform_L [264][0] ;			OUT_266 <= inform_L [265][0] ;			OUT_267 <= inform_L [266][0] ;			OUT_268 <= inform_L [267][0] ;			OUT_269 <= inform_L [268][0] ;			OUT_270 <= inform_L [269][0] ;			OUT_271 <= inform_L [270][0] ;			OUT_272 <= inform_L [271][0] ;			OUT_273 <= inform_L [272][0] ;			OUT_274 <= inform_L [273][0] ;			OUT_275 <= inform_L [274][0] ;			OUT_276 <= inform_L [275][0] ;			OUT_277 <= inform_L [276][0] ;			OUT_278 <= inform_L [277][0] ;			OUT_279 <= inform_L [278][0] ;			OUT_280 <= inform_L [279][0] ;			OUT_281 <= inform_L [280][0] ;			OUT_282 <= inform_L [281][0] ;			OUT_283 <= inform_L [282][0] ;			OUT_284 <= inform_L [283][0] ;			OUT_285 <= inform_L [284][0] ;			OUT_286 <= inform_L [285][0] ;			OUT_287 <= inform_L [286][0] ;			OUT_288 <= inform_L [287][0] ;			OUT_289 <= inform_L [288][0] ;			OUT_290 <= inform_L [289][0] ;			OUT_291 <= inform_L [290][0] ;			OUT_292 <= inform_L [291][0] ;			OUT_293 <= inform_L [292][0] ;			OUT_294 <= inform_L [293][0] ;			OUT_295 <= inform_L [294][0] ;			OUT_296 <= inform_L [295][0] ;			OUT_297 <= inform_L [296][0] ;			OUT_298 <= inform_L [297][0] ;			OUT_299 <= inform_L [298][0] ;			OUT_300 <= inform_L [299][0] ;			OUT_301 <= inform_L [300][0] ;			OUT_302 <= inform_L [301][0] ;			OUT_303 <= inform_L [302][0] ;			OUT_304 <= inform_L [303][0] ;			OUT_305 <= inform_L [304][0] ;			OUT_306 <= inform_L [305][0] ;			OUT_307 <= inform_L [306][0] ;			OUT_308 <= inform_L [307][0] ;			OUT_309 <= inform_L [308][0] ;			OUT_310 <= inform_L [309][0] ;			OUT_311 <= inform_L [310][0] ;			OUT_312 <= inform_L [311][0] ;			OUT_313 <= inform_L [312][0] ;			OUT_314 <= inform_L [313][0] ;			OUT_315 <= inform_L [314][0] ;			OUT_316 <= inform_L [315][0] ;			OUT_317 <= inform_L [316][0] ;			OUT_318 <= inform_L [317][0] ;			OUT_319 <= inform_L [318][0] ;			OUT_320 <= inform_L [319][0] ;			OUT_321 <= inform_L [320][0] ;			OUT_322 <= inform_L [321][0] ;			OUT_323 <= inform_L [322][0] ;			OUT_324 <= inform_L [323][0] ;			OUT_325 <= inform_L [324][0] ;			OUT_326 <= inform_L [325][0] ;			OUT_327 <= inform_L [326][0] ;			OUT_328 <= inform_L [327][0] ;			OUT_329 <= inform_L [328][0] ;			OUT_330 <= inform_L [329][0] ;			OUT_331 <= inform_L [330][0] ;			OUT_332 <= inform_L [331][0] ;			OUT_333 <= inform_L [332][0] ;			OUT_334 <= inform_L [333][0] ;			OUT_335 <= inform_L [334][0] ;			OUT_336 <= inform_L [335][0] ;			OUT_337 <= inform_L [336][0] ;			OUT_338 <= inform_L [337][0] ;			OUT_339 <= inform_L [338][0] ;			OUT_340 <= inform_L [339][0] ;			OUT_341 <= inform_L [340][0] ;			OUT_342 <= inform_L [341][0] ;			OUT_343 <= inform_L [342][0] ;			OUT_344 <= inform_L [343][0] ;			OUT_345 <= inform_L [344][0] ;			OUT_346 <= inform_L [345][0] ;			OUT_347 <= inform_L [346][0] ;			OUT_348 <= inform_L [347][0] ;			OUT_349 <= inform_L [348][0] ;			OUT_350 <= inform_L [349][0] ;			OUT_351 <= inform_L [350][0] ;			OUT_352 <= inform_L [351][0] ;			OUT_353 <= inform_L [352][0] ;			OUT_354 <= inform_L [353][0] ;			OUT_355 <= inform_L [354][0] ;			OUT_356 <= inform_L [355][0] ;			OUT_357 <= inform_L [356][0] ;			OUT_358 <= inform_L [357][0] ;			OUT_359 <= inform_L [358][0] ;			OUT_360 <= inform_L [359][0] ;			OUT_361 <= inform_L [360][0] ;			OUT_362 <= inform_L [361][0] ;			OUT_363 <= inform_L [362][0] ;			OUT_364 <= inform_L [363][0] ;			OUT_365 <= inform_L [364][0] ;			OUT_366 <= inform_L [365][0] ;			OUT_367 <= inform_L [366][0] ;			OUT_368 <= inform_L [367][0] ;			OUT_369 <= inform_L [368][0] ;			OUT_370 <= inform_L [369][0] ;			OUT_371 <= inform_L [370][0] ;			OUT_372 <= inform_L [371][0] ;			OUT_373 <= inform_L [372][0] ;			OUT_374 <= inform_L [373][0] ;			OUT_375 <= inform_L [374][0] ;			OUT_376 <= inform_L [375][0] ;			OUT_377 <= inform_L [376][0] ;			OUT_378 <= inform_L [377][0] ;			OUT_379 <= inform_L [378][0] ;			OUT_380 <= inform_L [379][0] ;			OUT_381 <= inform_L [380][0] ;			OUT_382 <= inform_L [381][0] ;			OUT_383 <= inform_L [382][0] ;			OUT_384 <= inform_L [383][0] ;			OUT_385 <= inform_L [384][0] ;			OUT_386 <= inform_L [385][0] ;			OUT_387 <= inform_L [386][0] ;			OUT_388 <= inform_L [387][0] ;			OUT_389 <= inform_L [388][0] ;			OUT_390 <= inform_L [389][0] ;			OUT_391 <= inform_L [390][0] ;			OUT_392 <= inform_L [391][0] ;			OUT_393 <= inform_L [392][0] ;			OUT_394 <= inform_L [393][0] ;			OUT_395 <= inform_L [394][0] ;			OUT_396 <= inform_L [395][0] ;			OUT_397 <= inform_L [396][0] ;			OUT_398 <= inform_L [397][0] ;			OUT_399 <= inform_L [398][0] ;			OUT_400 <= inform_L [399][0] ;			OUT_401 <= inform_L [400][0] ;			OUT_402 <= inform_L [401][0] ;			OUT_403 <= inform_L [402][0] ;			OUT_404 <= inform_L [403][0] ;			OUT_405 <= inform_L [404][0] ;			OUT_406 <= inform_L [405][0] ;			OUT_407 <= inform_L [406][0] ;			OUT_408 <= inform_L [407][0] ;			OUT_409 <= inform_L [408][0] ;			OUT_410 <= inform_L [409][0] ;			OUT_411 <= inform_L [410][0] ;			OUT_412 <= inform_L [411][0] ;			OUT_413 <= inform_L [412][0] ;			OUT_414 <= inform_L [413][0] ;			OUT_415 <= inform_L [414][0] ;			OUT_416 <= inform_L [415][0] ;			OUT_417 <= inform_L [416][0] ;			OUT_418 <= inform_L [417][0] ;			OUT_419 <= inform_L [418][0] ;			OUT_420 <= inform_L [419][0] ;			OUT_421 <= inform_L [420][0] ;			OUT_422 <= inform_L [421][0] ;			OUT_423 <= inform_L [422][0] ;			OUT_424 <= inform_L [423][0] ;			OUT_425 <= inform_L [424][0] ;			OUT_426 <= inform_L [425][0] ;			OUT_427 <= inform_L [426][0] ;			OUT_428 <= inform_L [427][0] ;			OUT_429 <= inform_L [428][0] ;			OUT_430 <= inform_L [429][0] ;			OUT_431 <= inform_L [430][0] ;			OUT_432 <= inform_L [431][0] ;			OUT_433 <= inform_L [432][0] ;			OUT_434 <= inform_L [433][0] ;			OUT_435 <= inform_L [434][0] ;			OUT_436 <= inform_L [435][0] ;			OUT_437 <= inform_L [436][0] ;			OUT_438 <= inform_L [437][0] ;			OUT_439 <= inform_L [438][0] ;			OUT_440 <= inform_L [439][0] ;			OUT_441 <= inform_L [440][0] ;			OUT_442 <= inform_L [441][0] ;			OUT_443 <= inform_L [442][0] ;			OUT_444 <= inform_L [443][0] ;			OUT_445 <= inform_L [444][0] ;			OUT_446 <= inform_L [445][0] ;			OUT_447 <= inform_L [446][0] ;			OUT_448 <= inform_L [447][0] ;			OUT_449 <= inform_L [448][0] ;			OUT_450 <= inform_L [449][0] ;			OUT_451 <= inform_L [450][0] ;			OUT_452 <= inform_L [451][0] ;			OUT_453 <= inform_L [452][0] ;			OUT_454 <= inform_L [453][0] ;			OUT_455 <= inform_L [454][0] ;			OUT_456 <= inform_L [455][0] ;			OUT_457 <= inform_L [456][0] ;			OUT_458 <= inform_L [457][0] ;			OUT_459 <= inform_L [458][0] ;			OUT_460 <= inform_L [459][0] ;			OUT_461 <= inform_L [460][0] ;			OUT_462 <= inform_L [461][0] ;			OUT_463 <= inform_L [462][0] ;			OUT_464 <= inform_L [463][0] ;			OUT_465 <= inform_L [464][0] ;			OUT_466 <= inform_L [465][0] ;			OUT_467 <= inform_L [466][0] ;			OUT_468 <= inform_L [467][0] ;			OUT_469 <= inform_L [468][0] ;			OUT_470 <= inform_L [469][0] ;			OUT_471 <= inform_L [470][0] ;			OUT_472 <= inform_L [471][0] ;			OUT_473 <= inform_L [472][0] ;			OUT_474 <= inform_L [473][0] ;			OUT_475 <= inform_L [474][0] ;			OUT_476 <= inform_L [475][0] ;			OUT_477 <= inform_L [476][0] ;			OUT_478 <= inform_L [477][0] ;			OUT_479 <= inform_L [478][0] ;			OUT_480 <= inform_L [479][0] ;			OUT_481 <= inform_L [480][0] ;			OUT_482 <= inform_L [481][0] ;			OUT_483 <= inform_L [482][0] ;			OUT_484 <= inform_L [483][0] ;			OUT_485 <= inform_L [484][0] ;			OUT_486 <= inform_L [485][0] ;			OUT_487 <= inform_L [486][0] ;			OUT_488 <= inform_L [487][0] ;			OUT_489 <= inform_L [488][0] ;			OUT_490 <= inform_L [489][0] ;			OUT_491 <= inform_L [490][0] ;			OUT_492 <= inform_L [491][0] ;			OUT_493 <= inform_L [492][0] ;			OUT_494 <= inform_L [493][0] ;			OUT_495 <= inform_L [494][0] ;			OUT_496 <= inform_L [495][0] ;			OUT_497 <= inform_L [496][0] ;			OUT_498 <= inform_L [497][0] ;			OUT_499 <= inform_L [498][0] ;			OUT_500 <= inform_L [499][0] ;			OUT_501 <= inform_L [500][0] ;			OUT_502 <= inform_L [501][0] ;			OUT_503 <= inform_L [502][0] ;			OUT_504 <= inform_L [503][0] ;			OUT_505 <= inform_L [504][0] ;			OUT_506 <= inform_L [505][0] ;			OUT_507 <= inform_L [506][0] ;			OUT_508 <= inform_L [507][0] ;			OUT_509 <= inform_L [508][0] ;			OUT_510 <= inform_L [509][0] ;			OUT_511 <= inform_L [510][0] ;			OUT_512 <= inform_L [511][0] ;			OUT_513 <= inform_L [512][0] ;			OUT_514 <= inform_L [513][0] ;			OUT_515 <= inform_L [514][0] ;			OUT_516 <= inform_L [515][0] ;			OUT_517 <= inform_L [516][0] ;			OUT_518 <= inform_L [517][0] ;			OUT_519 <= inform_L [518][0] ;			OUT_520 <= inform_L [519][0] ;			OUT_521 <= inform_L [520][0] ;			OUT_522 <= inform_L [521][0] ;			OUT_523 <= inform_L [522][0] ;			OUT_524 <= inform_L [523][0] ;			OUT_525 <= inform_L [524][0] ;			OUT_526 <= inform_L [525][0] ;			OUT_527 <= inform_L [526][0] ;			OUT_528 <= inform_L [527][0] ;			OUT_529 <= inform_L [528][0] ;			OUT_530 <= inform_L [529][0] ;			OUT_531 <= inform_L [530][0] ;			OUT_532 <= inform_L [531][0] ;			OUT_533 <= inform_L [532][0] ;			OUT_534 <= inform_L [533][0] ;			OUT_535 <= inform_L [534][0] ;			OUT_536 <= inform_L [535][0] ;			OUT_537 <= inform_L [536][0] ;			OUT_538 <= inform_L [537][0] ;			OUT_539 <= inform_L [538][0] ;			OUT_540 <= inform_L [539][0] ;			OUT_541 <= inform_L [540][0] ;			OUT_542 <= inform_L [541][0] ;			OUT_543 <= inform_L [542][0] ;			OUT_544 <= inform_L [543][0] ;			OUT_545 <= inform_L [544][0] ;			OUT_546 <= inform_L [545][0] ;			OUT_547 <= inform_L [546][0] ;			OUT_548 <= inform_L [547][0] ;			OUT_549 <= inform_L [548][0] ;			OUT_550 <= inform_L [549][0] ;			OUT_551 <= inform_L [550][0] ;			OUT_552 <= inform_L [551][0] ;			OUT_553 <= inform_L [552][0] ;			OUT_554 <= inform_L [553][0] ;			OUT_555 <= inform_L [554][0] ;			OUT_556 <= inform_L [555][0] ;			OUT_557 <= inform_L [556][0] ;			OUT_558 <= inform_L [557][0] ;			OUT_559 <= inform_L [558][0] ;			OUT_560 <= inform_L [559][0] ;			OUT_561 <= inform_L [560][0] ;			OUT_562 <= inform_L [561][0] ;			OUT_563 <= inform_L [562][0] ;			OUT_564 <= inform_L [563][0] ;			OUT_565 <= inform_L [564][0] ;			OUT_566 <= inform_L [565][0] ;			OUT_567 <= inform_L [566][0] ;			OUT_568 <= inform_L [567][0] ;			OUT_569 <= inform_L [568][0] ;			OUT_570 <= inform_L [569][0] ;			OUT_571 <= inform_L [570][0] ;			OUT_572 <= inform_L [571][0] ;			OUT_573 <= inform_L [572][0] ;			OUT_574 <= inform_L [573][0] ;			OUT_575 <= inform_L [574][0] ;			OUT_576 <= inform_L [575][0] ;			OUT_577 <= inform_L [576][0] ;			OUT_578 <= inform_L [577][0] ;			OUT_579 <= inform_L [578][0] ;			OUT_580 <= inform_L [579][0] ;			OUT_581 <= inform_L [580][0] ;			OUT_582 <= inform_L [581][0] ;			OUT_583 <= inform_L [582][0] ;			OUT_584 <= inform_L [583][0] ;			OUT_585 <= inform_L [584][0] ;			OUT_586 <= inform_L [585][0] ;			OUT_587 <= inform_L [586][0] ;			OUT_588 <= inform_L [587][0] ;			OUT_589 <= inform_L [588][0] ;			OUT_590 <= inform_L [589][0] ;			OUT_591 <= inform_L [590][0] ;			OUT_592 <= inform_L [591][0] ;			OUT_593 <= inform_L [592][0] ;			OUT_594 <= inform_L [593][0] ;			OUT_595 <= inform_L [594][0] ;			OUT_596 <= inform_L [595][0] ;			OUT_597 <= inform_L [596][0] ;			OUT_598 <= inform_L [597][0] ;			OUT_599 <= inform_L [598][0] ;			OUT_600 <= inform_L [599][0] ;			OUT_601 <= inform_L [600][0] ;			OUT_602 <= inform_L [601][0] ;			OUT_603 <= inform_L [602][0] ;			OUT_604 <= inform_L [603][0] ;			OUT_605 <= inform_L [604][0] ;			OUT_606 <= inform_L [605][0] ;			OUT_607 <= inform_L [606][0] ;			OUT_608 <= inform_L [607][0] ;			OUT_609 <= inform_L [608][0] ;			OUT_610 <= inform_L [609][0] ;			OUT_611 <= inform_L [610][0] ;			OUT_612 <= inform_L [611][0] ;			OUT_613 <= inform_L [612][0] ;			OUT_614 <= inform_L [613][0] ;			OUT_615 <= inform_L [614][0] ;			OUT_616 <= inform_L [615][0] ;			OUT_617 <= inform_L [616][0] ;			OUT_618 <= inform_L [617][0] ;			OUT_619 <= inform_L [618][0] ;			OUT_620 <= inform_L [619][0] ;			OUT_621 <= inform_L [620][0] ;			OUT_622 <= inform_L [621][0] ;			OUT_623 <= inform_L [622][0] ;			OUT_624 <= inform_L [623][0] ;			OUT_625 <= inform_L [624][0] ;			OUT_626 <= inform_L [625][0] ;			OUT_627 <= inform_L [626][0] ;			OUT_628 <= inform_L [627][0] ;			OUT_629 <= inform_L [628][0] ;			OUT_630 <= inform_L [629][0] ;			OUT_631 <= inform_L [630][0] ;			OUT_632 <= inform_L [631][0] ;			OUT_633 <= inform_L [632][0] ;			OUT_634 <= inform_L [633][0] ;			OUT_635 <= inform_L [634][0] ;			OUT_636 <= inform_L [635][0] ;			OUT_637 <= inform_L [636][0] ;			OUT_638 <= inform_L [637][0] ;			OUT_639 <= inform_L [638][0] ;			OUT_640 <= inform_L [639][0] ;			OUT_641 <= inform_L [640][0] ;			OUT_642 <= inform_L [641][0] ;			OUT_643 <= inform_L [642][0] ;			OUT_644 <= inform_L [643][0] ;			OUT_645 <= inform_L [644][0] ;			OUT_646 <= inform_L [645][0] ;			OUT_647 <= inform_L [646][0] ;			OUT_648 <= inform_L [647][0] ;			OUT_649 <= inform_L [648][0] ;			OUT_650 <= inform_L [649][0] ;			OUT_651 <= inform_L [650][0] ;			OUT_652 <= inform_L [651][0] ;			OUT_653 <= inform_L [652][0] ;			OUT_654 <= inform_L [653][0] ;			OUT_655 <= inform_L [654][0] ;			OUT_656 <= inform_L [655][0] ;			OUT_657 <= inform_L [656][0] ;			OUT_658 <= inform_L [657][0] ;			OUT_659 <= inform_L [658][0] ;			OUT_660 <= inform_L [659][0] ;			OUT_661 <= inform_L [660][0] ;			OUT_662 <= inform_L [661][0] ;			OUT_663 <= inform_L [662][0] ;			OUT_664 <= inform_L [663][0] ;			OUT_665 <= inform_L [664][0] ;			OUT_666 <= inform_L [665][0] ;			OUT_667 <= inform_L [666][0] ;			OUT_668 <= inform_L [667][0] ;			OUT_669 <= inform_L [668][0] ;			OUT_670 <= inform_L [669][0] ;			OUT_671 <= inform_L [670][0] ;			OUT_672 <= inform_L [671][0] ;			OUT_673 <= inform_L [672][0] ;			OUT_674 <= inform_L [673][0] ;			OUT_675 <= inform_L [674][0] ;			OUT_676 <= inform_L [675][0] ;			OUT_677 <= inform_L [676][0] ;			OUT_678 <= inform_L [677][0] ;			OUT_679 <= inform_L [678][0] ;			OUT_680 <= inform_L [679][0] ;			OUT_681 <= inform_L [680][0] ;			OUT_682 <= inform_L [681][0] ;			OUT_683 <= inform_L [682][0] ;			OUT_684 <= inform_L [683][0] ;			OUT_685 <= inform_L [684][0] ;			OUT_686 <= inform_L [685][0] ;			OUT_687 <= inform_L [686][0] ;			OUT_688 <= inform_L [687][0] ;			OUT_689 <= inform_L [688][0] ;			OUT_690 <= inform_L [689][0] ;			OUT_691 <= inform_L [690][0] ;			OUT_692 <= inform_L [691][0] ;			OUT_693 <= inform_L [692][0] ;			OUT_694 <= inform_L [693][0] ;			OUT_695 <= inform_L [694][0] ;			OUT_696 <= inform_L [695][0] ;			OUT_697 <= inform_L [696][0] ;			OUT_698 <= inform_L [697][0] ;			OUT_699 <= inform_L [698][0] ;			OUT_700 <= inform_L [699][0] ;			OUT_701 <= inform_L [700][0] ;			OUT_702 <= inform_L [701][0] ;			OUT_703 <= inform_L [702][0] ;			OUT_704 <= inform_L [703][0] ;			OUT_705 <= inform_L [704][0] ;			OUT_706 <= inform_L [705][0] ;			OUT_707 <= inform_L [706][0] ;			OUT_708 <= inform_L [707][0] ;			OUT_709 <= inform_L [708][0] ;			OUT_710 <= inform_L [709][0] ;			OUT_711 <= inform_L [710][0] ;			OUT_712 <= inform_L [711][0] ;			OUT_713 <= inform_L [712][0] ;			OUT_714 <= inform_L [713][0] ;			OUT_715 <= inform_L [714][0] ;			OUT_716 <= inform_L [715][0] ;			OUT_717 <= inform_L [716][0] ;			OUT_718 <= inform_L [717][0] ;			OUT_719 <= inform_L [718][0] ;			OUT_720 <= inform_L [719][0] ;			OUT_721 <= inform_L [720][0] ;			OUT_722 <= inform_L [721][0] ;			OUT_723 <= inform_L [722][0] ;			OUT_724 <= inform_L [723][0] ;			OUT_725 <= inform_L [724][0] ;			OUT_726 <= inform_L [725][0] ;			OUT_727 <= inform_L [726][0] ;			OUT_728 <= inform_L [727][0] ;			OUT_729 <= inform_L [728][0] ;			OUT_730 <= inform_L [729][0] ;			OUT_731 <= inform_L [730][0] ;			OUT_732 <= inform_L [731][0] ;			OUT_733 <= inform_L [732][0] ;			OUT_734 <= inform_L [733][0] ;			OUT_735 <= inform_L [734][0] ;			OUT_736 <= inform_L [735][0] ;			OUT_737 <= inform_L [736][0] ;			OUT_738 <= inform_L [737][0] ;			OUT_739 <= inform_L [738][0] ;			OUT_740 <= inform_L [739][0] ;			OUT_741 <= inform_L [740][0] ;			OUT_742 <= inform_L [741][0] ;			OUT_743 <= inform_L [742][0] ;			OUT_744 <= inform_L [743][0] ;			OUT_745 <= inform_L [744][0] ;			OUT_746 <= inform_L [745][0] ;			OUT_747 <= inform_L [746][0] ;			OUT_748 <= inform_L [747][0] ;			OUT_749 <= inform_L [748][0] ;			OUT_750 <= inform_L [749][0] ;			OUT_751 <= inform_L [750][0] ;			OUT_752 <= inform_L [751][0] ;			OUT_753 <= inform_L [752][0] ;			OUT_754 <= inform_L [753][0] ;			OUT_755 <= inform_L [754][0] ;			OUT_756 <= inform_L [755][0] ;			OUT_757 <= inform_L [756][0] ;			OUT_758 <= inform_L [757][0] ;			OUT_759 <= inform_L [758][0] ;			OUT_760 <= inform_L [759][0] ;			OUT_761 <= inform_L [760][0] ;			OUT_762 <= inform_L [761][0] ;			OUT_763 <= inform_L [762][0] ;			OUT_764 <= inform_L [763][0] ;			OUT_765 <= inform_L [764][0] ;			OUT_766 <= inform_L [765][0] ;			OUT_767 <= inform_L [766][0] ;			OUT_768 <= inform_L [767][0] ;			OUT_769 <= inform_L [768][0] ;			OUT_770 <= inform_L [769][0] ;			OUT_771 <= inform_L [770][0] ;			OUT_772 <= inform_L [771][0] ;			OUT_773 <= inform_L [772][0] ;			OUT_774 <= inform_L [773][0] ;			OUT_775 <= inform_L [774][0] ;			OUT_776 <= inform_L [775][0] ;			OUT_777 <= inform_L [776][0] ;			OUT_778 <= inform_L [777][0] ;			OUT_779 <= inform_L [778][0] ;			OUT_780 <= inform_L [779][0] ;			OUT_781 <= inform_L [780][0] ;			OUT_782 <= inform_L [781][0] ;			OUT_783 <= inform_L [782][0] ;			OUT_784 <= inform_L [783][0] ;			OUT_785 <= inform_L [784][0] ;			OUT_786 <= inform_L [785][0] ;			OUT_787 <= inform_L [786][0] ;			OUT_788 <= inform_L [787][0] ;			OUT_789 <= inform_L [788][0] ;			OUT_790 <= inform_L [789][0] ;			OUT_791 <= inform_L [790][0] ;			OUT_792 <= inform_L [791][0] ;			OUT_793 <= inform_L [792][0] ;			OUT_794 <= inform_L [793][0] ;			OUT_795 <= inform_L [794][0] ;			OUT_796 <= inform_L [795][0] ;			OUT_797 <= inform_L [796][0] ;			OUT_798 <= inform_L [797][0] ;			OUT_799 <= inform_L [798][0] ;			OUT_800 <= inform_L [799][0] ;			OUT_801 <= inform_L [800][0] ;			OUT_802 <= inform_L [801][0] ;			OUT_803 <= inform_L [802][0] ;			OUT_804 <= inform_L [803][0] ;			OUT_805 <= inform_L [804][0] ;			OUT_806 <= inform_L [805][0] ;			OUT_807 <= inform_L [806][0] ;			OUT_808 <= inform_L [807][0] ;			OUT_809 <= inform_L [808][0] ;			OUT_810 <= inform_L [809][0] ;			OUT_811 <= inform_L [810][0] ;			OUT_812 <= inform_L [811][0] ;			OUT_813 <= inform_L [812][0] ;			OUT_814 <= inform_L [813][0] ;			OUT_815 <= inform_L [814][0] ;			OUT_816 <= inform_L [815][0] ;			OUT_817 <= inform_L [816][0] ;			OUT_818 <= inform_L [817][0] ;			OUT_819 <= inform_L [818][0] ;			OUT_820 <= inform_L [819][0] ;			OUT_821 <= inform_L [820][0] ;			OUT_822 <= inform_L [821][0] ;			OUT_823 <= inform_L [822][0] ;			OUT_824 <= inform_L [823][0] ;			OUT_825 <= inform_L [824][0] ;			OUT_826 <= inform_L [825][0] ;			OUT_827 <= inform_L [826][0] ;			OUT_828 <= inform_L [827][0] ;			OUT_829 <= inform_L [828][0] ;			OUT_830 <= inform_L [829][0] ;			OUT_831 <= inform_L [830][0] ;			OUT_832 <= inform_L [831][0] ;			OUT_833 <= inform_L [832][0] ;			OUT_834 <= inform_L [833][0] ;			OUT_835 <= inform_L [834][0] ;			OUT_836 <= inform_L [835][0] ;			OUT_837 <= inform_L [836][0] ;			OUT_838 <= inform_L [837][0] ;			OUT_839 <= inform_L [838][0] ;			OUT_840 <= inform_L [839][0] ;			OUT_841 <= inform_L [840][0] ;			OUT_842 <= inform_L [841][0] ;			OUT_843 <= inform_L [842][0] ;			OUT_844 <= inform_L [843][0] ;			OUT_845 <= inform_L [844][0] ;			OUT_846 <= inform_L [845][0] ;			OUT_847 <= inform_L [846][0] ;			OUT_848 <= inform_L [847][0] ;			OUT_849 <= inform_L [848][0] ;			OUT_850 <= inform_L [849][0] ;			OUT_851 <= inform_L [850][0] ;			OUT_852 <= inform_L [851][0] ;			OUT_853 <= inform_L [852][0] ;			OUT_854 <= inform_L [853][0] ;			OUT_855 <= inform_L [854][0] ;			OUT_856 <= inform_L [855][0] ;			OUT_857 <= inform_L [856][0] ;			OUT_858 <= inform_L [857][0] ;			OUT_859 <= inform_L [858][0] ;			OUT_860 <= inform_L [859][0] ;			OUT_861 <= inform_L [860][0] ;			OUT_862 <= inform_L [861][0] ;			OUT_863 <= inform_L [862][0] ;			OUT_864 <= inform_L [863][0] ;			OUT_865 <= inform_L [864][0] ;			OUT_866 <= inform_L [865][0] ;			OUT_867 <= inform_L [866][0] ;			OUT_868 <= inform_L [867][0] ;			OUT_869 <= inform_L [868][0] ;			OUT_870 <= inform_L [869][0] ;			OUT_871 <= inform_L [870][0] ;			OUT_872 <= inform_L [871][0] ;			OUT_873 <= inform_L [872][0] ;			OUT_874 <= inform_L [873][0] ;			OUT_875 <= inform_L [874][0] ;			OUT_876 <= inform_L [875][0] ;			OUT_877 <= inform_L [876][0] ;			OUT_878 <= inform_L [877][0] ;			OUT_879 <= inform_L [878][0] ;			OUT_880 <= inform_L [879][0] ;			OUT_881 <= inform_L [880][0] ;			OUT_882 <= inform_L [881][0] ;			OUT_883 <= inform_L [882][0] ;			OUT_884 <= inform_L [883][0] ;			OUT_885 <= inform_L [884][0] ;			OUT_886 <= inform_L [885][0] ;			OUT_887 <= inform_L [886][0] ;			OUT_888 <= inform_L [887][0] ;			OUT_889 <= inform_L [888][0] ;			OUT_890 <= inform_L [889][0] ;			OUT_891 <= inform_L [890][0] ;			OUT_892 <= inform_L [891][0] ;			OUT_893 <= inform_L [892][0] ;			OUT_894 <= inform_L [893][0] ;			OUT_895 <= inform_L [894][0] ;			OUT_896 <= inform_L [895][0] ;			OUT_897 <= inform_L [896][0] ;			OUT_898 <= inform_L [897][0] ;			OUT_899 <= inform_L [898][0] ;			OUT_900 <= inform_L [899][0] ;			OUT_901 <= inform_L [900][0] ;			OUT_902 <= inform_L [901][0] ;			OUT_903 <= inform_L [902][0] ;			OUT_904 <= inform_L [903][0] ;			OUT_905 <= inform_L [904][0] ;			OUT_906 <= inform_L [905][0] ;			OUT_907 <= inform_L [906][0] ;			OUT_908 <= inform_L [907][0] ;			OUT_909 <= inform_L [908][0] ;			OUT_910 <= inform_L [909][0] ;			OUT_911 <= inform_L [910][0] ;			OUT_912 <= inform_L [911][0] ;			OUT_913 <= inform_L [912][0] ;			OUT_914 <= inform_L [913][0] ;			OUT_915 <= inform_L [914][0] ;			OUT_916 <= inform_L [915][0] ;			OUT_917 <= inform_L [916][0] ;			OUT_918 <= inform_L [917][0] ;			OUT_919 <= inform_L [918][0] ;			OUT_920 <= inform_L [919][0] ;			OUT_921 <= inform_L [920][0] ;			OUT_922 <= inform_L [921][0] ;			OUT_923 <= inform_L [922][0] ;			OUT_924 <= inform_L [923][0] ;			OUT_925 <= inform_L [924][0] ;			OUT_926 <= inform_L [925][0] ;			OUT_927 <= inform_L [926][0] ;			OUT_928 <= inform_L [927][0] ;			OUT_929 <= inform_L [928][0] ;			OUT_930 <= inform_L [929][0] ;			OUT_931 <= inform_L [930][0] ;			OUT_932 <= inform_L [931][0] ;			OUT_933 <= inform_L [932][0] ;			OUT_934 <= inform_L [933][0] ;			OUT_935 <= inform_L [934][0] ;			OUT_936 <= inform_L [935][0] ;			OUT_937 <= inform_L [936][0] ;			OUT_938 <= inform_L [937][0] ;			OUT_939 <= inform_L [938][0] ;			OUT_940 <= inform_L [939][0] ;			OUT_941 <= inform_L [940][0] ;			OUT_942 <= inform_L [941][0] ;			OUT_943 <= inform_L [942][0] ;			OUT_944 <= inform_L [943][0] ;			OUT_945 <= inform_L [944][0] ;			OUT_946 <= inform_L [945][0] ;			OUT_947 <= inform_L [946][0] ;			OUT_948 <= inform_L [947][0] ;			OUT_949 <= inform_L [948][0] ;			OUT_950 <= inform_L [949][0] ;			OUT_951 <= inform_L [950][0] ;			OUT_952 <= inform_L [951][0] ;			OUT_953 <= inform_L [952][0] ;			OUT_954 <= inform_L [953][0] ;			OUT_955 <= inform_L [954][0] ;			OUT_956 <= inform_L [955][0] ;			OUT_957 <= inform_L [956][0] ;			OUT_958 <= inform_L [957][0] ;			OUT_959 <= inform_L [958][0] ;			OUT_960 <= inform_L [959][0] ;			OUT_961 <= inform_L [960][0] ;			OUT_962 <= inform_L [961][0] ;			OUT_963 <= inform_L [962][0] ;			OUT_964 <= inform_L [963][0] ;			OUT_965 <= inform_L [964][0] ;			OUT_966 <= inform_L [965][0] ;			OUT_967 <= inform_L [966][0] ;			OUT_968 <= inform_L [967][0] ;			OUT_969 <= inform_L [968][0] ;			OUT_970 <= inform_L [969][0] ;			OUT_971 <= inform_L [970][0] ;			OUT_972 <= inform_L [971][0] ;			OUT_973 <= inform_L [972][0] ;			OUT_974 <= inform_L [973][0] ;			OUT_975 <= inform_L [974][0] ;			OUT_976 <= inform_L [975][0] ;			OUT_977 <= inform_L [976][0] ;			OUT_978 <= inform_L [977][0] ;			OUT_979 <= inform_L [978][0] ;			OUT_980 <= inform_L [979][0] ;			OUT_981 <= inform_L [980][0] ;			OUT_982 <= inform_L [981][0] ;			OUT_983 <= inform_L [982][0] ;			OUT_984 <= inform_L [983][0] ;			OUT_985 <= inform_L [984][0] ;			OUT_986 <= inform_L [985][0] ;			OUT_987 <= inform_L [986][0] ;			OUT_988 <= inform_L [987][0] ;			OUT_989 <= inform_L [988][0] ;			OUT_990 <= inform_L [989][0] ;			OUT_991 <= inform_L [990][0] ;			OUT_992 <= inform_L [991][0] ;			OUT_993 <= inform_L [992][0] ;			OUT_994 <= inform_L [993][0] ;			OUT_995 <= inform_L [994][0] ;			OUT_996 <= inform_L [995][0] ;			OUT_997 <= inform_L [996][0] ;			OUT_998 <= inform_L [997][0] ;			OUT_999 <= inform_L [998][0] ;			OUT_1000 <= inform_L [999][0] ;			OUT_1001 <= inform_L [1000][0] ;			OUT_1002 <= inform_L [1001][0] ;			OUT_1003 <= inform_L [1002][0] ;			OUT_1004 <= inform_L [1003][0] ;			OUT_1005 <= inform_L [1004][0] ;			OUT_1006 <= inform_L [1005][0] ;			OUT_1007 <= inform_L [1006][0] ;			OUT_1008 <= inform_L [1007][0] ;			OUT_1009 <= inform_L [1008][0] ;			OUT_1010 <= inform_L [1009][0] ;			OUT_1011 <= inform_L [1010][0] ;			OUT_1012 <= inform_L [1011][0] ;			OUT_1013 <= inform_L [1012][0] ;			OUT_1014 <= inform_L [1013][0] ;			OUT_1015 <= inform_L [1014][0] ;			OUT_1016 <= inform_L [1015][0] ;			OUT_1017 <= inform_L [1016][0] ;			OUT_1018 <= inform_L [1017][0] ;			OUT_1019 <= inform_L [1018][0] ;			OUT_1020 <= inform_L [1019][0] ;			OUT_1021 <= inform_L [1020][0] ;			OUT_1022 <= inform_L [1021][0] ;			OUT_1023 <= inform_L [1022][0] ;			OUT_1024 <= inform_L [1023][0] ;		end	end
endmodule