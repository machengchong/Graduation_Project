`define iteration_times 40 module bp_128_64 #(	parameter integer BIT = 8)(	input clk,	input rst_n,	input start,	output reg en_busy,	input [BIT - 1:0] LLR_1,	input [BIT - 1:0] LLR_2,	input [BIT - 1:0] LLR_3,	input [BIT - 1:0] LLR_4,	input [BIT - 1:0] LLR_5,	input [BIT - 1:0] LLR_6,	input [BIT - 1:0] LLR_7,	input [BIT - 1:0] LLR_8,	input [BIT - 1:0] LLR_9,	input [BIT - 1:0] LLR_10,	input [BIT - 1:0] LLR_11,	input [BIT - 1:0] LLR_12,	input [BIT - 1:0] LLR_13,	input [BIT - 1:0] LLR_14,	input [BIT - 1:0] LLR_15,	input [BIT - 1:0] LLR_16,	input [BIT - 1:0] LLR_17,	input [BIT - 1:0] LLR_18,	input [BIT - 1:0] LLR_19,	input [BIT - 1:0] LLR_20,	input [BIT - 1:0] LLR_21,	input [BIT - 1:0] LLR_22,	input [BIT - 1:0] LLR_23,	input [BIT - 1:0] LLR_24,	input [BIT - 1:0] LLR_25,	input [BIT - 1:0] LLR_26,	input [BIT - 1:0] LLR_27,	input [BIT - 1:0] LLR_28,	input [BIT - 1:0] LLR_29,	input [BIT - 1:0] LLR_30,	input [BIT - 1:0] LLR_31,	input [BIT - 1:0] LLR_32,	input [BIT - 1:0] LLR_33,	input [BIT - 1:0] LLR_34,	input [BIT - 1:0] LLR_35,	input [BIT - 1:0] LLR_36,	input [BIT - 1:0] LLR_37,	input [BIT - 1:0] LLR_38,	input [BIT - 1:0] LLR_39,	input [BIT - 1:0] LLR_40,	input [BIT - 1:0] LLR_41,	input [BIT - 1:0] LLR_42,	input [BIT - 1:0] LLR_43,	input [BIT - 1:0] LLR_44,	input [BIT - 1:0] LLR_45,	input [BIT - 1:0] LLR_46,	input [BIT - 1:0] LLR_47,	input [BIT - 1:0] LLR_48,	input [BIT - 1:0] LLR_49,	input [BIT - 1:0] LLR_50,	input [BIT - 1:0] LLR_51,	input [BIT - 1:0] LLR_52,	input [BIT - 1:0] LLR_53,	input [BIT - 1:0] LLR_54,	input [BIT - 1:0] LLR_55,	input [BIT - 1:0] LLR_56,	input [BIT - 1:0] LLR_57,	input [BIT - 1:0] LLR_58,	input [BIT - 1:0] LLR_59,	input [BIT - 1:0] LLR_60,	input [BIT - 1:0] LLR_61,	input [BIT - 1:0] LLR_62,	input [BIT - 1:0] LLR_63,	input [BIT - 1:0] LLR_64,	input [BIT - 1:0] LLR_65,	input [BIT - 1:0] LLR_66,	input [BIT - 1:0] LLR_67,	input [BIT - 1:0] LLR_68,	input [BIT - 1:0] LLR_69,	input [BIT - 1:0] LLR_70,	input [BIT - 1:0] LLR_71,	input [BIT - 1:0] LLR_72,	input [BIT - 1:0] LLR_73,	input [BIT - 1:0] LLR_74,	input [BIT - 1:0] LLR_75,	input [BIT - 1:0] LLR_76,	input [BIT - 1:0] LLR_77,	input [BIT - 1:0] LLR_78,	input [BIT - 1:0] LLR_79,	input [BIT - 1:0] LLR_80,	input [BIT - 1:0] LLR_81,	input [BIT - 1:0] LLR_82,	input [BIT - 1:0] LLR_83,	input [BIT - 1:0] LLR_84,	input [BIT - 1:0] LLR_85,	input [BIT - 1:0] LLR_86,	input [BIT - 1:0] LLR_87,	input [BIT - 1:0] LLR_88,	input [BIT - 1:0] LLR_89,	input [BIT - 1:0] LLR_90,	input [BIT - 1:0] LLR_91,	input [BIT - 1:0] LLR_92,	input [BIT - 1:0] LLR_93,	input [BIT - 1:0] LLR_94,	input [BIT - 1:0] LLR_95,	input [BIT - 1:0] LLR_96,	input [BIT - 1:0] LLR_97,	input [BIT - 1:0] LLR_98,	input [BIT - 1:0] LLR_99,	input [BIT - 1:0] LLR_100,	input [BIT - 1:0] LLR_101,	input [BIT - 1:0] LLR_102,	input [BIT - 1:0] LLR_103,	input [BIT - 1:0] LLR_104,	input [BIT - 1:0] LLR_105,	input [BIT - 1:0] LLR_106,	input [BIT - 1:0] LLR_107,	input [BIT - 1:0] LLR_108,	input [BIT - 1:0] LLR_109,	input [BIT - 1:0] LLR_110,	input [BIT - 1:0] LLR_111,	input [BIT - 1:0] LLR_112,	input [BIT - 1:0] LLR_113,	input [BIT - 1:0] LLR_114,	input [BIT - 1:0] LLR_115,	input [BIT - 1:0] LLR_116,	input [BIT - 1:0] LLR_117,	input [BIT - 1:0] LLR_118,	input [BIT - 1:0] LLR_119,	input [BIT - 1:0] LLR_120,	input [BIT - 1:0] LLR_121,	input [BIT - 1:0] LLR_122,	input [BIT - 1:0] LLR_123,	input [BIT - 1:0] LLR_124,	input [BIT - 1:0] LLR_125,	input [BIT - 1:0] LLR_126,	input [BIT - 1:0] LLR_127,	input [BIT - 1:0] LLR_128,	output reg [BIT - 1:0] OUT_1,	output reg [BIT - 1:0] OUT_2,	output reg [BIT - 1:0] OUT_3,	output reg [BIT - 1:0] OUT_4,	output reg [BIT - 1:0] OUT_5,	output reg [BIT - 1:0] OUT_6,	output reg [BIT - 1:0] OUT_7,	output reg [BIT - 1:0] OUT_8,	output reg [BIT - 1:0] OUT_9,	output reg [BIT - 1:0] OUT_10,	output reg [BIT - 1:0] OUT_11,	output reg [BIT - 1:0] OUT_12,	output reg [BIT - 1:0] OUT_13,	output reg [BIT - 1:0] OUT_14,	output reg [BIT - 1:0] OUT_15,	output reg [BIT - 1:0] OUT_16,	output reg [BIT - 1:0] OUT_17,	output reg [BIT - 1:0] OUT_18,	output reg [BIT - 1:0] OUT_19,	output reg [BIT - 1:0] OUT_20,	output reg [BIT - 1:0] OUT_21,	output reg [BIT - 1:0] OUT_22,	output reg [BIT - 1:0] OUT_23,	output reg [BIT - 1:0] OUT_24,	output reg [BIT - 1:0] OUT_25,	output reg [BIT - 1:0] OUT_26,	output reg [BIT - 1:0] OUT_27,	output reg [BIT - 1:0] OUT_28,	output reg [BIT - 1:0] OUT_29,	output reg [BIT - 1:0] OUT_30,	output reg [BIT - 1:0] OUT_31,	output reg [BIT - 1:0] OUT_32,	output reg [BIT - 1:0] OUT_33,	output reg [BIT - 1:0] OUT_34,	output reg [BIT - 1:0] OUT_35,	output reg [BIT - 1:0] OUT_36,	output reg [BIT - 1:0] OUT_37,	output reg [BIT - 1:0] OUT_38,	output reg [BIT - 1:0] OUT_39,	output reg [BIT - 1:0] OUT_40,	output reg [BIT - 1:0] OUT_41,	output reg [BIT - 1:0] OUT_42,	output reg [BIT - 1:0] OUT_43,	output reg [BIT - 1:0] OUT_44,	output reg [BIT - 1:0] OUT_45,	output reg [BIT - 1:0] OUT_46,	output reg [BIT - 1:0] OUT_47,	output reg [BIT - 1:0] OUT_48,	output reg [BIT - 1:0] OUT_49,	output reg [BIT - 1:0] OUT_50,	output reg [BIT - 1:0] OUT_51,	output reg [BIT - 1:0] OUT_52,	output reg [BIT - 1:0] OUT_53,	output reg [BIT - 1:0] OUT_54,	output reg [BIT - 1:0] OUT_55,	output reg [BIT - 1:0] OUT_56,	output reg [BIT - 1:0] OUT_57,	output reg [BIT - 1:0] OUT_58,	output reg [BIT - 1:0] OUT_59,	output reg [BIT - 1:0] OUT_60,	output reg [BIT - 1:0] OUT_61,	output reg [BIT - 1:0] OUT_62,	output reg [BIT - 1:0] OUT_63,	output reg [BIT - 1:0] OUT_64,	output reg [BIT - 1:0] OUT_65,	output reg [BIT - 1:0] OUT_66,	output reg [BIT - 1:0] OUT_67,	output reg [BIT - 1:0] OUT_68,	output reg [BIT - 1:0] OUT_69,	output reg [BIT - 1:0] OUT_70,	output reg [BIT - 1:0] OUT_71,	output reg [BIT - 1:0] OUT_72,	output reg [BIT - 1:0] OUT_73,	output reg [BIT - 1:0] OUT_74,	output reg [BIT - 1:0] OUT_75,	output reg [BIT - 1:0] OUT_76,	output reg [BIT - 1:0] OUT_77,	output reg [BIT - 1:0] OUT_78,	output reg [BIT - 1:0] OUT_79,	output reg [BIT - 1:0] OUT_80,	output reg [BIT - 1:0] OUT_81,	output reg [BIT - 1:0] OUT_82,	output reg [BIT - 1:0] OUT_83,	output reg [BIT - 1:0] OUT_84,	output reg [BIT - 1:0] OUT_85,	output reg [BIT - 1:0] OUT_86,	output reg [BIT - 1:0] OUT_87,	output reg [BIT - 1:0] OUT_88,	output reg [BIT - 1:0] OUT_89,	output reg [BIT - 1:0] OUT_90,	output reg [BIT - 1:0] OUT_91,	output reg [BIT - 1:0] OUT_92,	output reg [BIT - 1:0] OUT_93,	output reg [BIT - 1:0] OUT_94,	output reg [BIT - 1:0] OUT_95,	output reg [BIT - 1:0] OUT_96,	output reg [BIT - 1:0] OUT_97,	output reg [BIT - 1:0] OUT_98,	output reg [BIT - 1:0] OUT_99,	output reg [BIT - 1:0] OUT_100,	output reg [BIT - 1:0] OUT_101,	output reg [BIT - 1:0] OUT_102,	output reg [BIT - 1:0] OUT_103,	output reg [BIT - 1:0] OUT_104,	output reg [BIT - 1:0] OUT_105,	output reg [BIT - 1:0] OUT_106,	output reg [BIT - 1:0] OUT_107,	output reg [BIT - 1:0] OUT_108,	output reg [BIT - 1:0] OUT_109,	output reg [BIT - 1:0] OUT_110,	output reg [BIT - 1:0] OUT_111,	output reg [BIT - 1:0] OUT_112,	output reg [BIT - 1:0] OUT_113,	output reg [BIT - 1:0] OUT_114,	output reg [BIT - 1:0] OUT_115,	output reg [BIT - 1:0] OUT_116,	output reg [BIT - 1:0] OUT_117,	output reg [BIT - 1:0] OUT_118,	output reg [BIT - 1:0] OUT_119,	output reg [BIT - 1:0] OUT_120,	output reg [BIT - 1:0] OUT_121,	output reg [BIT - 1:0] OUT_122,	output reg [BIT - 1:0] OUT_123,	output reg [BIT - 1:0] OUT_124,	output reg [BIT - 1:0] OUT_125,	output reg [BIT - 1:0] OUT_126,	output reg [BIT - 1:0] OUT_127,	output reg [BIT - 1:0] OUT_128);	integer x, y;
	reg [BIT - 1:0] inform_R [128-1:0][8-1:0];	reg [BIT - 1:0] inform_L [128-1:0][8-1:0];	localparam IDLE = 2'b00;	localparam BUSY_LEFT = 2'b01;	localparam BUSY_RIGHT = 2'b10;	reg [1:0] bp_state,bp_next_state;	reg [7-1:0] cell_enable,w2r;	reg left_over_flag,right_over_flag,init_over_flag;	wire bp_over_flag;	reg [6:0]itera_time;
	always @(posedge clk or negedge rst_n) begin		if (!rst_n) begin			bp_state <= IDLE;		end		else begin			bp_state <= bp_next_state;		end	end
	always @(*) begin		case (bp_state)			IDLE:			if (init_over_flag) begin				bp_next_state <= BUSY_LEFT;			end			else begin				bp_next_state <= IDLE;			end
			BUSY_LEFT:			if (left_over_flag) begin				bp_next_state <= BUSY_RIGHT;			end			else begin				 bp_next_state <= BUSY_LEFT;			end
			BUSY_RIGHT:			if (bp_over_flag) begin				bp_next_state <= IDLE;			end			else if (right_over_flag) begin				bp_next_state <= BUSY_LEFT;			end			else begin				 bp_next_state <= BUSY_RIGHT;			end
			default: bp_next_state <= IDLE;		endcase	end
	reg [1:0] clk_counter;
	always @(posedge clk) begin		case (bp_next_state)			IDLE:			begin				left_over_flag <= 0;				right_over_flag <= 0;				itera_time <= 7'b0;				clk_counter <= 2'b0;				if (start) begin					cell_enable <=7'b1;					w2r <= 7;					init_over_flag <= 1;					en_busy <= 1;				end				else begin					cell_enable <=7'b0;					w2r <= 0;					init_over_flag <= 0;					en_busy <= 0;				end			end
			BUSY_LEFT:			begin				init_over_flag <= 0;				en_busy <= 1;				right_over_flag <= 0;				if (clk_counter == 2'b11) begin					clk_counter <= 2'b00;					if (cell_enable == 64) begin						left_over_flag <= 1;						cell_enable <= cell_enable >> 1;						w2r <= w2r + 1;					end					else begin						left_over_flag <= 0;						cell_enable <= cell_enable << 1;						w2r <= w2r - 1;					end				end				else begin					clk_counter <= clk_counter + 1;				end			end
			BUSY_RIGHT:			begin				en_busy <= 1;				left_over_flag <= 0;				if (clk_counter == 2'b11) begin					clk_counter <= 2'b00;					if (cell_enable == 1) begin						right_over_flag <= 1;						itera_time <= itera_time + 1;						cell_enable <= cell_enable << 1;						w2r <= w2r - 1;					end					else begin						right_over_flag <= 0;						cell_enable <= cell_enable >> 1;						w2r <= w2r + 1;					end				end				else begin					clk_counter <= clk_counter + 1;				end			end
			default:			begin				left_over_flag <= 0;				right_over_flag <= 0;				itera_time <= 7'b0;				clk_counter <= 2'b0;				if (start) begin					cell_enable <=7'b1;					w2r <= 7;					init_over_flag <= 1;					en_busy <= 1;				end				else begin					cell_enable <=7'b0;					w2r <= 0;					init_over_flag <= 0;					en_busy <= 0;				end			end
		endcase	end
	reg[BIT - 1:0] r_cell_reg[128-1:0];	reg[BIT - 1:0] l_cell_reg[128-1:0];	wire[BIT - 1:0] r_cell_wire[128-1:0];	wire[BIT - 1:0] l_cell_wire[128-1:0];
	always @(posedge clk) begin		case (bp_next_state)			IDLE:			begin				if (start) begin					inform_R [0][0] <= 8'b0111_1111;					inform_R [1][0] <= 8'b0111_1111;					inform_R [2][0] <= 8'b0111_1111;					inform_R [3][0] <= 8'b0111_1111;					inform_R [4][0] <= 8'b0111_1111;					inform_R [5][0] <= 8'b0111_1111;					inform_R [6][0] <= 8'b0111_1111;					inform_R [7][0] <= 8'b0111_1111;					inform_R [8][0] <= 8'b0111_1111;					inform_R [9][0] <= 8'b0111_1111;					inform_R [10][0] <= 8'b0111_1111;					inform_R [11][0] <= 8'b0111_1111;					inform_R [12][0] <= 8'b0111_1111;					inform_R [13][0] <= 8'b0111_1111;					inform_R [14][0] <= 8'b0111_1111;					inform_R [15][0] <= 8'b0111_1111;					inform_R [16][0] <= 8'b0111_1111;					inform_R [17][0] <= 8'b0111_1111;					inform_R [18][0] <= 8'b0111_1111;					inform_R [19][0] <= 8'b0111_1111;					inform_R [20][0] <= 8'b0111_1111;					inform_R [21][0] <= 8'b0111_1111;					inform_R [22][0] <= 8'b0111_1111;					inform_R [23][0] <= 8'b0111_1111;					inform_R [24][0] <= 8'b0111_1111;					inform_R [25][0] <= 8'b0111_1111;					inform_R [26][0] <= 8'b0111_1111;					inform_R [27][0] <= 8'b0111_1111;					inform_R [28][0] <= 8'b0111_1111;					inform_R [29][0] <= 8'b0111_1111;					inform_R [30][0] <= 8'b0111_1111;					inform_R [31][0] <= 8'b0000_0000;					inform_R [32][0] <= 8'b0111_1111;					inform_R [33][0] <= 8'b0111_1111;					inform_R [34][0] <= 8'b0111_1111;					inform_R [35][0] <= 8'b0111_1111;					inform_R [36][0] <= 8'b0111_1111;					inform_R [37][0] <= 8'b0111_1111;					inform_R [38][0] <= 8'b0111_1111;					inform_R [39][0] <= 8'b0111_1111;					inform_R [40][0] <= 8'b0111_1111;					inform_R [41][0] <= 8'b0111_1111;					inform_R [42][0] <= 8'b0111_1111;					inform_R [43][0] <= 8'b0111_1111;					inform_R [44][0] <= 8'b0111_1111;					inform_R [45][0] <= 8'b0000_0000;					inform_R [46][0] <= 8'b0000_0000;					inform_R [47][0] <= 8'b0000_0000;					inform_R [48][0] <= 8'b0111_1111;					inform_R [49][0] <= 8'b0111_1111;					inform_R [50][0] <= 8'b0111_1111;					inform_R [51][0] <= 8'b0000_0000;					inform_R [52][0] <= 8'b0111_1111;					inform_R [53][0] <= 8'b0000_0000;					inform_R [54][0] <= 8'b0000_0000;					inform_R [55][0] <= 8'b0000_0000;					inform_R [56][0] <= 8'b0111_1111;					inform_R [57][0] <= 8'b0000_0000;					inform_R [58][0] <= 8'b0000_0000;					inform_R [59][0] <= 8'b0000_0000;					inform_R [60][0] <= 8'b0000_0000;					inform_R [61][0] <= 8'b0000_0000;					inform_R [62][0] <= 8'b0000_0000;					inform_R [63][0] <= 8'b0000_0000;					inform_R [64][0] <= 8'b0111_1111;					inform_R [65][0] <= 8'b0111_1111;					inform_R [66][0] <= 8'b0111_1111;					inform_R [67][0] <= 8'b0111_1111;					inform_R [68][0] <= 8'b0111_1111;					inform_R [69][0] <= 8'b0111_1111;					inform_R [70][0] <= 8'b0111_1111;					inform_R [71][0] <= 8'b0000_0000;					inform_R [72][0] <= 8'b0111_1111;					inform_R [73][0] <= 8'b0111_1111;					inform_R [74][0] <= 8'b0111_1111;					inform_R [75][0] <= 8'b0000_0000;					inform_R [76][0] <= 8'b0111_1111;					inform_R [77][0] <= 8'b0000_0000;					inform_R [78][0] <= 8'b0000_0000;					inform_R [79][0] <= 8'b0000_0000;					inform_R [80][0] <= 8'b0111_1111;					inform_R [81][0] <= 8'b0111_1111;					inform_R [82][0] <= 8'b0111_1111;					inform_R [83][0] <= 8'b0000_0000;					inform_R [84][0] <= 8'b0000_0000;					inform_R [85][0] <= 8'b0000_0000;					inform_R [86][0] <= 8'b0000_0000;					inform_R [87][0] <= 8'b0000_0000;					inform_R [88][0] <= 8'b0000_0000;					inform_R [89][0] <= 8'b0000_0000;					inform_R [90][0] <= 8'b0000_0000;					inform_R [91][0] <= 8'b0000_0000;					inform_R [92][0] <= 8'b0000_0000;					inform_R [93][0] <= 8'b0000_0000;					inform_R [94][0] <= 8'b0000_0000;					inform_R [95][0] <= 8'b0000_0000;					inform_R [96][0] <= 8'b0111_1111;					inform_R [97][0] <= 8'b0000_0000;					inform_R [98][0] <= 8'b0000_0000;					inform_R [99][0] <= 8'b0000_0000;					inform_R [100][0] <= 8'b0000_0000;					inform_R [101][0] <= 8'b0000_0000;					inform_R [102][0] <= 8'b0000_0000;					inform_R [103][0] <= 8'b0000_0000;					inform_R [104][0] <= 8'b0000_0000;					inform_R [105][0] <= 8'b0000_0000;					inform_R [106][0] <= 8'b0000_0000;					inform_R [107][0] <= 8'b0000_0000;					inform_R [108][0] <= 8'b0000_0000;					inform_R [109][0] <= 8'b0000_0000;					inform_R [110][0] <= 8'b0000_0000;					inform_R [111][0] <= 8'b0000_0000;					inform_R [112][0] <= 8'b0000_0000;					inform_R [113][0] <= 8'b0000_0000;					inform_R [114][0] <= 8'b0000_0000;					inform_R [115][0] <= 8'b0000_0000;					inform_R [116][0] <= 8'b0000_0000;					inform_R [117][0] <= 8'b0000_0000;					inform_R [118][0] <= 8'b0000_0000;					inform_R [119][0] <= 8'b0000_0000;					inform_R [120][0] <= 8'b0000_0000;					inform_R [121][0] <= 8'b0000_0000;					inform_R [122][0] <= 8'b0000_0000;					inform_R [123][0] <= 8'b0000_0000;					inform_R [124][0] <= 8'b0000_0000;					inform_R [125][0] <= 8'b0000_0000;					inform_R [126][0] <= 8'b0000_0000;					inform_R [127][0] <= 8'b0000_0000;					inform_L [0][7] <= LLR_1;					inform_L [1][7] <= LLR_2;					inform_L [2][7] <= LLR_3;					inform_L [3][7] <= LLR_4;					inform_L [4][7] <= LLR_5;					inform_L [5][7] <= LLR_6;					inform_L [6][7] <= LLR_7;					inform_L [7][7] <= LLR_8;					inform_L [8][7] <= LLR_9;					inform_L [9][7] <= LLR_10;					inform_L [10][7] <= LLR_11;					inform_L [11][7] <= LLR_12;					inform_L [12][7] <= LLR_13;					inform_L [13][7] <= LLR_14;					inform_L [14][7] <= LLR_15;					inform_L [15][7] <= LLR_16;					inform_L [16][7] <= LLR_17;					inform_L [17][7] <= LLR_18;					inform_L [18][7] <= LLR_19;					inform_L [19][7] <= LLR_20;					inform_L [20][7] <= LLR_21;					inform_L [21][7] <= LLR_22;					inform_L [22][7] <= LLR_23;					inform_L [23][7] <= LLR_24;					inform_L [24][7] <= LLR_25;					inform_L [25][7] <= LLR_26;					inform_L [26][7] <= LLR_27;					inform_L [27][7] <= LLR_28;					inform_L [28][7] <= LLR_29;					inform_L [29][7] <= LLR_30;					inform_L [30][7] <= LLR_31;					inform_L [31][7] <= LLR_32;					inform_L [32][7] <= LLR_33;					inform_L [33][7] <= LLR_34;					inform_L [34][7] <= LLR_35;					inform_L [35][7] <= LLR_36;					inform_L [36][7] <= LLR_37;					inform_L [37][7] <= LLR_38;					inform_L [38][7] <= LLR_39;					inform_L [39][7] <= LLR_40;					inform_L [40][7] <= LLR_41;					inform_L [41][7] <= LLR_42;					inform_L [42][7] <= LLR_43;					inform_L [43][7] <= LLR_44;					inform_L [44][7] <= LLR_45;					inform_L [45][7] <= LLR_46;					inform_L [46][7] <= LLR_47;					inform_L [47][7] <= LLR_48;					inform_L [48][7] <= LLR_49;					inform_L [49][7] <= LLR_50;					inform_L [50][7] <= LLR_51;					inform_L [51][7] <= LLR_52;					inform_L [52][7] <= LLR_53;					inform_L [53][7] <= LLR_54;					inform_L [54][7] <= LLR_55;					inform_L [55][7] <= LLR_56;					inform_L [56][7] <= LLR_57;					inform_L [57][7] <= LLR_58;					inform_L [58][7] <= LLR_59;					inform_L [59][7] <= LLR_60;					inform_L [60][7] <= LLR_61;					inform_L [61][7] <= LLR_62;					inform_L [62][7] <= LLR_63;					inform_L [63][7] <= LLR_64;					inform_L [64][7] <= LLR_65;					inform_L [65][7] <= LLR_66;					inform_L [66][7] <= LLR_67;					inform_L [67][7] <= LLR_68;					inform_L [68][7] <= LLR_69;					inform_L [69][7] <= LLR_70;					inform_L [70][7] <= LLR_71;					inform_L [71][7] <= LLR_72;					inform_L [72][7] <= LLR_73;					inform_L [73][7] <= LLR_74;					inform_L [74][7] <= LLR_75;					inform_L [75][7] <= LLR_76;					inform_L [76][7] <= LLR_77;					inform_L [77][7] <= LLR_78;					inform_L [78][7] <= LLR_79;					inform_L [79][7] <= LLR_80;					inform_L [80][7] <= LLR_81;					inform_L [81][7] <= LLR_82;					inform_L [82][7] <= LLR_83;					inform_L [83][7] <= LLR_84;					inform_L [84][7] <= LLR_85;					inform_L [85][7] <= LLR_86;					inform_L [86][7] <= LLR_87;					inform_L [87][7] <= LLR_88;					inform_L [88][7] <= LLR_89;					inform_L [89][7] <= LLR_90;					inform_L [90][7] <= LLR_91;					inform_L [91][7] <= LLR_92;					inform_L [92][7] <= LLR_93;					inform_L [93][7] <= LLR_94;					inform_L [94][7] <= LLR_95;					inform_L [95][7] <= LLR_96;					inform_L [96][7] <= LLR_97;					inform_L [97][7] <= LLR_98;					inform_L [98][7] <= LLR_99;					inform_L [99][7] <= LLR_100;					inform_L [100][7] <= LLR_101;					inform_L [101][7] <= LLR_102;					inform_L [102][7] <= LLR_103;					inform_L [103][7] <= LLR_104;					inform_L [104][7] <= LLR_105;					inform_L [105][7] <= LLR_106;					inform_L [106][7] <= LLR_107;					inform_L [107][7] <= LLR_108;					inform_L [108][7] <= LLR_109;					inform_L [109][7] <= LLR_110;					inform_L [110][7] <= LLR_111;					inform_L [111][7] <= LLR_112;					inform_L [112][7] <= LLR_113;					inform_L [113][7] <= LLR_114;					inform_L [114][7] <= LLR_115;					inform_L [115][7] <= LLR_116;					inform_L [116][7] <= LLR_117;					inform_L [117][7] <= LLR_118;					inform_L [118][7] <= LLR_119;					inform_L [119][7] <= LLR_120;					inform_L [120][7] <= LLR_121;					inform_L [121][7] <= LLR_122;					inform_L [122][7] <= LLR_123;					inform_L [123][7] <= LLR_124;					inform_L [124][7] <= LLR_125;					inform_L [125][7] <= LLR_126;					inform_L [126][7] <= LLR_127;					inform_L [127][7] <= LLR_128;				end				for (x = 0; x < 128; x = x + 1)					for (y = 0; y < 7; y = y + 1)					begin						inform_R[x][y+1] <= 8'd0;						inform_L[x][y] <= 8'd0;					end			end
			BUSY_LEFT:			begin				if(clk_counter == 2'b11)begin					case (w2r)						1:						begin							inform_R[0][1] = r_cell_wire[0];							inform_R[1][1] = r_cell_wire[1];							inform_R[2][1] = r_cell_wire[2];							inform_R[3][1] = r_cell_wire[3];							inform_R[4][1] = r_cell_wire[4];							inform_R[5][1] = r_cell_wire[5];							inform_R[6][1] = r_cell_wire[6];							inform_R[7][1] = r_cell_wire[7];							inform_R[8][1] = r_cell_wire[8];							inform_R[9][1] = r_cell_wire[9];							inform_R[10][1] = r_cell_wire[10];							inform_R[11][1] = r_cell_wire[11];							inform_R[12][1] = r_cell_wire[12];							inform_R[13][1] = r_cell_wire[13];							inform_R[14][1] = r_cell_wire[14];							inform_R[15][1] = r_cell_wire[15];							inform_R[16][1] = r_cell_wire[16];							inform_R[17][1] = r_cell_wire[17];							inform_R[18][1] = r_cell_wire[18];							inform_R[19][1] = r_cell_wire[19];							inform_R[20][1] = r_cell_wire[20];							inform_R[21][1] = r_cell_wire[21];							inform_R[22][1] = r_cell_wire[22];							inform_R[23][1] = r_cell_wire[23];							inform_R[24][1] = r_cell_wire[24];							inform_R[25][1] = r_cell_wire[25];							inform_R[26][1] = r_cell_wire[26];							inform_R[27][1] = r_cell_wire[27];							inform_R[28][1] = r_cell_wire[28];							inform_R[29][1] = r_cell_wire[29];							inform_R[30][1] = r_cell_wire[30];							inform_R[31][1] = r_cell_wire[31];							inform_R[32][1] = r_cell_wire[32];							inform_R[33][1] = r_cell_wire[33];							inform_R[34][1] = r_cell_wire[34];							inform_R[35][1] = r_cell_wire[35];							inform_R[36][1] = r_cell_wire[36];							inform_R[37][1] = r_cell_wire[37];							inform_R[38][1] = r_cell_wire[38];							inform_R[39][1] = r_cell_wire[39];							inform_R[40][1] = r_cell_wire[40];							inform_R[41][1] = r_cell_wire[41];							inform_R[42][1] = r_cell_wire[42];							inform_R[43][1] = r_cell_wire[43];							inform_R[44][1] = r_cell_wire[44];							inform_R[45][1] = r_cell_wire[45];							inform_R[46][1] = r_cell_wire[46];							inform_R[47][1] = r_cell_wire[47];							inform_R[48][1] = r_cell_wire[48];							inform_R[49][1] = r_cell_wire[49];							inform_R[50][1] = r_cell_wire[50];							inform_R[51][1] = r_cell_wire[51];							inform_R[52][1] = r_cell_wire[52];							inform_R[53][1] = r_cell_wire[53];							inform_R[54][1] = r_cell_wire[54];							inform_R[55][1] = r_cell_wire[55];							inform_R[56][1] = r_cell_wire[56];							inform_R[57][1] = r_cell_wire[57];							inform_R[58][1] = r_cell_wire[58];							inform_R[59][1] = r_cell_wire[59];							inform_R[60][1] = r_cell_wire[60];							inform_R[61][1] = r_cell_wire[61];							inform_R[62][1] = r_cell_wire[62];							inform_R[63][1] = r_cell_wire[63];							inform_R[64][1] = r_cell_wire[64];							inform_R[65][1] = r_cell_wire[65];							inform_R[66][1] = r_cell_wire[66];							inform_R[67][1] = r_cell_wire[67];							inform_R[68][1] = r_cell_wire[68];							inform_R[69][1] = r_cell_wire[69];							inform_R[70][1] = r_cell_wire[70];							inform_R[71][1] = r_cell_wire[71];							inform_R[72][1] = r_cell_wire[72];							inform_R[73][1] = r_cell_wire[73];							inform_R[74][1] = r_cell_wire[74];							inform_R[75][1] = r_cell_wire[75];							inform_R[76][1] = r_cell_wire[76];							inform_R[77][1] = r_cell_wire[77];							inform_R[78][1] = r_cell_wire[78];							inform_R[79][1] = r_cell_wire[79];							inform_R[80][1] = r_cell_wire[80];							inform_R[81][1] = r_cell_wire[81];							inform_R[82][1] = r_cell_wire[82];							inform_R[83][1] = r_cell_wire[83];							inform_R[84][1] = r_cell_wire[84];							inform_R[85][1] = r_cell_wire[85];							inform_R[86][1] = r_cell_wire[86];							inform_R[87][1] = r_cell_wire[87];							inform_R[88][1] = r_cell_wire[88];							inform_R[89][1] = r_cell_wire[89];							inform_R[90][1] = r_cell_wire[90];							inform_R[91][1] = r_cell_wire[91];							inform_R[92][1] = r_cell_wire[92];							inform_R[93][1] = r_cell_wire[93];							inform_R[94][1] = r_cell_wire[94];							inform_R[95][1] = r_cell_wire[95];							inform_R[96][1] = r_cell_wire[96];							inform_R[97][1] = r_cell_wire[97];							inform_R[98][1] = r_cell_wire[98];							inform_R[99][1] = r_cell_wire[99];							inform_R[100][1] = r_cell_wire[100];							inform_R[101][1] = r_cell_wire[101];							inform_R[102][1] = r_cell_wire[102];							inform_R[103][1] = r_cell_wire[103];							inform_R[104][1] = r_cell_wire[104];							inform_R[105][1] = r_cell_wire[105];							inform_R[106][1] = r_cell_wire[106];							inform_R[107][1] = r_cell_wire[107];							inform_R[108][1] = r_cell_wire[108];							inform_R[109][1] = r_cell_wire[109];							inform_R[110][1] = r_cell_wire[110];							inform_R[111][1] = r_cell_wire[111];							inform_R[112][1] = r_cell_wire[112];							inform_R[113][1] = r_cell_wire[113];							inform_R[114][1] = r_cell_wire[114];							inform_R[115][1] = r_cell_wire[115];							inform_R[116][1] = r_cell_wire[116];							inform_R[117][1] = r_cell_wire[117];							inform_R[118][1] = r_cell_wire[118];							inform_R[119][1] = r_cell_wire[119];							inform_R[120][1] = r_cell_wire[120];							inform_R[121][1] = r_cell_wire[121];							inform_R[122][1] = r_cell_wire[122];							inform_R[123][1] = r_cell_wire[123];							inform_R[124][1] = r_cell_wire[124];							inform_R[125][1] = r_cell_wire[125];							inform_R[126][1] = r_cell_wire[126];							inform_R[127][1] = r_cell_wire[127];							inform_L[0][0] = l_cell_wire[0];							inform_L[1][0] = l_cell_wire[1];							inform_L[2][0] = l_cell_wire[2];							inform_L[3][0] = l_cell_wire[3];							inform_L[4][0] = l_cell_wire[4];							inform_L[5][0] = l_cell_wire[5];							inform_L[6][0] = l_cell_wire[6];							inform_L[7][0] = l_cell_wire[7];							inform_L[8][0] = l_cell_wire[8];							inform_L[9][0] = l_cell_wire[9];							inform_L[10][0] = l_cell_wire[10];							inform_L[11][0] = l_cell_wire[11];							inform_L[12][0] = l_cell_wire[12];							inform_L[13][0] = l_cell_wire[13];							inform_L[14][0] = l_cell_wire[14];							inform_L[15][0] = l_cell_wire[15];							inform_L[16][0] = l_cell_wire[16];							inform_L[17][0] = l_cell_wire[17];							inform_L[18][0] = l_cell_wire[18];							inform_L[19][0] = l_cell_wire[19];							inform_L[20][0] = l_cell_wire[20];							inform_L[21][0] = l_cell_wire[21];							inform_L[22][0] = l_cell_wire[22];							inform_L[23][0] = l_cell_wire[23];							inform_L[24][0] = l_cell_wire[24];							inform_L[25][0] = l_cell_wire[25];							inform_L[26][0] = l_cell_wire[26];							inform_L[27][0] = l_cell_wire[27];							inform_L[28][0] = l_cell_wire[28];							inform_L[29][0] = l_cell_wire[29];							inform_L[30][0] = l_cell_wire[30];							inform_L[31][0] = l_cell_wire[31];							inform_L[32][0] = l_cell_wire[32];							inform_L[33][0] = l_cell_wire[33];							inform_L[34][0] = l_cell_wire[34];							inform_L[35][0] = l_cell_wire[35];							inform_L[36][0] = l_cell_wire[36];							inform_L[37][0] = l_cell_wire[37];							inform_L[38][0] = l_cell_wire[38];							inform_L[39][0] = l_cell_wire[39];							inform_L[40][0] = l_cell_wire[40];							inform_L[41][0] = l_cell_wire[41];							inform_L[42][0] = l_cell_wire[42];							inform_L[43][0] = l_cell_wire[43];							inform_L[44][0] = l_cell_wire[44];							inform_L[45][0] = l_cell_wire[45];							inform_L[46][0] = l_cell_wire[46];							inform_L[47][0] = l_cell_wire[47];							inform_L[48][0] = l_cell_wire[48];							inform_L[49][0] = l_cell_wire[49];							inform_L[50][0] = l_cell_wire[50];							inform_L[51][0] = l_cell_wire[51];							inform_L[52][0] = l_cell_wire[52];							inform_L[53][0] = l_cell_wire[53];							inform_L[54][0] = l_cell_wire[54];							inform_L[55][0] = l_cell_wire[55];							inform_L[56][0] = l_cell_wire[56];							inform_L[57][0] = l_cell_wire[57];							inform_L[58][0] = l_cell_wire[58];							inform_L[59][0] = l_cell_wire[59];							inform_L[60][0] = l_cell_wire[60];							inform_L[61][0] = l_cell_wire[61];							inform_L[62][0] = l_cell_wire[62];							inform_L[63][0] = l_cell_wire[63];							inform_L[64][0] = l_cell_wire[64];							inform_L[65][0] = l_cell_wire[65];							inform_L[66][0] = l_cell_wire[66];							inform_L[67][0] = l_cell_wire[67];							inform_L[68][0] = l_cell_wire[68];							inform_L[69][0] = l_cell_wire[69];							inform_L[70][0] = l_cell_wire[70];							inform_L[71][0] = l_cell_wire[71];							inform_L[72][0] = l_cell_wire[72];							inform_L[73][0] = l_cell_wire[73];							inform_L[74][0] = l_cell_wire[74];							inform_L[75][0] = l_cell_wire[75];							inform_L[76][0] = l_cell_wire[76];							inform_L[77][0] = l_cell_wire[77];							inform_L[78][0] = l_cell_wire[78];							inform_L[79][0] = l_cell_wire[79];							inform_L[80][0] = l_cell_wire[80];							inform_L[81][0] = l_cell_wire[81];							inform_L[82][0] = l_cell_wire[82];							inform_L[83][0] = l_cell_wire[83];							inform_L[84][0] = l_cell_wire[84];							inform_L[85][0] = l_cell_wire[85];							inform_L[86][0] = l_cell_wire[86];							inform_L[87][0] = l_cell_wire[87];							inform_L[88][0] = l_cell_wire[88];							inform_L[89][0] = l_cell_wire[89];							inform_L[90][0] = l_cell_wire[90];							inform_L[91][0] = l_cell_wire[91];							inform_L[92][0] = l_cell_wire[92];							inform_L[93][0] = l_cell_wire[93];							inform_L[94][0] = l_cell_wire[94];							inform_L[95][0] = l_cell_wire[95];							inform_L[96][0] = l_cell_wire[96];							inform_L[97][0] = l_cell_wire[97];							inform_L[98][0] = l_cell_wire[98];							inform_L[99][0] = l_cell_wire[99];							inform_L[100][0] = l_cell_wire[100];							inform_L[101][0] = l_cell_wire[101];							inform_L[102][0] = l_cell_wire[102];							inform_L[103][0] = l_cell_wire[103];							inform_L[104][0] = l_cell_wire[104];							inform_L[105][0] = l_cell_wire[105];							inform_L[106][0] = l_cell_wire[106];							inform_L[107][0] = l_cell_wire[107];							inform_L[108][0] = l_cell_wire[108];							inform_L[109][0] = l_cell_wire[109];							inform_L[110][0] = l_cell_wire[110];							inform_L[111][0] = l_cell_wire[111];							inform_L[112][0] = l_cell_wire[112];							inform_L[113][0] = l_cell_wire[113];							inform_L[114][0] = l_cell_wire[114];							inform_L[115][0] = l_cell_wire[115];							inform_L[116][0] = l_cell_wire[116];							inform_L[117][0] = l_cell_wire[117];							inform_L[118][0] = l_cell_wire[118];							inform_L[119][0] = l_cell_wire[119];							inform_L[120][0] = l_cell_wire[120];							inform_L[121][0] = l_cell_wire[121];							inform_L[122][0] = l_cell_wire[122];							inform_L[123][0] = l_cell_wire[123];							inform_L[124][0] = l_cell_wire[124];							inform_L[125][0] = l_cell_wire[125];							inform_L[126][0] = l_cell_wire[126];							inform_L[127][0] = l_cell_wire[127];						end
						2:						begin							inform_R[0][2] = r_cell_wire[0];							inform_R[2][2] = r_cell_wire[1];							inform_R[1][2] = r_cell_wire[2];							inform_R[3][2] = r_cell_wire[3];							inform_R[4][2] = r_cell_wire[4];							inform_R[6][2] = r_cell_wire[5];							inform_R[5][2] = r_cell_wire[6];							inform_R[7][2] = r_cell_wire[7];							inform_R[8][2] = r_cell_wire[8];							inform_R[10][2] = r_cell_wire[9];							inform_R[9][2] = r_cell_wire[10];							inform_R[11][2] = r_cell_wire[11];							inform_R[12][2] = r_cell_wire[12];							inform_R[14][2] = r_cell_wire[13];							inform_R[13][2] = r_cell_wire[14];							inform_R[15][2] = r_cell_wire[15];							inform_R[16][2] = r_cell_wire[16];							inform_R[18][2] = r_cell_wire[17];							inform_R[17][2] = r_cell_wire[18];							inform_R[19][2] = r_cell_wire[19];							inform_R[20][2] = r_cell_wire[20];							inform_R[22][2] = r_cell_wire[21];							inform_R[21][2] = r_cell_wire[22];							inform_R[23][2] = r_cell_wire[23];							inform_R[24][2] = r_cell_wire[24];							inform_R[26][2] = r_cell_wire[25];							inform_R[25][2] = r_cell_wire[26];							inform_R[27][2] = r_cell_wire[27];							inform_R[28][2] = r_cell_wire[28];							inform_R[30][2] = r_cell_wire[29];							inform_R[29][2] = r_cell_wire[30];							inform_R[31][2] = r_cell_wire[31];							inform_R[32][2] = r_cell_wire[32];							inform_R[34][2] = r_cell_wire[33];							inform_R[33][2] = r_cell_wire[34];							inform_R[35][2] = r_cell_wire[35];							inform_R[36][2] = r_cell_wire[36];							inform_R[38][2] = r_cell_wire[37];							inform_R[37][2] = r_cell_wire[38];							inform_R[39][2] = r_cell_wire[39];							inform_R[40][2] = r_cell_wire[40];							inform_R[42][2] = r_cell_wire[41];							inform_R[41][2] = r_cell_wire[42];							inform_R[43][2] = r_cell_wire[43];							inform_R[44][2] = r_cell_wire[44];							inform_R[46][2] = r_cell_wire[45];							inform_R[45][2] = r_cell_wire[46];							inform_R[47][2] = r_cell_wire[47];							inform_R[48][2] = r_cell_wire[48];							inform_R[50][2] = r_cell_wire[49];							inform_R[49][2] = r_cell_wire[50];							inform_R[51][2] = r_cell_wire[51];							inform_R[52][2] = r_cell_wire[52];							inform_R[54][2] = r_cell_wire[53];							inform_R[53][2] = r_cell_wire[54];							inform_R[55][2] = r_cell_wire[55];							inform_R[56][2] = r_cell_wire[56];							inform_R[58][2] = r_cell_wire[57];							inform_R[57][2] = r_cell_wire[58];							inform_R[59][2] = r_cell_wire[59];							inform_R[60][2] = r_cell_wire[60];							inform_R[62][2] = r_cell_wire[61];							inform_R[61][2] = r_cell_wire[62];							inform_R[63][2] = r_cell_wire[63];							inform_R[64][2] = r_cell_wire[64];							inform_R[66][2] = r_cell_wire[65];							inform_R[65][2] = r_cell_wire[66];							inform_R[67][2] = r_cell_wire[67];							inform_R[68][2] = r_cell_wire[68];							inform_R[70][2] = r_cell_wire[69];							inform_R[69][2] = r_cell_wire[70];							inform_R[71][2] = r_cell_wire[71];							inform_R[72][2] = r_cell_wire[72];							inform_R[74][2] = r_cell_wire[73];							inform_R[73][2] = r_cell_wire[74];							inform_R[75][2] = r_cell_wire[75];							inform_R[76][2] = r_cell_wire[76];							inform_R[78][2] = r_cell_wire[77];							inform_R[77][2] = r_cell_wire[78];							inform_R[79][2] = r_cell_wire[79];							inform_R[80][2] = r_cell_wire[80];							inform_R[82][2] = r_cell_wire[81];							inform_R[81][2] = r_cell_wire[82];							inform_R[83][2] = r_cell_wire[83];							inform_R[84][2] = r_cell_wire[84];							inform_R[86][2] = r_cell_wire[85];							inform_R[85][2] = r_cell_wire[86];							inform_R[87][2] = r_cell_wire[87];							inform_R[88][2] = r_cell_wire[88];							inform_R[90][2] = r_cell_wire[89];							inform_R[89][2] = r_cell_wire[90];							inform_R[91][2] = r_cell_wire[91];							inform_R[92][2] = r_cell_wire[92];							inform_R[94][2] = r_cell_wire[93];							inform_R[93][2] = r_cell_wire[94];							inform_R[95][2] = r_cell_wire[95];							inform_R[96][2] = r_cell_wire[96];							inform_R[98][2] = r_cell_wire[97];							inform_R[97][2] = r_cell_wire[98];							inform_R[99][2] = r_cell_wire[99];							inform_R[100][2] = r_cell_wire[100];							inform_R[102][2] = r_cell_wire[101];							inform_R[101][2] = r_cell_wire[102];							inform_R[103][2] = r_cell_wire[103];							inform_R[104][2] = r_cell_wire[104];							inform_R[106][2] = r_cell_wire[105];							inform_R[105][2] = r_cell_wire[106];							inform_R[107][2] = r_cell_wire[107];							inform_R[108][2] = r_cell_wire[108];							inform_R[110][2] = r_cell_wire[109];							inform_R[109][2] = r_cell_wire[110];							inform_R[111][2] = r_cell_wire[111];							inform_R[112][2] = r_cell_wire[112];							inform_R[114][2] = r_cell_wire[113];							inform_R[113][2] = r_cell_wire[114];							inform_R[115][2] = r_cell_wire[115];							inform_R[116][2] = r_cell_wire[116];							inform_R[118][2] = r_cell_wire[117];							inform_R[117][2] = r_cell_wire[118];							inform_R[119][2] = r_cell_wire[119];							inform_R[120][2] = r_cell_wire[120];							inform_R[122][2] = r_cell_wire[121];							inform_R[121][2] = r_cell_wire[122];							inform_R[123][2] = r_cell_wire[123];							inform_R[124][2] = r_cell_wire[124];							inform_R[126][2] = r_cell_wire[125];							inform_R[125][2] = r_cell_wire[126];							inform_R[127][2] = r_cell_wire[127];							inform_L[0][1] = l_cell_wire[0];							inform_L[2][1] = l_cell_wire[1];							inform_L[1][1] = l_cell_wire[2];							inform_L[3][1] = l_cell_wire[3];							inform_L[4][1] = l_cell_wire[4];							inform_L[6][1] = l_cell_wire[5];							inform_L[5][1] = l_cell_wire[6];							inform_L[7][1] = l_cell_wire[7];							inform_L[8][1] = l_cell_wire[8];							inform_L[10][1] = l_cell_wire[9];							inform_L[9][1] = l_cell_wire[10];							inform_L[11][1] = l_cell_wire[11];							inform_L[12][1] = l_cell_wire[12];							inform_L[14][1] = l_cell_wire[13];							inform_L[13][1] = l_cell_wire[14];							inform_L[15][1] = l_cell_wire[15];							inform_L[16][1] = l_cell_wire[16];							inform_L[18][1] = l_cell_wire[17];							inform_L[17][1] = l_cell_wire[18];							inform_L[19][1] = l_cell_wire[19];							inform_L[20][1] = l_cell_wire[20];							inform_L[22][1] = l_cell_wire[21];							inform_L[21][1] = l_cell_wire[22];							inform_L[23][1] = l_cell_wire[23];							inform_L[24][1] = l_cell_wire[24];							inform_L[26][1] = l_cell_wire[25];							inform_L[25][1] = l_cell_wire[26];							inform_L[27][1] = l_cell_wire[27];							inform_L[28][1] = l_cell_wire[28];							inform_L[30][1] = l_cell_wire[29];							inform_L[29][1] = l_cell_wire[30];							inform_L[31][1] = l_cell_wire[31];							inform_L[32][1] = l_cell_wire[32];							inform_L[34][1] = l_cell_wire[33];							inform_L[33][1] = l_cell_wire[34];							inform_L[35][1] = l_cell_wire[35];							inform_L[36][1] = l_cell_wire[36];							inform_L[38][1] = l_cell_wire[37];							inform_L[37][1] = l_cell_wire[38];							inform_L[39][1] = l_cell_wire[39];							inform_L[40][1] = l_cell_wire[40];							inform_L[42][1] = l_cell_wire[41];							inform_L[41][1] = l_cell_wire[42];							inform_L[43][1] = l_cell_wire[43];							inform_L[44][1] = l_cell_wire[44];							inform_L[46][1] = l_cell_wire[45];							inform_L[45][1] = l_cell_wire[46];							inform_L[47][1] = l_cell_wire[47];							inform_L[48][1] = l_cell_wire[48];							inform_L[50][1] = l_cell_wire[49];							inform_L[49][1] = l_cell_wire[50];							inform_L[51][1] = l_cell_wire[51];							inform_L[52][1] = l_cell_wire[52];							inform_L[54][1] = l_cell_wire[53];							inform_L[53][1] = l_cell_wire[54];							inform_L[55][1] = l_cell_wire[55];							inform_L[56][1] = l_cell_wire[56];							inform_L[58][1] = l_cell_wire[57];							inform_L[57][1] = l_cell_wire[58];							inform_L[59][1] = l_cell_wire[59];							inform_L[60][1] = l_cell_wire[60];							inform_L[62][1] = l_cell_wire[61];							inform_L[61][1] = l_cell_wire[62];							inform_L[63][1] = l_cell_wire[63];							inform_L[64][1] = l_cell_wire[64];							inform_L[66][1] = l_cell_wire[65];							inform_L[65][1] = l_cell_wire[66];							inform_L[67][1] = l_cell_wire[67];							inform_L[68][1] = l_cell_wire[68];							inform_L[70][1] = l_cell_wire[69];							inform_L[69][1] = l_cell_wire[70];							inform_L[71][1] = l_cell_wire[71];							inform_L[72][1] = l_cell_wire[72];							inform_L[74][1] = l_cell_wire[73];							inform_L[73][1] = l_cell_wire[74];							inform_L[75][1] = l_cell_wire[75];							inform_L[76][1] = l_cell_wire[76];							inform_L[78][1] = l_cell_wire[77];							inform_L[77][1] = l_cell_wire[78];							inform_L[79][1] = l_cell_wire[79];							inform_L[80][1] = l_cell_wire[80];							inform_L[82][1] = l_cell_wire[81];							inform_L[81][1] = l_cell_wire[82];							inform_L[83][1] = l_cell_wire[83];							inform_L[84][1] = l_cell_wire[84];							inform_L[86][1] = l_cell_wire[85];							inform_L[85][1] = l_cell_wire[86];							inform_L[87][1] = l_cell_wire[87];							inform_L[88][1] = l_cell_wire[88];							inform_L[90][1] = l_cell_wire[89];							inform_L[89][1] = l_cell_wire[90];							inform_L[91][1] = l_cell_wire[91];							inform_L[92][1] = l_cell_wire[92];							inform_L[94][1] = l_cell_wire[93];							inform_L[93][1] = l_cell_wire[94];							inform_L[95][1] = l_cell_wire[95];							inform_L[96][1] = l_cell_wire[96];							inform_L[98][1] = l_cell_wire[97];							inform_L[97][1] = l_cell_wire[98];							inform_L[99][1] = l_cell_wire[99];							inform_L[100][1] = l_cell_wire[100];							inform_L[102][1] = l_cell_wire[101];							inform_L[101][1] = l_cell_wire[102];							inform_L[103][1] = l_cell_wire[103];							inform_L[104][1] = l_cell_wire[104];							inform_L[106][1] = l_cell_wire[105];							inform_L[105][1] = l_cell_wire[106];							inform_L[107][1] = l_cell_wire[107];							inform_L[108][1] = l_cell_wire[108];							inform_L[110][1] = l_cell_wire[109];							inform_L[109][1] = l_cell_wire[110];							inform_L[111][1] = l_cell_wire[111];							inform_L[112][1] = l_cell_wire[112];							inform_L[114][1] = l_cell_wire[113];							inform_L[113][1] = l_cell_wire[114];							inform_L[115][1] = l_cell_wire[115];							inform_L[116][1] = l_cell_wire[116];							inform_L[118][1] = l_cell_wire[117];							inform_L[117][1] = l_cell_wire[118];							inform_L[119][1] = l_cell_wire[119];							inform_L[120][1] = l_cell_wire[120];							inform_L[122][1] = l_cell_wire[121];							inform_L[121][1] = l_cell_wire[122];							inform_L[123][1] = l_cell_wire[123];							inform_L[124][1] = l_cell_wire[124];							inform_L[126][1] = l_cell_wire[125];							inform_L[125][1] = l_cell_wire[126];							inform_L[127][1] = l_cell_wire[127];						end
						3:						begin							inform_R[0][3] = r_cell_wire[0];							inform_R[4][3] = r_cell_wire[1];							inform_R[1][3] = r_cell_wire[2];							inform_R[5][3] = r_cell_wire[3];							inform_R[2][3] = r_cell_wire[4];							inform_R[6][3] = r_cell_wire[5];							inform_R[3][3] = r_cell_wire[6];							inform_R[7][3] = r_cell_wire[7];							inform_R[8][3] = r_cell_wire[8];							inform_R[12][3] = r_cell_wire[9];							inform_R[9][3] = r_cell_wire[10];							inform_R[13][3] = r_cell_wire[11];							inform_R[10][3] = r_cell_wire[12];							inform_R[14][3] = r_cell_wire[13];							inform_R[11][3] = r_cell_wire[14];							inform_R[15][3] = r_cell_wire[15];							inform_R[16][3] = r_cell_wire[16];							inform_R[20][3] = r_cell_wire[17];							inform_R[17][3] = r_cell_wire[18];							inform_R[21][3] = r_cell_wire[19];							inform_R[18][3] = r_cell_wire[20];							inform_R[22][3] = r_cell_wire[21];							inform_R[19][3] = r_cell_wire[22];							inform_R[23][3] = r_cell_wire[23];							inform_R[24][3] = r_cell_wire[24];							inform_R[28][3] = r_cell_wire[25];							inform_R[25][3] = r_cell_wire[26];							inform_R[29][3] = r_cell_wire[27];							inform_R[26][3] = r_cell_wire[28];							inform_R[30][3] = r_cell_wire[29];							inform_R[27][3] = r_cell_wire[30];							inform_R[31][3] = r_cell_wire[31];							inform_R[32][3] = r_cell_wire[32];							inform_R[36][3] = r_cell_wire[33];							inform_R[33][3] = r_cell_wire[34];							inform_R[37][3] = r_cell_wire[35];							inform_R[34][3] = r_cell_wire[36];							inform_R[38][3] = r_cell_wire[37];							inform_R[35][3] = r_cell_wire[38];							inform_R[39][3] = r_cell_wire[39];							inform_R[40][3] = r_cell_wire[40];							inform_R[44][3] = r_cell_wire[41];							inform_R[41][3] = r_cell_wire[42];							inform_R[45][3] = r_cell_wire[43];							inform_R[42][3] = r_cell_wire[44];							inform_R[46][3] = r_cell_wire[45];							inform_R[43][3] = r_cell_wire[46];							inform_R[47][3] = r_cell_wire[47];							inform_R[48][3] = r_cell_wire[48];							inform_R[52][3] = r_cell_wire[49];							inform_R[49][3] = r_cell_wire[50];							inform_R[53][3] = r_cell_wire[51];							inform_R[50][3] = r_cell_wire[52];							inform_R[54][3] = r_cell_wire[53];							inform_R[51][3] = r_cell_wire[54];							inform_R[55][3] = r_cell_wire[55];							inform_R[56][3] = r_cell_wire[56];							inform_R[60][3] = r_cell_wire[57];							inform_R[57][3] = r_cell_wire[58];							inform_R[61][3] = r_cell_wire[59];							inform_R[58][3] = r_cell_wire[60];							inform_R[62][3] = r_cell_wire[61];							inform_R[59][3] = r_cell_wire[62];							inform_R[63][3] = r_cell_wire[63];							inform_R[64][3] = r_cell_wire[64];							inform_R[68][3] = r_cell_wire[65];							inform_R[65][3] = r_cell_wire[66];							inform_R[69][3] = r_cell_wire[67];							inform_R[66][3] = r_cell_wire[68];							inform_R[70][3] = r_cell_wire[69];							inform_R[67][3] = r_cell_wire[70];							inform_R[71][3] = r_cell_wire[71];							inform_R[72][3] = r_cell_wire[72];							inform_R[76][3] = r_cell_wire[73];							inform_R[73][3] = r_cell_wire[74];							inform_R[77][3] = r_cell_wire[75];							inform_R[74][3] = r_cell_wire[76];							inform_R[78][3] = r_cell_wire[77];							inform_R[75][3] = r_cell_wire[78];							inform_R[79][3] = r_cell_wire[79];							inform_R[80][3] = r_cell_wire[80];							inform_R[84][3] = r_cell_wire[81];							inform_R[81][3] = r_cell_wire[82];							inform_R[85][3] = r_cell_wire[83];							inform_R[82][3] = r_cell_wire[84];							inform_R[86][3] = r_cell_wire[85];							inform_R[83][3] = r_cell_wire[86];							inform_R[87][3] = r_cell_wire[87];							inform_R[88][3] = r_cell_wire[88];							inform_R[92][3] = r_cell_wire[89];							inform_R[89][3] = r_cell_wire[90];							inform_R[93][3] = r_cell_wire[91];							inform_R[90][3] = r_cell_wire[92];							inform_R[94][3] = r_cell_wire[93];							inform_R[91][3] = r_cell_wire[94];							inform_R[95][3] = r_cell_wire[95];							inform_R[96][3] = r_cell_wire[96];							inform_R[100][3] = r_cell_wire[97];							inform_R[97][3] = r_cell_wire[98];							inform_R[101][3] = r_cell_wire[99];							inform_R[98][3] = r_cell_wire[100];							inform_R[102][3] = r_cell_wire[101];							inform_R[99][3] = r_cell_wire[102];							inform_R[103][3] = r_cell_wire[103];							inform_R[104][3] = r_cell_wire[104];							inform_R[108][3] = r_cell_wire[105];							inform_R[105][3] = r_cell_wire[106];							inform_R[109][3] = r_cell_wire[107];							inform_R[106][3] = r_cell_wire[108];							inform_R[110][3] = r_cell_wire[109];							inform_R[107][3] = r_cell_wire[110];							inform_R[111][3] = r_cell_wire[111];							inform_R[112][3] = r_cell_wire[112];							inform_R[116][3] = r_cell_wire[113];							inform_R[113][3] = r_cell_wire[114];							inform_R[117][3] = r_cell_wire[115];							inform_R[114][3] = r_cell_wire[116];							inform_R[118][3] = r_cell_wire[117];							inform_R[115][3] = r_cell_wire[118];							inform_R[119][3] = r_cell_wire[119];							inform_R[120][3] = r_cell_wire[120];							inform_R[124][3] = r_cell_wire[121];							inform_R[121][3] = r_cell_wire[122];							inform_R[125][3] = r_cell_wire[123];							inform_R[122][3] = r_cell_wire[124];							inform_R[126][3] = r_cell_wire[125];							inform_R[123][3] = r_cell_wire[126];							inform_R[127][3] = r_cell_wire[127];							inform_L[0][2] = l_cell_wire[0];							inform_L[4][2] = l_cell_wire[1];							inform_L[1][2] = l_cell_wire[2];							inform_L[5][2] = l_cell_wire[3];							inform_L[2][2] = l_cell_wire[4];							inform_L[6][2] = l_cell_wire[5];							inform_L[3][2] = l_cell_wire[6];							inform_L[7][2] = l_cell_wire[7];							inform_L[8][2] = l_cell_wire[8];							inform_L[12][2] = l_cell_wire[9];							inform_L[9][2] = l_cell_wire[10];							inform_L[13][2] = l_cell_wire[11];							inform_L[10][2] = l_cell_wire[12];							inform_L[14][2] = l_cell_wire[13];							inform_L[11][2] = l_cell_wire[14];							inform_L[15][2] = l_cell_wire[15];							inform_L[16][2] = l_cell_wire[16];							inform_L[20][2] = l_cell_wire[17];							inform_L[17][2] = l_cell_wire[18];							inform_L[21][2] = l_cell_wire[19];							inform_L[18][2] = l_cell_wire[20];							inform_L[22][2] = l_cell_wire[21];							inform_L[19][2] = l_cell_wire[22];							inform_L[23][2] = l_cell_wire[23];							inform_L[24][2] = l_cell_wire[24];							inform_L[28][2] = l_cell_wire[25];							inform_L[25][2] = l_cell_wire[26];							inform_L[29][2] = l_cell_wire[27];							inform_L[26][2] = l_cell_wire[28];							inform_L[30][2] = l_cell_wire[29];							inform_L[27][2] = l_cell_wire[30];							inform_L[31][2] = l_cell_wire[31];							inform_L[32][2] = l_cell_wire[32];							inform_L[36][2] = l_cell_wire[33];							inform_L[33][2] = l_cell_wire[34];							inform_L[37][2] = l_cell_wire[35];							inform_L[34][2] = l_cell_wire[36];							inform_L[38][2] = l_cell_wire[37];							inform_L[35][2] = l_cell_wire[38];							inform_L[39][2] = l_cell_wire[39];							inform_L[40][2] = l_cell_wire[40];							inform_L[44][2] = l_cell_wire[41];							inform_L[41][2] = l_cell_wire[42];							inform_L[45][2] = l_cell_wire[43];							inform_L[42][2] = l_cell_wire[44];							inform_L[46][2] = l_cell_wire[45];							inform_L[43][2] = l_cell_wire[46];							inform_L[47][2] = l_cell_wire[47];							inform_L[48][2] = l_cell_wire[48];							inform_L[52][2] = l_cell_wire[49];							inform_L[49][2] = l_cell_wire[50];							inform_L[53][2] = l_cell_wire[51];							inform_L[50][2] = l_cell_wire[52];							inform_L[54][2] = l_cell_wire[53];							inform_L[51][2] = l_cell_wire[54];							inform_L[55][2] = l_cell_wire[55];							inform_L[56][2] = l_cell_wire[56];							inform_L[60][2] = l_cell_wire[57];							inform_L[57][2] = l_cell_wire[58];							inform_L[61][2] = l_cell_wire[59];							inform_L[58][2] = l_cell_wire[60];							inform_L[62][2] = l_cell_wire[61];							inform_L[59][2] = l_cell_wire[62];							inform_L[63][2] = l_cell_wire[63];							inform_L[64][2] = l_cell_wire[64];							inform_L[68][2] = l_cell_wire[65];							inform_L[65][2] = l_cell_wire[66];							inform_L[69][2] = l_cell_wire[67];							inform_L[66][2] = l_cell_wire[68];							inform_L[70][2] = l_cell_wire[69];							inform_L[67][2] = l_cell_wire[70];							inform_L[71][2] = l_cell_wire[71];							inform_L[72][2] = l_cell_wire[72];							inform_L[76][2] = l_cell_wire[73];							inform_L[73][2] = l_cell_wire[74];							inform_L[77][2] = l_cell_wire[75];							inform_L[74][2] = l_cell_wire[76];							inform_L[78][2] = l_cell_wire[77];							inform_L[75][2] = l_cell_wire[78];							inform_L[79][2] = l_cell_wire[79];							inform_L[80][2] = l_cell_wire[80];							inform_L[84][2] = l_cell_wire[81];							inform_L[81][2] = l_cell_wire[82];							inform_L[85][2] = l_cell_wire[83];							inform_L[82][2] = l_cell_wire[84];							inform_L[86][2] = l_cell_wire[85];							inform_L[83][2] = l_cell_wire[86];							inform_L[87][2] = l_cell_wire[87];							inform_L[88][2] = l_cell_wire[88];							inform_L[92][2] = l_cell_wire[89];							inform_L[89][2] = l_cell_wire[90];							inform_L[93][2] = l_cell_wire[91];							inform_L[90][2] = l_cell_wire[92];							inform_L[94][2] = l_cell_wire[93];							inform_L[91][2] = l_cell_wire[94];							inform_L[95][2] = l_cell_wire[95];							inform_L[96][2] = l_cell_wire[96];							inform_L[100][2] = l_cell_wire[97];							inform_L[97][2] = l_cell_wire[98];							inform_L[101][2] = l_cell_wire[99];							inform_L[98][2] = l_cell_wire[100];							inform_L[102][2] = l_cell_wire[101];							inform_L[99][2] = l_cell_wire[102];							inform_L[103][2] = l_cell_wire[103];							inform_L[104][2] = l_cell_wire[104];							inform_L[108][2] = l_cell_wire[105];							inform_L[105][2] = l_cell_wire[106];							inform_L[109][2] = l_cell_wire[107];							inform_L[106][2] = l_cell_wire[108];							inform_L[110][2] = l_cell_wire[109];							inform_L[107][2] = l_cell_wire[110];							inform_L[111][2] = l_cell_wire[111];							inform_L[112][2] = l_cell_wire[112];							inform_L[116][2] = l_cell_wire[113];							inform_L[113][2] = l_cell_wire[114];							inform_L[117][2] = l_cell_wire[115];							inform_L[114][2] = l_cell_wire[116];							inform_L[118][2] = l_cell_wire[117];							inform_L[115][2] = l_cell_wire[118];							inform_L[119][2] = l_cell_wire[119];							inform_L[120][2] = l_cell_wire[120];							inform_L[124][2] = l_cell_wire[121];							inform_L[121][2] = l_cell_wire[122];							inform_L[125][2] = l_cell_wire[123];							inform_L[122][2] = l_cell_wire[124];							inform_L[126][2] = l_cell_wire[125];							inform_L[123][2] = l_cell_wire[126];							inform_L[127][2] = l_cell_wire[127];						end
						4:						begin							inform_R[0][4] = r_cell_wire[0];							inform_R[8][4] = r_cell_wire[1];							inform_R[1][4] = r_cell_wire[2];							inform_R[9][4] = r_cell_wire[3];							inform_R[2][4] = r_cell_wire[4];							inform_R[10][4] = r_cell_wire[5];							inform_R[3][4] = r_cell_wire[6];							inform_R[11][4] = r_cell_wire[7];							inform_R[4][4] = r_cell_wire[8];							inform_R[12][4] = r_cell_wire[9];							inform_R[5][4] = r_cell_wire[10];							inform_R[13][4] = r_cell_wire[11];							inform_R[6][4] = r_cell_wire[12];							inform_R[14][4] = r_cell_wire[13];							inform_R[7][4] = r_cell_wire[14];							inform_R[15][4] = r_cell_wire[15];							inform_R[16][4] = r_cell_wire[16];							inform_R[24][4] = r_cell_wire[17];							inform_R[17][4] = r_cell_wire[18];							inform_R[25][4] = r_cell_wire[19];							inform_R[18][4] = r_cell_wire[20];							inform_R[26][4] = r_cell_wire[21];							inform_R[19][4] = r_cell_wire[22];							inform_R[27][4] = r_cell_wire[23];							inform_R[20][4] = r_cell_wire[24];							inform_R[28][4] = r_cell_wire[25];							inform_R[21][4] = r_cell_wire[26];							inform_R[29][4] = r_cell_wire[27];							inform_R[22][4] = r_cell_wire[28];							inform_R[30][4] = r_cell_wire[29];							inform_R[23][4] = r_cell_wire[30];							inform_R[31][4] = r_cell_wire[31];							inform_R[32][4] = r_cell_wire[32];							inform_R[40][4] = r_cell_wire[33];							inform_R[33][4] = r_cell_wire[34];							inform_R[41][4] = r_cell_wire[35];							inform_R[34][4] = r_cell_wire[36];							inform_R[42][4] = r_cell_wire[37];							inform_R[35][4] = r_cell_wire[38];							inform_R[43][4] = r_cell_wire[39];							inform_R[36][4] = r_cell_wire[40];							inform_R[44][4] = r_cell_wire[41];							inform_R[37][4] = r_cell_wire[42];							inform_R[45][4] = r_cell_wire[43];							inform_R[38][4] = r_cell_wire[44];							inform_R[46][4] = r_cell_wire[45];							inform_R[39][4] = r_cell_wire[46];							inform_R[47][4] = r_cell_wire[47];							inform_R[48][4] = r_cell_wire[48];							inform_R[56][4] = r_cell_wire[49];							inform_R[49][4] = r_cell_wire[50];							inform_R[57][4] = r_cell_wire[51];							inform_R[50][4] = r_cell_wire[52];							inform_R[58][4] = r_cell_wire[53];							inform_R[51][4] = r_cell_wire[54];							inform_R[59][4] = r_cell_wire[55];							inform_R[52][4] = r_cell_wire[56];							inform_R[60][4] = r_cell_wire[57];							inform_R[53][4] = r_cell_wire[58];							inform_R[61][4] = r_cell_wire[59];							inform_R[54][4] = r_cell_wire[60];							inform_R[62][4] = r_cell_wire[61];							inform_R[55][4] = r_cell_wire[62];							inform_R[63][4] = r_cell_wire[63];							inform_R[64][4] = r_cell_wire[64];							inform_R[72][4] = r_cell_wire[65];							inform_R[65][4] = r_cell_wire[66];							inform_R[73][4] = r_cell_wire[67];							inform_R[66][4] = r_cell_wire[68];							inform_R[74][4] = r_cell_wire[69];							inform_R[67][4] = r_cell_wire[70];							inform_R[75][4] = r_cell_wire[71];							inform_R[68][4] = r_cell_wire[72];							inform_R[76][4] = r_cell_wire[73];							inform_R[69][4] = r_cell_wire[74];							inform_R[77][4] = r_cell_wire[75];							inform_R[70][4] = r_cell_wire[76];							inform_R[78][4] = r_cell_wire[77];							inform_R[71][4] = r_cell_wire[78];							inform_R[79][4] = r_cell_wire[79];							inform_R[80][4] = r_cell_wire[80];							inform_R[88][4] = r_cell_wire[81];							inform_R[81][4] = r_cell_wire[82];							inform_R[89][4] = r_cell_wire[83];							inform_R[82][4] = r_cell_wire[84];							inform_R[90][4] = r_cell_wire[85];							inform_R[83][4] = r_cell_wire[86];							inform_R[91][4] = r_cell_wire[87];							inform_R[84][4] = r_cell_wire[88];							inform_R[92][4] = r_cell_wire[89];							inform_R[85][4] = r_cell_wire[90];							inform_R[93][4] = r_cell_wire[91];							inform_R[86][4] = r_cell_wire[92];							inform_R[94][4] = r_cell_wire[93];							inform_R[87][4] = r_cell_wire[94];							inform_R[95][4] = r_cell_wire[95];							inform_R[96][4] = r_cell_wire[96];							inform_R[104][4] = r_cell_wire[97];							inform_R[97][4] = r_cell_wire[98];							inform_R[105][4] = r_cell_wire[99];							inform_R[98][4] = r_cell_wire[100];							inform_R[106][4] = r_cell_wire[101];							inform_R[99][4] = r_cell_wire[102];							inform_R[107][4] = r_cell_wire[103];							inform_R[100][4] = r_cell_wire[104];							inform_R[108][4] = r_cell_wire[105];							inform_R[101][4] = r_cell_wire[106];							inform_R[109][4] = r_cell_wire[107];							inform_R[102][4] = r_cell_wire[108];							inform_R[110][4] = r_cell_wire[109];							inform_R[103][4] = r_cell_wire[110];							inform_R[111][4] = r_cell_wire[111];							inform_R[112][4] = r_cell_wire[112];							inform_R[120][4] = r_cell_wire[113];							inform_R[113][4] = r_cell_wire[114];							inform_R[121][4] = r_cell_wire[115];							inform_R[114][4] = r_cell_wire[116];							inform_R[122][4] = r_cell_wire[117];							inform_R[115][4] = r_cell_wire[118];							inform_R[123][4] = r_cell_wire[119];							inform_R[116][4] = r_cell_wire[120];							inform_R[124][4] = r_cell_wire[121];							inform_R[117][4] = r_cell_wire[122];							inform_R[125][4] = r_cell_wire[123];							inform_R[118][4] = r_cell_wire[124];							inform_R[126][4] = r_cell_wire[125];							inform_R[119][4] = r_cell_wire[126];							inform_R[127][4] = r_cell_wire[127];							inform_L[0][3] = l_cell_wire[0];							inform_L[8][3] = l_cell_wire[1];							inform_L[1][3] = l_cell_wire[2];							inform_L[9][3] = l_cell_wire[3];							inform_L[2][3] = l_cell_wire[4];							inform_L[10][3] = l_cell_wire[5];							inform_L[3][3] = l_cell_wire[6];							inform_L[11][3] = l_cell_wire[7];							inform_L[4][3] = l_cell_wire[8];							inform_L[12][3] = l_cell_wire[9];							inform_L[5][3] = l_cell_wire[10];							inform_L[13][3] = l_cell_wire[11];							inform_L[6][3] = l_cell_wire[12];							inform_L[14][3] = l_cell_wire[13];							inform_L[7][3] = l_cell_wire[14];							inform_L[15][3] = l_cell_wire[15];							inform_L[16][3] = l_cell_wire[16];							inform_L[24][3] = l_cell_wire[17];							inform_L[17][3] = l_cell_wire[18];							inform_L[25][3] = l_cell_wire[19];							inform_L[18][3] = l_cell_wire[20];							inform_L[26][3] = l_cell_wire[21];							inform_L[19][3] = l_cell_wire[22];							inform_L[27][3] = l_cell_wire[23];							inform_L[20][3] = l_cell_wire[24];							inform_L[28][3] = l_cell_wire[25];							inform_L[21][3] = l_cell_wire[26];							inform_L[29][3] = l_cell_wire[27];							inform_L[22][3] = l_cell_wire[28];							inform_L[30][3] = l_cell_wire[29];							inform_L[23][3] = l_cell_wire[30];							inform_L[31][3] = l_cell_wire[31];							inform_L[32][3] = l_cell_wire[32];							inform_L[40][3] = l_cell_wire[33];							inform_L[33][3] = l_cell_wire[34];							inform_L[41][3] = l_cell_wire[35];							inform_L[34][3] = l_cell_wire[36];							inform_L[42][3] = l_cell_wire[37];							inform_L[35][3] = l_cell_wire[38];							inform_L[43][3] = l_cell_wire[39];							inform_L[36][3] = l_cell_wire[40];							inform_L[44][3] = l_cell_wire[41];							inform_L[37][3] = l_cell_wire[42];							inform_L[45][3] = l_cell_wire[43];							inform_L[38][3] = l_cell_wire[44];							inform_L[46][3] = l_cell_wire[45];							inform_L[39][3] = l_cell_wire[46];							inform_L[47][3] = l_cell_wire[47];							inform_L[48][3] = l_cell_wire[48];							inform_L[56][3] = l_cell_wire[49];							inform_L[49][3] = l_cell_wire[50];							inform_L[57][3] = l_cell_wire[51];							inform_L[50][3] = l_cell_wire[52];							inform_L[58][3] = l_cell_wire[53];							inform_L[51][3] = l_cell_wire[54];							inform_L[59][3] = l_cell_wire[55];							inform_L[52][3] = l_cell_wire[56];							inform_L[60][3] = l_cell_wire[57];							inform_L[53][3] = l_cell_wire[58];							inform_L[61][3] = l_cell_wire[59];							inform_L[54][3] = l_cell_wire[60];							inform_L[62][3] = l_cell_wire[61];							inform_L[55][3] = l_cell_wire[62];							inform_L[63][3] = l_cell_wire[63];							inform_L[64][3] = l_cell_wire[64];							inform_L[72][3] = l_cell_wire[65];							inform_L[65][3] = l_cell_wire[66];							inform_L[73][3] = l_cell_wire[67];							inform_L[66][3] = l_cell_wire[68];							inform_L[74][3] = l_cell_wire[69];							inform_L[67][3] = l_cell_wire[70];							inform_L[75][3] = l_cell_wire[71];							inform_L[68][3] = l_cell_wire[72];							inform_L[76][3] = l_cell_wire[73];							inform_L[69][3] = l_cell_wire[74];							inform_L[77][3] = l_cell_wire[75];							inform_L[70][3] = l_cell_wire[76];							inform_L[78][3] = l_cell_wire[77];							inform_L[71][3] = l_cell_wire[78];							inform_L[79][3] = l_cell_wire[79];							inform_L[80][3] = l_cell_wire[80];							inform_L[88][3] = l_cell_wire[81];							inform_L[81][3] = l_cell_wire[82];							inform_L[89][3] = l_cell_wire[83];							inform_L[82][3] = l_cell_wire[84];							inform_L[90][3] = l_cell_wire[85];							inform_L[83][3] = l_cell_wire[86];							inform_L[91][3] = l_cell_wire[87];							inform_L[84][3] = l_cell_wire[88];							inform_L[92][3] = l_cell_wire[89];							inform_L[85][3] = l_cell_wire[90];							inform_L[93][3] = l_cell_wire[91];							inform_L[86][3] = l_cell_wire[92];							inform_L[94][3] = l_cell_wire[93];							inform_L[87][3] = l_cell_wire[94];							inform_L[95][3] = l_cell_wire[95];							inform_L[96][3] = l_cell_wire[96];							inform_L[104][3] = l_cell_wire[97];							inform_L[97][3] = l_cell_wire[98];							inform_L[105][3] = l_cell_wire[99];							inform_L[98][3] = l_cell_wire[100];							inform_L[106][3] = l_cell_wire[101];							inform_L[99][3] = l_cell_wire[102];							inform_L[107][3] = l_cell_wire[103];							inform_L[100][3] = l_cell_wire[104];							inform_L[108][3] = l_cell_wire[105];							inform_L[101][3] = l_cell_wire[106];							inform_L[109][3] = l_cell_wire[107];							inform_L[102][3] = l_cell_wire[108];							inform_L[110][3] = l_cell_wire[109];							inform_L[103][3] = l_cell_wire[110];							inform_L[111][3] = l_cell_wire[111];							inform_L[112][3] = l_cell_wire[112];							inform_L[120][3] = l_cell_wire[113];							inform_L[113][3] = l_cell_wire[114];							inform_L[121][3] = l_cell_wire[115];							inform_L[114][3] = l_cell_wire[116];							inform_L[122][3] = l_cell_wire[117];							inform_L[115][3] = l_cell_wire[118];							inform_L[123][3] = l_cell_wire[119];							inform_L[116][3] = l_cell_wire[120];							inform_L[124][3] = l_cell_wire[121];							inform_L[117][3] = l_cell_wire[122];							inform_L[125][3] = l_cell_wire[123];							inform_L[118][3] = l_cell_wire[124];							inform_L[126][3] = l_cell_wire[125];							inform_L[119][3] = l_cell_wire[126];							inform_L[127][3] = l_cell_wire[127];						end
						5:						begin							inform_R[0][5] = r_cell_wire[0];							inform_R[16][5] = r_cell_wire[1];							inform_R[1][5] = r_cell_wire[2];							inform_R[17][5] = r_cell_wire[3];							inform_R[2][5] = r_cell_wire[4];							inform_R[18][5] = r_cell_wire[5];							inform_R[3][5] = r_cell_wire[6];							inform_R[19][5] = r_cell_wire[7];							inform_R[4][5] = r_cell_wire[8];							inform_R[20][5] = r_cell_wire[9];							inform_R[5][5] = r_cell_wire[10];							inform_R[21][5] = r_cell_wire[11];							inform_R[6][5] = r_cell_wire[12];							inform_R[22][5] = r_cell_wire[13];							inform_R[7][5] = r_cell_wire[14];							inform_R[23][5] = r_cell_wire[15];							inform_R[8][5] = r_cell_wire[16];							inform_R[24][5] = r_cell_wire[17];							inform_R[9][5] = r_cell_wire[18];							inform_R[25][5] = r_cell_wire[19];							inform_R[10][5] = r_cell_wire[20];							inform_R[26][5] = r_cell_wire[21];							inform_R[11][5] = r_cell_wire[22];							inform_R[27][5] = r_cell_wire[23];							inform_R[12][5] = r_cell_wire[24];							inform_R[28][5] = r_cell_wire[25];							inform_R[13][5] = r_cell_wire[26];							inform_R[29][5] = r_cell_wire[27];							inform_R[14][5] = r_cell_wire[28];							inform_R[30][5] = r_cell_wire[29];							inform_R[15][5] = r_cell_wire[30];							inform_R[31][5] = r_cell_wire[31];							inform_R[32][5] = r_cell_wire[32];							inform_R[48][5] = r_cell_wire[33];							inform_R[33][5] = r_cell_wire[34];							inform_R[49][5] = r_cell_wire[35];							inform_R[34][5] = r_cell_wire[36];							inform_R[50][5] = r_cell_wire[37];							inform_R[35][5] = r_cell_wire[38];							inform_R[51][5] = r_cell_wire[39];							inform_R[36][5] = r_cell_wire[40];							inform_R[52][5] = r_cell_wire[41];							inform_R[37][5] = r_cell_wire[42];							inform_R[53][5] = r_cell_wire[43];							inform_R[38][5] = r_cell_wire[44];							inform_R[54][5] = r_cell_wire[45];							inform_R[39][5] = r_cell_wire[46];							inform_R[55][5] = r_cell_wire[47];							inform_R[40][5] = r_cell_wire[48];							inform_R[56][5] = r_cell_wire[49];							inform_R[41][5] = r_cell_wire[50];							inform_R[57][5] = r_cell_wire[51];							inform_R[42][5] = r_cell_wire[52];							inform_R[58][5] = r_cell_wire[53];							inform_R[43][5] = r_cell_wire[54];							inform_R[59][5] = r_cell_wire[55];							inform_R[44][5] = r_cell_wire[56];							inform_R[60][5] = r_cell_wire[57];							inform_R[45][5] = r_cell_wire[58];							inform_R[61][5] = r_cell_wire[59];							inform_R[46][5] = r_cell_wire[60];							inform_R[62][5] = r_cell_wire[61];							inform_R[47][5] = r_cell_wire[62];							inform_R[63][5] = r_cell_wire[63];							inform_R[64][5] = r_cell_wire[64];							inform_R[80][5] = r_cell_wire[65];							inform_R[65][5] = r_cell_wire[66];							inform_R[81][5] = r_cell_wire[67];							inform_R[66][5] = r_cell_wire[68];							inform_R[82][5] = r_cell_wire[69];							inform_R[67][5] = r_cell_wire[70];							inform_R[83][5] = r_cell_wire[71];							inform_R[68][5] = r_cell_wire[72];							inform_R[84][5] = r_cell_wire[73];							inform_R[69][5] = r_cell_wire[74];							inform_R[85][5] = r_cell_wire[75];							inform_R[70][5] = r_cell_wire[76];							inform_R[86][5] = r_cell_wire[77];							inform_R[71][5] = r_cell_wire[78];							inform_R[87][5] = r_cell_wire[79];							inform_R[72][5] = r_cell_wire[80];							inform_R[88][5] = r_cell_wire[81];							inform_R[73][5] = r_cell_wire[82];							inform_R[89][5] = r_cell_wire[83];							inform_R[74][5] = r_cell_wire[84];							inform_R[90][5] = r_cell_wire[85];							inform_R[75][5] = r_cell_wire[86];							inform_R[91][5] = r_cell_wire[87];							inform_R[76][5] = r_cell_wire[88];							inform_R[92][5] = r_cell_wire[89];							inform_R[77][5] = r_cell_wire[90];							inform_R[93][5] = r_cell_wire[91];							inform_R[78][5] = r_cell_wire[92];							inform_R[94][5] = r_cell_wire[93];							inform_R[79][5] = r_cell_wire[94];							inform_R[95][5] = r_cell_wire[95];							inform_R[96][5] = r_cell_wire[96];							inform_R[112][5] = r_cell_wire[97];							inform_R[97][5] = r_cell_wire[98];							inform_R[113][5] = r_cell_wire[99];							inform_R[98][5] = r_cell_wire[100];							inform_R[114][5] = r_cell_wire[101];							inform_R[99][5] = r_cell_wire[102];							inform_R[115][5] = r_cell_wire[103];							inform_R[100][5] = r_cell_wire[104];							inform_R[116][5] = r_cell_wire[105];							inform_R[101][5] = r_cell_wire[106];							inform_R[117][5] = r_cell_wire[107];							inform_R[102][5] = r_cell_wire[108];							inform_R[118][5] = r_cell_wire[109];							inform_R[103][5] = r_cell_wire[110];							inform_R[119][5] = r_cell_wire[111];							inform_R[104][5] = r_cell_wire[112];							inform_R[120][5] = r_cell_wire[113];							inform_R[105][5] = r_cell_wire[114];							inform_R[121][5] = r_cell_wire[115];							inform_R[106][5] = r_cell_wire[116];							inform_R[122][5] = r_cell_wire[117];							inform_R[107][5] = r_cell_wire[118];							inform_R[123][5] = r_cell_wire[119];							inform_R[108][5] = r_cell_wire[120];							inform_R[124][5] = r_cell_wire[121];							inform_R[109][5] = r_cell_wire[122];							inform_R[125][5] = r_cell_wire[123];							inform_R[110][5] = r_cell_wire[124];							inform_R[126][5] = r_cell_wire[125];							inform_R[111][5] = r_cell_wire[126];							inform_R[127][5] = r_cell_wire[127];							inform_L[0][4] = l_cell_wire[0];							inform_L[16][4] = l_cell_wire[1];							inform_L[1][4] = l_cell_wire[2];							inform_L[17][4] = l_cell_wire[3];							inform_L[2][4] = l_cell_wire[4];							inform_L[18][4] = l_cell_wire[5];							inform_L[3][4] = l_cell_wire[6];							inform_L[19][4] = l_cell_wire[7];							inform_L[4][4] = l_cell_wire[8];							inform_L[20][4] = l_cell_wire[9];							inform_L[5][4] = l_cell_wire[10];							inform_L[21][4] = l_cell_wire[11];							inform_L[6][4] = l_cell_wire[12];							inform_L[22][4] = l_cell_wire[13];							inform_L[7][4] = l_cell_wire[14];							inform_L[23][4] = l_cell_wire[15];							inform_L[8][4] = l_cell_wire[16];							inform_L[24][4] = l_cell_wire[17];							inform_L[9][4] = l_cell_wire[18];							inform_L[25][4] = l_cell_wire[19];							inform_L[10][4] = l_cell_wire[20];							inform_L[26][4] = l_cell_wire[21];							inform_L[11][4] = l_cell_wire[22];							inform_L[27][4] = l_cell_wire[23];							inform_L[12][4] = l_cell_wire[24];							inform_L[28][4] = l_cell_wire[25];							inform_L[13][4] = l_cell_wire[26];							inform_L[29][4] = l_cell_wire[27];							inform_L[14][4] = l_cell_wire[28];							inform_L[30][4] = l_cell_wire[29];							inform_L[15][4] = l_cell_wire[30];							inform_L[31][4] = l_cell_wire[31];							inform_L[32][4] = l_cell_wire[32];							inform_L[48][4] = l_cell_wire[33];							inform_L[33][4] = l_cell_wire[34];							inform_L[49][4] = l_cell_wire[35];							inform_L[34][4] = l_cell_wire[36];							inform_L[50][4] = l_cell_wire[37];							inform_L[35][4] = l_cell_wire[38];							inform_L[51][4] = l_cell_wire[39];							inform_L[36][4] = l_cell_wire[40];							inform_L[52][4] = l_cell_wire[41];							inform_L[37][4] = l_cell_wire[42];							inform_L[53][4] = l_cell_wire[43];							inform_L[38][4] = l_cell_wire[44];							inform_L[54][4] = l_cell_wire[45];							inform_L[39][4] = l_cell_wire[46];							inform_L[55][4] = l_cell_wire[47];							inform_L[40][4] = l_cell_wire[48];							inform_L[56][4] = l_cell_wire[49];							inform_L[41][4] = l_cell_wire[50];							inform_L[57][4] = l_cell_wire[51];							inform_L[42][4] = l_cell_wire[52];							inform_L[58][4] = l_cell_wire[53];							inform_L[43][4] = l_cell_wire[54];							inform_L[59][4] = l_cell_wire[55];							inform_L[44][4] = l_cell_wire[56];							inform_L[60][4] = l_cell_wire[57];							inform_L[45][4] = l_cell_wire[58];							inform_L[61][4] = l_cell_wire[59];							inform_L[46][4] = l_cell_wire[60];							inform_L[62][4] = l_cell_wire[61];							inform_L[47][4] = l_cell_wire[62];							inform_L[63][4] = l_cell_wire[63];							inform_L[64][4] = l_cell_wire[64];							inform_L[80][4] = l_cell_wire[65];							inform_L[65][4] = l_cell_wire[66];							inform_L[81][4] = l_cell_wire[67];							inform_L[66][4] = l_cell_wire[68];							inform_L[82][4] = l_cell_wire[69];							inform_L[67][4] = l_cell_wire[70];							inform_L[83][4] = l_cell_wire[71];							inform_L[68][4] = l_cell_wire[72];							inform_L[84][4] = l_cell_wire[73];							inform_L[69][4] = l_cell_wire[74];							inform_L[85][4] = l_cell_wire[75];							inform_L[70][4] = l_cell_wire[76];							inform_L[86][4] = l_cell_wire[77];							inform_L[71][4] = l_cell_wire[78];							inform_L[87][4] = l_cell_wire[79];							inform_L[72][4] = l_cell_wire[80];							inform_L[88][4] = l_cell_wire[81];							inform_L[73][4] = l_cell_wire[82];							inform_L[89][4] = l_cell_wire[83];							inform_L[74][4] = l_cell_wire[84];							inform_L[90][4] = l_cell_wire[85];							inform_L[75][4] = l_cell_wire[86];							inform_L[91][4] = l_cell_wire[87];							inform_L[76][4] = l_cell_wire[88];							inform_L[92][4] = l_cell_wire[89];							inform_L[77][4] = l_cell_wire[90];							inform_L[93][4] = l_cell_wire[91];							inform_L[78][4] = l_cell_wire[92];							inform_L[94][4] = l_cell_wire[93];							inform_L[79][4] = l_cell_wire[94];							inform_L[95][4] = l_cell_wire[95];							inform_L[96][4] = l_cell_wire[96];							inform_L[112][4] = l_cell_wire[97];							inform_L[97][4] = l_cell_wire[98];							inform_L[113][4] = l_cell_wire[99];							inform_L[98][4] = l_cell_wire[100];							inform_L[114][4] = l_cell_wire[101];							inform_L[99][4] = l_cell_wire[102];							inform_L[115][4] = l_cell_wire[103];							inform_L[100][4] = l_cell_wire[104];							inform_L[116][4] = l_cell_wire[105];							inform_L[101][4] = l_cell_wire[106];							inform_L[117][4] = l_cell_wire[107];							inform_L[102][4] = l_cell_wire[108];							inform_L[118][4] = l_cell_wire[109];							inform_L[103][4] = l_cell_wire[110];							inform_L[119][4] = l_cell_wire[111];							inform_L[104][4] = l_cell_wire[112];							inform_L[120][4] = l_cell_wire[113];							inform_L[105][4] = l_cell_wire[114];							inform_L[121][4] = l_cell_wire[115];							inform_L[106][4] = l_cell_wire[116];							inform_L[122][4] = l_cell_wire[117];							inform_L[107][4] = l_cell_wire[118];							inform_L[123][4] = l_cell_wire[119];							inform_L[108][4] = l_cell_wire[120];							inform_L[124][4] = l_cell_wire[121];							inform_L[109][4] = l_cell_wire[122];							inform_L[125][4] = l_cell_wire[123];							inform_L[110][4] = l_cell_wire[124];							inform_L[126][4] = l_cell_wire[125];							inform_L[111][4] = l_cell_wire[126];							inform_L[127][4] = l_cell_wire[127];						end
						6:						begin							inform_R[0][6] = r_cell_wire[0];							inform_R[32][6] = r_cell_wire[1];							inform_R[1][6] = r_cell_wire[2];							inform_R[33][6] = r_cell_wire[3];							inform_R[2][6] = r_cell_wire[4];							inform_R[34][6] = r_cell_wire[5];							inform_R[3][6] = r_cell_wire[6];							inform_R[35][6] = r_cell_wire[7];							inform_R[4][6] = r_cell_wire[8];							inform_R[36][6] = r_cell_wire[9];							inform_R[5][6] = r_cell_wire[10];							inform_R[37][6] = r_cell_wire[11];							inform_R[6][6] = r_cell_wire[12];							inform_R[38][6] = r_cell_wire[13];							inform_R[7][6] = r_cell_wire[14];							inform_R[39][6] = r_cell_wire[15];							inform_R[8][6] = r_cell_wire[16];							inform_R[40][6] = r_cell_wire[17];							inform_R[9][6] = r_cell_wire[18];							inform_R[41][6] = r_cell_wire[19];							inform_R[10][6] = r_cell_wire[20];							inform_R[42][6] = r_cell_wire[21];							inform_R[11][6] = r_cell_wire[22];							inform_R[43][6] = r_cell_wire[23];							inform_R[12][6] = r_cell_wire[24];							inform_R[44][6] = r_cell_wire[25];							inform_R[13][6] = r_cell_wire[26];							inform_R[45][6] = r_cell_wire[27];							inform_R[14][6] = r_cell_wire[28];							inform_R[46][6] = r_cell_wire[29];							inform_R[15][6] = r_cell_wire[30];							inform_R[47][6] = r_cell_wire[31];							inform_R[16][6] = r_cell_wire[32];							inform_R[48][6] = r_cell_wire[33];							inform_R[17][6] = r_cell_wire[34];							inform_R[49][6] = r_cell_wire[35];							inform_R[18][6] = r_cell_wire[36];							inform_R[50][6] = r_cell_wire[37];							inform_R[19][6] = r_cell_wire[38];							inform_R[51][6] = r_cell_wire[39];							inform_R[20][6] = r_cell_wire[40];							inform_R[52][6] = r_cell_wire[41];							inform_R[21][6] = r_cell_wire[42];							inform_R[53][6] = r_cell_wire[43];							inform_R[22][6] = r_cell_wire[44];							inform_R[54][6] = r_cell_wire[45];							inform_R[23][6] = r_cell_wire[46];							inform_R[55][6] = r_cell_wire[47];							inform_R[24][6] = r_cell_wire[48];							inform_R[56][6] = r_cell_wire[49];							inform_R[25][6] = r_cell_wire[50];							inform_R[57][6] = r_cell_wire[51];							inform_R[26][6] = r_cell_wire[52];							inform_R[58][6] = r_cell_wire[53];							inform_R[27][6] = r_cell_wire[54];							inform_R[59][6] = r_cell_wire[55];							inform_R[28][6] = r_cell_wire[56];							inform_R[60][6] = r_cell_wire[57];							inform_R[29][6] = r_cell_wire[58];							inform_R[61][6] = r_cell_wire[59];							inform_R[30][6] = r_cell_wire[60];							inform_R[62][6] = r_cell_wire[61];							inform_R[31][6] = r_cell_wire[62];							inform_R[63][6] = r_cell_wire[63];							inform_R[64][6] = r_cell_wire[64];							inform_R[96][6] = r_cell_wire[65];							inform_R[65][6] = r_cell_wire[66];							inform_R[97][6] = r_cell_wire[67];							inform_R[66][6] = r_cell_wire[68];							inform_R[98][6] = r_cell_wire[69];							inform_R[67][6] = r_cell_wire[70];							inform_R[99][6] = r_cell_wire[71];							inform_R[68][6] = r_cell_wire[72];							inform_R[100][6] = r_cell_wire[73];							inform_R[69][6] = r_cell_wire[74];							inform_R[101][6] = r_cell_wire[75];							inform_R[70][6] = r_cell_wire[76];							inform_R[102][6] = r_cell_wire[77];							inform_R[71][6] = r_cell_wire[78];							inform_R[103][6] = r_cell_wire[79];							inform_R[72][6] = r_cell_wire[80];							inform_R[104][6] = r_cell_wire[81];							inform_R[73][6] = r_cell_wire[82];							inform_R[105][6] = r_cell_wire[83];							inform_R[74][6] = r_cell_wire[84];							inform_R[106][6] = r_cell_wire[85];							inform_R[75][6] = r_cell_wire[86];							inform_R[107][6] = r_cell_wire[87];							inform_R[76][6] = r_cell_wire[88];							inform_R[108][6] = r_cell_wire[89];							inform_R[77][6] = r_cell_wire[90];							inform_R[109][6] = r_cell_wire[91];							inform_R[78][6] = r_cell_wire[92];							inform_R[110][6] = r_cell_wire[93];							inform_R[79][6] = r_cell_wire[94];							inform_R[111][6] = r_cell_wire[95];							inform_R[80][6] = r_cell_wire[96];							inform_R[112][6] = r_cell_wire[97];							inform_R[81][6] = r_cell_wire[98];							inform_R[113][6] = r_cell_wire[99];							inform_R[82][6] = r_cell_wire[100];							inform_R[114][6] = r_cell_wire[101];							inform_R[83][6] = r_cell_wire[102];							inform_R[115][6] = r_cell_wire[103];							inform_R[84][6] = r_cell_wire[104];							inform_R[116][6] = r_cell_wire[105];							inform_R[85][6] = r_cell_wire[106];							inform_R[117][6] = r_cell_wire[107];							inform_R[86][6] = r_cell_wire[108];							inform_R[118][6] = r_cell_wire[109];							inform_R[87][6] = r_cell_wire[110];							inform_R[119][6] = r_cell_wire[111];							inform_R[88][6] = r_cell_wire[112];							inform_R[120][6] = r_cell_wire[113];							inform_R[89][6] = r_cell_wire[114];							inform_R[121][6] = r_cell_wire[115];							inform_R[90][6] = r_cell_wire[116];							inform_R[122][6] = r_cell_wire[117];							inform_R[91][6] = r_cell_wire[118];							inform_R[123][6] = r_cell_wire[119];							inform_R[92][6] = r_cell_wire[120];							inform_R[124][6] = r_cell_wire[121];							inform_R[93][6] = r_cell_wire[122];							inform_R[125][6] = r_cell_wire[123];							inform_R[94][6] = r_cell_wire[124];							inform_R[126][6] = r_cell_wire[125];							inform_R[95][6] = r_cell_wire[126];							inform_R[127][6] = r_cell_wire[127];							inform_L[0][5] = l_cell_wire[0];							inform_L[32][5] = l_cell_wire[1];							inform_L[1][5] = l_cell_wire[2];							inform_L[33][5] = l_cell_wire[3];							inform_L[2][5] = l_cell_wire[4];							inform_L[34][5] = l_cell_wire[5];							inform_L[3][5] = l_cell_wire[6];							inform_L[35][5] = l_cell_wire[7];							inform_L[4][5] = l_cell_wire[8];							inform_L[36][5] = l_cell_wire[9];							inform_L[5][5] = l_cell_wire[10];							inform_L[37][5] = l_cell_wire[11];							inform_L[6][5] = l_cell_wire[12];							inform_L[38][5] = l_cell_wire[13];							inform_L[7][5] = l_cell_wire[14];							inform_L[39][5] = l_cell_wire[15];							inform_L[8][5] = l_cell_wire[16];							inform_L[40][5] = l_cell_wire[17];							inform_L[9][5] = l_cell_wire[18];							inform_L[41][5] = l_cell_wire[19];							inform_L[10][5] = l_cell_wire[20];							inform_L[42][5] = l_cell_wire[21];							inform_L[11][5] = l_cell_wire[22];							inform_L[43][5] = l_cell_wire[23];							inform_L[12][5] = l_cell_wire[24];							inform_L[44][5] = l_cell_wire[25];							inform_L[13][5] = l_cell_wire[26];							inform_L[45][5] = l_cell_wire[27];							inform_L[14][5] = l_cell_wire[28];							inform_L[46][5] = l_cell_wire[29];							inform_L[15][5] = l_cell_wire[30];							inform_L[47][5] = l_cell_wire[31];							inform_L[16][5] = l_cell_wire[32];							inform_L[48][5] = l_cell_wire[33];							inform_L[17][5] = l_cell_wire[34];							inform_L[49][5] = l_cell_wire[35];							inform_L[18][5] = l_cell_wire[36];							inform_L[50][5] = l_cell_wire[37];							inform_L[19][5] = l_cell_wire[38];							inform_L[51][5] = l_cell_wire[39];							inform_L[20][5] = l_cell_wire[40];							inform_L[52][5] = l_cell_wire[41];							inform_L[21][5] = l_cell_wire[42];							inform_L[53][5] = l_cell_wire[43];							inform_L[22][5] = l_cell_wire[44];							inform_L[54][5] = l_cell_wire[45];							inform_L[23][5] = l_cell_wire[46];							inform_L[55][5] = l_cell_wire[47];							inform_L[24][5] = l_cell_wire[48];							inform_L[56][5] = l_cell_wire[49];							inform_L[25][5] = l_cell_wire[50];							inform_L[57][5] = l_cell_wire[51];							inform_L[26][5] = l_cell_wire[52];							inform_L[58][5] = l_cell_wire[53];							inform_L[27][5] = l_cell_wire[54];							inform_L[59][5] = l_cell_wire[55];							inform_L[28][5] = l_cell_wire[56];							inform_L[60][5] = l_cell_wire[57];							inform_L[29][5] = l_cell_wire[58];							inform_L[61][5] = l_cell_wire[59];							inform_L[30][5] = l_cell_wire[60];							inform_L[62][5] = l_cell_wire[61];							inform_L[31][5] = l_cell_wire[62];							inform_L[63][5] = l_cell_wire[63];							inform_L[64][5] = l_cell_wire[64];							inform_L[96][5] = l_cell_wire[65];							inform_L[65][5] = l_cell_wire[66];							inform_L[97][5] = l_cell_wire[67];							inform_L[66][5] = l_cell_wire[68];							inform_L[98][5] = l_cell_wire[69];							inform_L[67][5] = l_cell_wire[70];							inform_L[99][5] = l_cell_wire[71];							inform_L[68][5] = l_cell_wire[72];							inform_L[100][5] = l_cell_wire[73];							inform_L[69][5] = l_cell_wire[74];							inform_L[101][5] = l_cell_wire[75];							inform_L[70][5] = l_cell_wire[76];							inform_L[102][5] = l_cell_wire[77];							inform_L[71][5] = l_cell_wire[78];							inform_L[103][5] = l_cell_wire[79];							inform_L[72][5] = l_cell_wire[80];							inform_L[104][5] = l_cell_wire[81];							inform_L[73][5] = l_cell_wire[82];							inform_L[105][5] = l_cell_wire[83];							inform_L[74][5] = l_cell_wire[84];							inform_L[106][5] = l_cell_wire[85];							inform_L[75][5] = l_cell_wire[86];							inform_L[107][5] = l_cell_wire[87];							inform_L[76][5] = l_cell_wire[88];							inform_L[108][5] = l_cell_wire[89];							inform_L[77][5] = l_cell_wire[90];							inform_L[109][5] = l_cell_wire[91];							inform_L[78][5] = l_cell_wire[92];							inform_L[110][5] = l_cell_wire[93];							inform_L[79][5] = l_cell_wire[94];							inform_L[111][5] = l_cell_wire[95];							inform_L[80][5] = l_cell_wire[96];							inform_L[112][5] = l_cell_wire[97];							inform_L[81][5] = l_cell_wire[98];							inform_L[113][5] = l_cell_wire[99];							inform_L[82][5] = l_cell_wire[100];							inform_L[114][5] = l_cell_wire[101];							inform_L[83][5] = l_cell_wire[102];							inform_L[115][5] = l_cell_wire[103];							inform_L[84][5] = l_cell_wire[104];							inform_L[116][5] = l_cell_wire[105];							inform_L[85][5] = l_cell_wire[106];							inform_L[117][5] = l_cell_wire[107];							inform_L[86][5] = l_cell_wire[108];							inform_L[118][5] = l_cell_wire[109];							inform_L[87][5] = l_cell_wire[110];							inform_L[119][5] = l_cell_wire[111];							inform_L[88][5] = l_cell_wire[112];							inform_L[120][5] = l_cell_wire[113];							inform_L[89][5] = l_cell_wire[114];							inform_L[121][5] = l_cell_wire[115];							inform_L[90][5] = l_cell_wire[116];							inform_L[122][5] = l_cell_wire[117];							inform_L[91][5] = l_cell_wire[118];							inform_L[123][5] = l_cell_wire[119];							inform_L[92][5] = l_cell_wire[120];							inform_L[124][5] = l_cell_wire[121];							inform_L[93][5] = l_cell_wire[122];							inform_L[125][5] = l_cell_wire[123];							inform_L[94][5] = l_cell_wire[124];							inform_L[126][5] = l_cell_wire[125];							inform_L[95][5] = l_cell_wire[126];							inform_L[127][5] = l_cell_wire[127];						end
						7:						begin							inform_R[0][7] = r_cell_wire[0];							inform_R[64][7] = r_cell_wire[1];							inform_R[1][7] = r_cell_wire[2];							inform_R[65][7] = r_cell_wire[3];							inform_R[2][7] = r_cell_wire[4];							inform_R[66][7] = r_cell_wire[5];							inform_R[3][7] = r_cell_wire[6];							inform_R[67][7] = r_cell_wire[7];							inform_R[4][7] = r_cell_wire[8];							inform_R[68][7] = r_cell_wire[9];							inform_R[5][7] = r_cell_wire[10];							inform_R[69][7] = r_cell_wire[11];							inform_R[6][7] = r_cell_wire[12];							inform_R[70][7] = r_cell_wire[13];							inform_R[7][7] = r_cell_wire[14];							inform_R[71][7] = r_cell_wire[15];							inform_R[8][7] = r_cell_wire[16];							inform_R[72][7] = r_cell_wire[17];							inform_R[9][7] = r_cell_wire[18];							inform_R[73][7] = r_cell_wire[19];							inform_R[10][7] = r_cell_wire[20];							inform_R[74][7] = r_cell_wire[21];							inform_R[11][7] = r_cell_wire[22];							inform_R[75][7] = r_cell_wire[23];							inform_R[12][7] = r_cell_wire[24];							inform_R[76][7] = r_cell_wire[25];							inform_R[13][7] = r_cell_wire[26];							inform_R[77][7] = r_cell_wire[27];							inform_R[14][7] = r_cell_wire[28];							inform_R[78][7] = r_cell_wire[29];							inform_R[15][7] = r_cell_wire[30];							inform_R[79][7] = r_cell_wire[31];							inform_R[16][7] = r_cell_wire[32];							inform_R[80][7] = r_cell_wire[33];							inform_R[17][7] = r_cell_wire[34];							inform_R[81][7] = r_cell_wire[35];							inform_R[18][7] = r_cell_wire[36];							inform_R[82][7] = r_cell_wire[37];							inform_R[19][7] = r_cell_wire[38];							inform_R[83][7] = r_cell_wire[39];							inform_R[20][7] = r_cell_wire[40];							inform_R[84][7] = r_cell_wire[41];							inform_R[21][7] = r_cell_wire[42];							inform_R[85][7] = r_cell_wire[43];							inform_R[22][7] = r_cell_wire[44];							inform_R[86][7] = r_cell_wire[45];							inform_R[23][7] = r_cell_wire[46];							inform_R[87][7] = r_cell_wire[47];							inform_R[24][7] = r_cell_wire[48];							inform_R[88][7] = r_cell_wire[49];							inform_R[25][7] = r_cell_wire[50];							inform_R[89][7] = r_cell_wire[51];							inform_R[26][7] = r_cell_wire[52];							inform_R[90][7] = r_cell_wire[53];							inform_R[27][7] = r_cell_wire[54];							inform_R[91][7] = r_cell_wire[55];							inform_R[28][7] = r_cell_wire[56];							inform_R[92][7] = r_cell_wire[57];							inform_R[29][7] = r_cell_wire[58];							inform_R[93][7] = r_cell_wire[59];							inform_R[30][7] = r_cell_wire[60];							inform_R[94][7] = r_cell_wire[61];							inform_R[31][7] = r_cell_wire[62];							inform_R[95][7] = r_cell_wire[63];							inform_R[32][7] = r_cell_wire[64];							inform_R[96][7] = r_cell_wire[65];							inform_R[33][7] = r_cell_wire[66];							inform_R[97][7] = r_cell_wire[67];							inform_R[34][7] = r_cell_wire[68];							inform_R[98][7] = r_cell_wire[69];							inform_R[35][7] = r_cell_wire[70];							inform_R[99][7] = r_cell_wire[71];							inform_R[36][7] = r_cell_wire[72];							inform_R[100][7] = r_cell_wire[73];							inform_R[37][7] = r_cell_wire[74];							inform_R[101][7] = r_cell_wire[75];							inform_R[38][7] = r_cell_wire[76];							inform_R[102][7] = r_cell_wire[77];							inform_R[39][7] = r_cell_wire[78];							inform_R[103][7] = r_cell_wire[79];							inform_R[40][7] = r_cell_wire[80];							inform_R[104][7] = r_cell_wire[81];							inform_R[41][7] = r_cell_wire[82];							inform_R[105][7] = r_cell_wire[83];							inform_R[42][7] = r_cell_wire[84];							inform_R[106][7] = r_cell_wire[85];							inform_R[43][7] = r_cell_wire[86];							inform_R[107][7] = r_cell_wire[87];							inform_R[44][7] = r_cell_wire[88];							inform_R[108][7] = r_cell_wire[89];							inform_R[45][7] = r_cell_wire[90];							inform_R[109][7] = r_cell_wire[91];							inform_R[46][7] = r_cell_wire[92];							inform_R[110][7] = r_cell_wire[93];							inform_R[47][7] = r_cell_wire[94];							inform_R[111][7] = r_cell_wire[95];							inform_R[48][7] = r_cell_wire[96];							inform_R[112][7] = r_cell_wire[97];							inform_R[49][7] = r_cell_wire[98];							inform_R[113][7] = r_cell_wire[99];							inform_R[50][7] = r_cell_wire[100];							inform_R[114][7] = r_cell_wire[101];							inform_R[51][7] = r_cell_wire[102];							inform_R[115][7] = r_cell_wire[103];							inform_R[52][7] = r_cell_wire[104];							inform_R[116][7] = r_cell_wire[105];							inform_R[53][7] = r_cell_wire[106];							inform_R[117][7] = r_cell_wire[107];							inform_R[54][7] = r_cell_wire[108];							inform_R[118][7] = r_cell_wire[109];							inform_R[55][7] = r_cell_wire[110];							inform_R[119][7] = r_cell_wire[111];							inform_R[56][7] = r_cell_wire[112];							inform_R[120][7] = r_cell_wire[113];							inform_R[57][7] = r_cell_wire[114];							inform_R[121][7] = r_cell_wire[115];							inform_R[58][7] = r_cell_wire[116];							inform_R[122][7] = r_cell_wire[117];							inform_R[59][7] = r_cell_wire[118];							inform_R[123][7] = r_cell_wire[119];							inform_R[60][7] = r_cell_wire[120];							inform_R[124][7] = r_cell_wire[121];							inform_R[61][7] = r_cell_wire[122];							inform_R[125][7] = r_cell_wire[123];							inform_R[62][7] = r_cell_wire[124];							inform_R[126][7] = r_cell_wire[125];							inform_R[63][7] = r_cell_wire[126];							inform_R[127][7] = r_cell_wire[127];							inform_L[0][6] = l_cell_wire[0];							inform_L[64][6] = l_cell_wire[1];							inform_L[1][6] = l_cell_wire[2];							inform_L[65][6] = l_cell_wire[3];							inform_L[2][6] = l_cell_wire[4];							inform_L[66][6] = l_cell_wire[5];							inform_L[3][6] = l_cell_wire[6];							inform_L[67][6] = l_cell_wire[7];							inform_L[4][6] = l_cell_wire[8];							inform_L[68][6] = l_cell_wire[9];							inform_L[5][6] = l_cell_wire[10];							inform_L[69][6] = l_cell_wire[11];							inform_L[6][6] = l_cell_wire[12];							inform_L[70][6] = l_cell_wire[13];							inform_L[7][6] = l_cell_wire[14];							inform_L[71][6] = l_cell_wire[15];							inform_L[8][6] = l_cell_wire[16];							inform_L[72][6] = l_cell_wire[17];							inform_L[9][6] = l_cell_wire[18];							inform_L[73][6] = l_cell_wire[19];							inform_L[10][6] = l_cell_wire[20];							inform_L[74][6] = l_cell_wire[21];							inform_L[11][6] = l_cell_wire[22];							inform_L[75][6] = l_cell_wire[23];							inform_L[12][6] = l_cell_wire[24];							inform_L[76][6] = l_cell_wire[25];							inform_L[13][6] = l_cell_wire[26];							inform_L[77][6] = l_cell_wire[27];							inform_L[14][6] = l_cell_wire[28];							inform_L[78][6] = l_cell_wire[29];							inform_L[15][6] = l_cell_wire[30];							inform_L[79][6] = l_cell_wire[31];							inform_L[16][6] = l_cell_wire[32];							inform_L[80][6] = l_cell_wire[33];							inform_L[17][6] = l_cell_wire[34];							inform_L[81][6] = l_cell_wire[35];							inform_L[18][6] = l_cell_wire[36];							inform_L[82][6] = l_cell_wire[37];							inform_L[19][6] = l_cell_wire[38];							inform_L[83][6] = l_cell_wire[39];							inform_L[20][6] = l_cell_wire[40];							inform_L[84][6] = l_cell_wire[41];							inform_L[21][6] = l_cell_wire[42];							inform_L[85][6] = l_cell_wire[43];							inform_L[22][6] = l_cell_wire[44];							inform_L[86][6] = l_cell_wire[45];							inform_L[23][6] = l_cell_wire[46];							inform_L[87][6] = l_cell_wire[47];							inform_L[24][6] = l_cell_wire[48];							inform_L[88][6] = l_cell_wire[49];							inform_L[25][6] = l_cell_wire[50];							inform_L[89][6] = l_cell_wire[51];							inform_L[26][6] = l_cell_wire[52];							inform_L[90][6] = l_cell_wire[53];							inform_L[27][6] = l_cell_wire[54];							inform_L[91][6] = l_cell_wire[55];							inform_L[28][6] = l_cell_wire[56];							inform_L[92][6] = l_cell_wire[57];							inform_L[29][6] = l_cell_wire[58];							inform_L[93][6] = l_cell_wire[59];							inform_L[30][6] = l_cell_wire[60];							inform_L[94][6] = l_cell_wire[61];							inform_L[31][6] = l_cell_wire[62];							inform_L[95][6] = l_cell_wire[63];							inform_L[32][6] = l_cell_wire[64];							inform_L[96][6] = l_cell_wire[65];							inform_L[33][6] = l_cell_wire[66];							inform_L[97][6] = l_cell_wire[67];							inform_L[34][6] = l_cell_wire[68];							inform_L[98][6] = l_cell_wire[69];							inform_L[35][6] = l_cell_wire[70];							inform_L[99][6] = l_cell_wire[71];							inform_L[36][6] = l_cell_wire[72];							inform_L[100][6] = l_cell_wire[73];							inform_L[37][6] = l_cell_wire[74];							inform_L[101][6] = l_cell_wire[75];							inform_L[38][6] = l_cell_wire[76];							inform_L[102][6] = l_cell_wire[77];							inform_L[39][6] = l_cell_wire[78];							inform_L[103][6] = l_cell_wire[79];							inform_L[40][6] = l_cell_wire[80];							inform_L[104][6] = l_cell_wire[81];							inform_L[41][6] = l_cell_wire[82];							inform_L[105][6] = l_cell_wire[83];							inform_L[42][6] = l_cell_wire[84];							inform_L[106][6] = l_cell_wire[85];							inform_L[43][6] = l_cell_wire[86];							inform_L[107][6] = l_cell_wire[87];							inform_L[44][6] = l_cell_wire[88];							inform_L[108][6] = l_cell_wire[89];							inform_L[45][6] = l_cell_wire[90];							inform_L[109][6] = l_cell_wire[91];							inform_L[46][6] = l_cell_wire[92];							inform_L[110][6] = l_cell_wire[93];							inform_L[47][6] = l_cell_wire[94];							inform_L[111][6] = l_cell_wire[95];							inform_L[48][6] = l_cell_wire[96];							inform_L[112][6] = l_cell_wire[97];							inform_L[49][6] = l_cell_wire[98];							inform_L[113][6] = l_cell_wire[99];							inform_L[50][6] = l_cell_wire[100];							inform_L[114][6] = l_cell_wire[101];							inform_L[51][6] = l_cell_wire[102];							inform_L[115][6] = l_cell_wire[103];							inform_L[52][6] = l_cell_wire[104];							inform_L[116][6] = l_cell_wire[105];							inform_L[53][6] = l_cell_wire[106];							inform_L[117][6] = l_cell_wire[107];							inform_L[54][6] = l_cell_wire[108];							inform_L[118][6] = l_cell_wire[109];							inform_L[55][6] = l_cell_wire[110];							inform_L[119][6] = l_cell_wire[111];							inform_L[56][6] = l_cell_wire[112];							inform_L[120][6] = l_cell_wire[113];							inform_L[57][6] = l_cell_wire[114];							inform_L[121][6] = l_cell_wire[115];							inform_L[58][6] = l_cell_wire[116];							inform_L[122][6] = l_cell_wire[117];							inform_L[59][6] = l_cell_wire[118];							inform_L[123][6] = l_cell_wire[119];							inform_L[60][6] = l_cell_wire[120];							inform_L[124][6] = l_cell_wire[121];							inform_L[61][6] = l_cell_wire[122];							inform_L[125][6] = l_cell_wire[123];							inform_L[62][6] = l_cell_wire[124];							inform_L[126][6] = l_cell_wire[125];							inform_L[63][6] = l_cell_wire[126];							inform_L[127][6] = l_cell_wire[127];						end
						default:							for (x = 0; x < 128; x = x + 1)								for (y = 0; y < 7; y = y + 1)								begin									inform_R[x][y+1] <= 8'd0;									inform_L[x][y] <= 8'd0;								end					endcase				end			end
			BUSY_RIGHT:			begin				if(clk_counter == 2'b11)begin					case (w2r)						1:						begin							inform_R[0][1] = r_cell_wire[0];							inform_R[1][1] = r_cell_wire[1];							inform_R[2][1] = r_cell_wire[2];							inform_R[3][1] = r_cell_wire[3];							inform_R[4][1] = r_cell_wire[4];							inform_R[5][1] = r_cell_wire[5];							inform_R[6][1] = r_cell_wire[6];							inform_R[7][1] = r_cell_wire[7];							inform_R[8][1] = r_cell_wire[8];							inform_R[9][1] = r_cell_wire[9];							inform_R[10][1] = r_cell_wire[10];							inform_R[11][1] = r_cell_wire[11];							inform_R[12][1] = r_cell_wire[12];							inform_R[13][1] = r_cell_wire[13];							inform_R[14][1] = r_cell_wire[14];							inform_R[15][1] = r_cell_wire[15];							inform_R[16][1] = r_cell_wire[16];							inform_R[17][1] = r_cell_wire[17];							inform_R[18][1] = r_cell_wire[18];							inform_R[19][1] = r_cell_wire[19];							inform_R[20][1] = r_cell_wire[20];							inform_R[21][1] = r_cell_wire[21];							inform_R[22][1] = r_cell_wire[22];							inform_R[23][1] = r_cell_wire[23];							inform_R[24][1] = r_cell_wire[24];							inform_R[25][1] = r_cell_wire[25];							inform_R[26][1] = r_cell_wire[26];							inform_R[27][1] = r_cell_wire[27];							inform_R[28][1] = r_cell_wire[28];							inform_R[29][1] = r_cell_wire[29];							inform_R[30][1] = r_cell_wire[30];							inform_R[31][1] = r_cell_wire[31];							inform_R[32][1] = r_cell_wire[32];							inform_R[33][1] = r_cell_wire[33];							inform_R[34][1] = r_cell_wire[34];							inform_R[35][1] = r_cell_wire[35];							inform_R[36][1] = r_cell_wire[36];							inform_R[37][1] = r_cell_wire[37];							inform_R[38][1] = r_cell_wire[38];							inform_R[39][1] = r_cell_wire[39];							inform_R[40][1] = r_cell_wire[40];							inform_R[41][1] = r_cell_wire[41];							inform_R[42][1] = r_cell_wire[42];							inform_R[43][1] = r_cell_wire[43];							inform_R[44][1] = r_cell_wire[44];							inform_R[45][1] = r_cell_wire[45];							inform_R[46][1] = r_cell_wire[46];							inform_R[47][1] = r_cell_wire[47];							inform_R[48][1] = r_cell_wire[48];							inform_R[49][1] = r_cell_wire[49];							inform_R[50][1] = r_cell_wire[50];							inform_R[51][1] = r_cell_wire[51];							inform_R[52][1] = r_cell_wire[52];							inform_R[53][1] = r_cell_wire[53];							inform_R[54][1] = r_cell_wire[54];							inform_R[55][1] = r_cell_wire[55];							inform_R[56][1] = r_cell_wire[56];							inform_R[57][1] = r_cell_wire[57];							inform_R[58][1] = r_cell_wire[58];							inform_R[59][1] = r_cell_wire[59];							inform_R[60][1] = r_cell_wire[60];							inform_R[61][1] = r_cell_wire[61];							inform_R[62][1] = r_cell_wire[62];							inform_R[63][1] = r_cell_wire[63];							inform_R[64][1] = r_cell_wire[64];							inform_R[65][1] = r_cell_wire[65];							inform_R[66][1] = r_cell_wire[66];							inform_R[67][1] = r_cell_wire[67];							inform_R[68][1] = r_cell_wire[68];							inform_R[69][1] = r_cell_wire[69];							inform_R[70][1] = r_cell_wire[70];							inform_R[71][1] = r_cell_wire[71];							inform_R[72][1] = r_cell_wire[72];							inform_R[73][1] = r_cell_wire[73];							inform_R[74][1] = r_cell_wire[74];							inform_R[75][1] = r_cell_wire[75];							inform_R[76][1] = r_cell_wire[76];							inform_R[77][1] = r_cell_wire[77];							inform_R[78][1] = r_cell_wire[78];							inform_R[79][1] = r_cell_wire[79];							inform_R[80][1] = r_cell_wire[80];							inform_R[81][1] = r_cell_wire[81];							inform_R[82][1] = r_cell_wire[82];							inform_R[83][1] = r_cell_wire[83];							inform_R[84][1] = r_cell_wire[84];							inform_R[85][1] = r_cell_wire[85];							inform_R[86][1] = r_cell_wire[86];							inform_R[87][1] = r_cell_wire[87];							inform_R[88][1] = r_cell_wire[88];							inform_R[89][1] = r_cell_wire[89];							inform_R[90][1] = r_cell_wire[90];							inform_R[91][1] = r_cell_wire[91];							inform_R[92][1] = r_cell_wire[92];							inform_R[93][1] = r_cell_wire[93];							inform_R[94][1] = r_cell_wire[94];							inform_R[95][1] = r_cell_wire[95];							inform_R[96][1] = r_cell_wire[96];							inform_R[97][1] = r_cell_wire[97];							inform_R[98][1] = r_cell_wire[98];							inform_R[99][1] = r_cell_wire[99];							inform_R[100][1] = r_cell_wire[100];							inform_R[101][1] = r_cell_wire[101];							inform_R[102][1] = r_cell_wire[102];							inform_R[103][1] = r_cell_wire[103];							inform_R[104][1] = r_cell_wire[104];							inform_R[105][1] = r_cell_wire[105];							inform_R[106][1] = r_cell_wire[106];							inform_R[107][1] = r_cell_wire[107];							inform_R[108][1] = r_cell_wire[108];							inform_R[109][1] = r_cell_wire[109];							inform_R[110][1] = r_cell_wire[110];							inform_R[111][1] = r_cell_wire[111];							inform_R[112][1] = r_cell_wire[112];							inform_R[113][1] = r_cell_wire[113];							inform_R[114][1] = r_cell_wire[114];							inform_R[115][1] = r_cell_wire[115];							inform_R[116][1] = r_cell_wire[116];							inform_R[117][1] = r_cell_wire[117];							inform_R[118][1] = r_cell_wire[118];							inform_R[119][1] = r_cell_wire[119];							inform_R[120][1] = r_cell_wire[120];							inform_R[121][1] = r_cell_wire[121];							inform_R[122][1] = r_cell_wire[122];							inform_R[123][1] = r_cell_wire[123];							inform_R[124][1] = r_cell_wire[124];							inform_R[125][1] = r_cell_wire[125];							inform_R[126][1] = r_cell_wire[126];							inform_R[127][1] = r_cell_wire[127];							inform_L[0][0] = l_cell_wire[0];							inform_L[1][0] = l_cell_wire[1];							inform_L[2][0] = l_cell_wire[2];							inform_L[3][0] = l_cell_wire[3];							inform_L[4][0] = l_cell_wire[4];							inform_L[5][0] = l_cell_wire[5];							inform_L[6][0] = l_cell_wire[6];							inform_L[7][0] = l_cell_wire[7];							inform_L[8][0] = l_cell_wire[8];							inform_L[9][0] = l_cell_wire[9];							inform_L[10][0] = l_cell_wire[10];							inform_L[11][0] = l_cell_wire[11];							inform_L[12][0] = l_cell_wire[12];							inform_L[13][0] = l_cell_wire[13];							inform_L[14][0] = l_cell_wire[14];							inform_L[15][0] = l_cell_wire[15];							inform_L[16][0] = l_cell_wire[16];							inform_L[17][0] = l_cell_wire[17];							inform_L[18][0] = l_cell_wire[18];							inform_L[19][0] = l_cell_wire[19];							inform_L[20][0] = l_cell_wire[20];							inform_L[21][0] = l_cell_wire[21];							inform_L[22][0] = l_cell_wire[22];							inform_L[23][0] = l_cell_wire[23];							inform_L[24][0] = l_cell_wire[24];							inform_L[25][0] = l_cell_wire[25];							inform_L[26][0] = l_cell_wire[26];							inform_L[27][0] = l_cell_wire[27];							inform_L[28][0] = l_cell_wire[28];							inform_L[29][0] = l_cell_wire[29];							inform_L[30][0] = l_cell_wire[30];							inform_L[31][0] = l_cell_wire[31];							inform_L[32][0] = l_cell_wire[32];							inform_L[33][0] = l_cell_wire[33];							inform_L[34][0] = l_cell_wire[34];							inform_L[35][0] = l_cell_wire[35];							inform_L[36][0] = l_cell_wire[36];							inform_L[37][0] = l_cell_wire[37];							inform_L[38][0] = l_cell_wire[38];							inform_L[39][0] = l_cell_wire[39];							inform_L[40][0] = l_cell_wire[40];							inform_L[41][0] = l_cell_wire[41];							inform_L[42][0] = l_cell_wire[42];							inform_L[43][0] = l_cell_wire[43];							inform_L[44][0] = l_cell_wire[44];							inform_L[45][0] = l_cell_wire[45];							inform_L[46][0] = l_cell_wire[46];							inform_L[47][0] = l_cell_wire[47];							inform_L[48][0] = l_cell_wire[48];							inform_L[49][0] = l_cell_wire[49];							inform_L[50][0] = l_cell_wire[50];							inform_L[51][0] = l_cell_wire[51];							inform_L[52][0] = l_cell_wire[52];							inform_L[53][0] = l_cell_wire[53];							inform_L[54][0] = l_cell_wire[54];							inform_L[55][0] = l_cell_wire[55];							inform_L[56][0] = l_cell_wire[56];							inform_L[57][0] = l_cell_wire[57];							inform_L[58][0] = l_cell_wire[58];							inform_L[59][0] = l_cell_wire[59];							inform_L[60][0] = l_cell_wire[60];							inform_L[61][0] = l_cell_wire[61];							inform_L[62][0] = l_cell_wire[62];							inform_L[63][0] = l_cell_wire[63];							inform_L[64][0] = l_cell_wire[64];							inform_L[65][0] = l_cell_wire[65];							inform_L[66][0] = l_cell_wire[66];							inform_L[67][0] = l_cell_wire[67];							inform_L[68][0] = l_cell_wire[68];							inform_L[69][0] = l_cell_wire[69];							inform_L[70][0] = l_cell_wire[70];							inform_L[71][0] = l_cell_wire[71];							inform_L[72][0] = l_cell_wire[72];							inform_L[73][0] = l_cell_wire[73];							inform_L[74][0] = l_cell_wire[74];							inform_L[75][0] = l_cell_wire[75];							inform_L[76][0] = l_cell_wire[76];							inform_L[77][0] = l_cell_wire[77];							inform_L[78][0] = l_cell_wire[78];							inform_L[79][0] = l_cell_wire[79];							inform_L[80][0] = l_cell_wire[80];							inform_L[81][0] = l_cell_wire[81];							inform_L[82][0] = l_cell_wire[82];							inform_L[83][0] = l_cell_wire[83];							inform_L[84][0] = l_cell_wire[84];							inform_L[85][0] = l_cell_wire[85];							inform_L[86][0] = l_cell_wire[86];							inform_L[87][0] = l_cell_wire[87];							inform_L[88][0] = l_cell_wire[88];							inform_L[89][0] = l_cell_wire[89];							inform_L[90][0] = l_cell_wire[90];							inform_L[91][0] = l_cell_wire[91];							inform_L[92][0] = l_cell_wire[92];							inform_L[93][0] = l_cell_wire[93];							inform_L[94][0] = l_cell_wire[94];							inform_L[95][0] = l_cell_wire[95];							inform_L[96][0] = l_cell_wire[96];							inform_L[97][0] = l_cell_wire[97];							inform_L[98][0] = l_cell_wire[98];							inform_L[99][0] = l_cell_wire[99];							inform_L[100][0] = l_cell_wire[100];							inform_L[101][0] = l_cell_wire[101];							inform_L[102][0] = l_cell_wire[102];							inform_L[103][0] = l_cell_wire[103];							inform_L[104][0] = l_cell_wire[104];							inform_L[105][0] = l_cell_wire[105];							inform_L[106][0] = l_cell_wire[106];							inform_L[107][0] = l_cell_wire[107];							inform_L[108][0] = l_cell_wire[108];							inform_L[109][0] = l_cell_wire[109];							inform_L[110][0] = l_cell_wire[110];							inform_L[111][0] = l_cell_wire[111];							inform_L[112][0] = l_cell_wire[112];							inform_L[113][0] = l_cell_wire[113];							inform_L[114][0] = l_cell_wire[114];							inform_L[115][0] = l_cell_wire[115];							inform_L[116][0] = l_cell_wire[116];							inform_L[117][0] = l_cell_wire[117];							inform_L[118][0] = l_cell_wire[118];							inform_L[119][0] = l_cell_wire[119];							inform_L[120][0] = l_cell_wire[120];							inform_L[121][0] = l_cell_wire[121];							inform_L[122][0] = l_cell_wire[122];							inform_L[123][0] = l_cell_wire[123];							inform_L[124][0] = l_cell_wire[124];							inform_L[125][0] = l_cell_wire[125];							inform_L[126][0] = l_cell_wire[126];							inform_L[127][0] = l_cell_wire[127];						end
						2:						begin							inform_R[0][2] = r_cell_wire[0];							inform_R[2][2] = r_cell_wire[1];							inform_R[1][2] = r_cell_wire[2];							inform_R[3][2] = r_cell_wire[3];							inform_R[4][2] = r_cell_wire[4];							inform_R[6][2] = r_cell_wire[5];							inform_R[5][2] = r_cell_wire[6];							inform_R[7][2] = r_cell_wire[7];							inform_R[8][2] = r_cell_wire[8];							inform_R[10][2] = r_cell_wire[9];							inform_R[9][2] = r_cell_wire[10];							inform_R[11][2] = r_cell_wire[11];							inform_R[12][2] = r_cell_wire[12];							inform_R[14][2] = r_cell_wire[13];							inform_R[13][2] = r_cell_wire[14];							inform_R[15][2] = r_cell_wire[15];							inform_R[16][2] = r_cell_wire[16];							inform_R[18][2] = r_cell_wire[17];							inform_R[17][2] = r_cell_wire[18];							inform_R[19][2] = r_cell_wire[19];							inform_R[20][2] = r_cell_wire[20];							inform_R[22][2] = r_cell_wire[21];							inform_R[21][2] = r_cell_wire[22];							inform_R[23][2] = r_cell_wire[23];							inform_R[24][2] = r_cell_wire[24];							inform_R[26][2] = r_cell_wire[25];							inform_R[25][2] = r_cell_wire[26];							inform_R[27][2] = r_cell_wire[27];							inform_R[28][2] = r_cell_wire[28];							inform_R[30][2] = r_cell_wire[29];							inform_R[29][2] = r_cell_wire[30];							inform_R[31][2] = r_cell_wire[31];							inform_R[32][2] = r_cell_wire[32];							inform_R[34][2] = r_cell_wire[33];							inform_R[33][2] = r_cell_wire[34];							inform_R[35][2] = r_cell_wire[35];							inform_R[36][2] = r_cell_wire[36];							inform_R[38][2] = r_cell_wire[37];							inform_R[37][2] = r_cell_wire[38];							inform_R[39][2] = r_cell_wire[39];							inform_R[40][2] = r_cell_wire[40];							inform_R[42][2] = r_cell_wire[41];							inform_R[41][2] = r_cell_wire[42];							inform_R[43][2] = r_cell_wire[43];							inform_R[44][2] = r_cell_wire[44];							inform_R[46][2] = r_cell_wire[45];							inform_R[45][2] = r_cell_wire[46];							inform_R[47][2] = r_cell_wire[47];							inform_R[48][2] = r_cell_wire[48];							inform_R[50][2] = r_cell_wire[49];							inform_R[49][2] = r_cell_wire[50];							inform_R[51][2] = r_cell_wire[51];							inform_R[52][2] = r_cell_wire[52];							inform_R[54][2] = r_cell_wire[53];							inform_R[53][2] = r_cell_wire[54];							inform_R[55][2] = r_cell_wire[55];							inform_R[56][2] = r_cell_wire[56];							inform_R[58][2] = r_cell_wire[57];							inform_R[57][2] = r_cell_wire[58];							inform_R[59][2] = r_cell_wire[59];							inform_R[60][2] = r_cell_wire[60];							inform_R[62][2] = r_cell_wire[61];							inform_R[61][2] = r_cell_wire[62];							inform_R[63][2] = r_cell_wire[63];							inform_R[64][2] = r_cell_wire[64];							inform_R[66][2] = r_cell_wire[65];							inform_R[65][2] = r_cell_wire[66];							inform_R[67][2] = r_cell_wire[67];							inform_R[68][2] = r_cell_wire[68];							inform_R[70][2] = r_cell_wire[69];							inform_R[69][2] = r_cell_wire[70];							inform_R[71][2] = r_cell_wire[71];							inform_R[72][2] = r_cell_wire[72];							inform_R[74][2] = r_cell_wire[73];							inform_R[73][2] = r_cell_wire[74];							inform_R[75][2] = r_cell_wire[75];							inform_R[76][2] = r_cell_wire[76];							inform_R[78][2] = r_cell_wire[77];							inform_R[77][2] = r_cell_wire[78];							inform_R[79][2] = r_cell_wire[79];							inform_R[80][2] = r_cell_wire[80];							inform_R[82][2] = r_cell_wire[81];							inform_R[81][2] = r_cell_wire[82];							inform_R[83][2] = r_cell_wire[83];							inform_R[84][2] = r_cell_wire[84];							inform_R[86][2] = r_cell_wire[85];							inform_R[85][2] = r_cell_wire[86];							inform_R[87][2] = r_cell_wire[87];							inform_R[88][2] = r_cell_wire[88];							inform_R[90][2] = r_cell_wire[89];							inform_R[89][2] = r_cell_wire[90];							inform_R[91][2] = r_cell_wire[91];							inform_R[92][2] = r_cell_wire[92];							inform_R[94][2] = r_cell_wire[93];							inform_R[93][2] = r_cell_wire[94];							inform_R[95][2] = r_cell_wire[95];							inform_R[96][2] = r_cell_wire[96];							inform_R[98][2] = r_cell_wire[97];							inform_R[97][2] = r_cell_wire[98];							inform_R[99][2] = r_cell_wire[99];							inform_R[100][2] = r_cell_wire[100];							inform_R[102][2] = r_cell_wire[101];							inform_R[101][2] = r_cell_wire[102];							inform_R[103][2] = r_cell_wire[103];							inform_R[104][2] = r_cell_wire[104];							inform_R[106][2] = r_cell_wire[105];							inform_R[105][2] = r_cell_wire[106];							inform_R[107][2] = r_cell_wire[107];							inform_R[108][2] = r_cell_wire[108];							inform_R[110][2] = r_cell_wire[109];							inform_R[109][2] = r_cell_wire[110];							inform_R[111][2] = r_cell_wire[111];							inform_R[112][2] = r_cell_wire[112];							inform_R[114][2] = r_cell_wire[113];							inform_R[113][2] = r_cell_wire[114];							inform_R[115][2] = r_cell_wire[115];							inform_R[116][2] = r_cell_wire[116];							inform_R[118][2] = r_cell_wire[117];							inform_R[117][2] = r_cell_wire[118];							inform_R[119][2] = r_cell_wire[119];							inform_R[120][2] = r_cell_wire[120];							inform_R[122][2] = r_cell_wire[121];							inform_R[121][2] = r_cell_wire[122];							inform_R[123][2] = r_cell_wire[123];							inform_R[124][2] = r_cell_wire[124];							inform_R[126][2] = r_cell_wire[125];							inform_R[125][2] = r_cell_wire[126];							inform_R[127][2] = r_cell_wire[127];							inform_L[0][1] = l_cell_wire[0];							inform_L[2][1] = l_cell_wire[1];							inform_L[1][1] = l_cell_wire[2];							inform_L[3][1] = l_cell_wire[3];							inform_L[4][1] = l_cell_wire[4];							inform_L[6][1] = l_cell_wire[5];							inform_L[5][1] = l_cell_wire[6];							inform_L[7][1] = l_cell_wire[7];							inform_L[8][1] = l_cell_wire[8];							inform_L[10][1] = l_cell_wire[9];							inform_L[9][1] = l_cell_wire[10];							inform_L[11][1] = l_cell_wire[11];							inform_L[12][1] = l_cell_wire[12];							inform_L[14][1] = l_cell_wire[13];							inform_L[13][1] = l_cell_wire[14];							inform_L[15][1] = l_cell_wire[15];							inform_L[16][1] = l_cell_wire[16];							inform_L[18][1] = l_cell_wire[17];							inform_L[17][1] = l_cell_wire[18];							inform_L[19][1] = l_cell_wire[19];							inform_L[20][1] = l_cell_wire[20];							inform_L[22][1] = l_cell_wire[21];							inform_L[21][1] = l_cell_wire[22];							inform_L[23][1] = l_cell_wire[23];							inform_L[24][1] = l_cell_wire[24];							inform_L[26][1] = l_cell_wire[25];							inform_L[25][1] = l_cell_wire[26];							inform_L[27][1] = l_cell_wire[27];							inform_L[28][1] = l_cell_wire[28];							inform_L[30][1] = l_cell_wire[29];							inform_L[29][1] = l_cell_wire[30];							inform_L[31][1] = l_cell_wire[31];							inform_L[32][1] = l_cell_wire[32];							inform_L[34][1] = l_cell_wire[33];							inform_L[33][1] = l_cell_wire[34];							inform_L[35][1] = l_cell_wire[35];							inform_L[36][1] = l_cell_wire[36];							inform_L[38][1] = l_cell_wire[37];							inform_L[37][1] = l_cell_wire[38];							inform_L[39][1] = l_cell_wire[39];							inform_L[40][1] = l_cell_wire[40];							inform_L[42][1] = l_cell_wire[41];							inform_L[41][1] = l_cell_wire[42];							inform_L[43][1] = l_cell_wire[43];							inform_L[44][1] = l_cell_wire[44];							inform_L[46][1] = l_cell_wire[45];							inform_L[45][1] = l_cell_wire[46];							inform_L[47][1] = l_cell_wire[47];							inform_L[48][1] = l_cell_wire[48];							inform_L[50][1] = l_cell_wire[49];							inform_L[49][1] = l_cell_wire[50];							inform_L[51][1] = l_cell_wire[51];							inform_L[52][1] = l_cell_wire[52];							inform_L[54][1] = l_cell_wire[53];							inform_L[53][1] = l_cell_wire[54];							inform_L[55][1] = l_cell_wire[55];							inform_L[56][1] = l_cell_wire[56];							inform_L[58][1] = l_cell_wire[57];							inform_L[57][1] = l_cell_wire[58];							inform_L[59][1] = l_cell_wire[59];							inform_L[60][1] = l_cell_wire[60];							inform_L[62][1] = l_cell_wire[61];							inform_L[61][1] = l_cell_wire[62];							inform_L[63][1] = l_cell_wire[63];							inform_L[64][1] = l_cell_wire[64];							inform_L[66][1] = l_cell_wire[65];							inform_L[65][1] = l_cell_wire[66];							inform_L[67][1] = l_cell_wire[67];							inform_L[68][1] = l_cell_wire[68];							inform_L[70][1] = l_cell_wire[69];							inform_L[69][1] = l_cell_wire[70];							inform_L[71][1] = l_cell_wire[71];							inform_L[72][1] = l_cell_wire[72];							inform_L[74][1] = l_cell_wire[73];							inform_L[73][1] = l_cell_wire[74];							inform_L[75][1] = l_cell_wire[75];							inform_L[76][1] = l_cell_wire[76];							inform_L[78][1] = l_cell_wire[77];							inform_L[77][1] = l_cell_wire[78];							inform_L[79][1] = l_cell_wire[79];							inform_L[80][1] = l_cell_wire[80];							inform_L[82][1] = l_cell_wire[81];							inform_L[81][1] = l_cell_wire[82];							inform_L[83][1] = l_cell_wire[83];							inform_L[84][1] = l_cell_wire[84];							inform_L[86][1] = l_cell_wire[85];							inform_L[85][1] = l_cell_wire[86];							inform_L[87][1] = l_cell_wire[87];							inform_L[88][1] = l_cell_wire[88];							inform_L[90][1] = l_cell_wire[89];							inform_L[89][1] = l_cell_wire[90];							inform_L[91][1] = l_cell_wire[91];							inform_L[92][1] = l_cell_wire[92];							inform_L[94][1] = l_cell_wire[93];							inform_L[93][1] = l_cell_wire[94];							inform_L[95][1] = l_cell_wire[95];							inform_L[96][1] = l_cell_wire[96];							inform_L[98][1] = l_cell_wire[97];							inform_L[97][1] = l_cell_wire[98];							inform_L[99][1] = l_cell_wire[99];							inform_L[100][1] = l_cell_wire[100];							inform_L[102][1] = l_cell_wire[101];							inform_L[101][1] = l_cell_wire[102];							inform_L[103][1] = l_cell_wire[103];							inform_L[104][1] = l_cell_wire[104];							inform_L[106][1] = l_cell_wire[105];							inform_L[105][1] = l_cell_wire[106];							inform_L[107][1] = l_cell_wire[107];							inform_L[108][1] = l_cell_wire[108];							inform_L[110][1] = l_cell_wire[109];							inform_L[109][1] = l_cell_wire[110];							inform_L[111][1] = l_cell_wire[111];							inform_L[112][1] = l_cell_wire[112];							inform_L[114][1] = l_cell_wire[113];							inform_L[113][1] = l_cell_wire[114];							inform_L[115][1] = l_cell_wire[115];							inform_L[116][1] = l_cell_wire[116];							inform_L[118][1] = l_cell_wire[117];							inform_L[117][1] = l_cell_wire[118];							inform_L[119][1] = l_cell_wire[119];							inform_L[120][1] = l_cell_wire[120];							inform_L[122][1] = l_cell_wire[121];							inform_L[121][1] = l_cell_wire[122];							inform_L[123][1] = l_cell_wire[123];							inform_L[124][1] = l_cell_wire[124];							inform_L[126][1] = l_cell_wire[125];							inform_L[125][1] = l_cell_wire[126];							inform_L[127][1] = l_cell_wire[127];						end
						3:						begin							inform_R[0][3] = r_cell_wire[0];							inform_R[4][3] = r_cell_wire[1];							inform_R[1][3] = r_cell_wire[2];							inform_R[5][3] = r_cell_wire[3];							inform_R[2][3] = r_cell_wire[4];							inform_R[6][3] = r_cell_wire[5];							inform_R[3][3] = r_cell_wire[6];							inform_R[7][3] = r_cell_wire[7];							inform_R[8][3] = r_cell_wire[8];							inform_R[12][3] = r_cell_wire[9];							inform_R[9][3] = r_cell_wire[10];							inform_R[13][3] = r_cell_wire[11];							inform_R[10][3] = r_cell_wire[12];							inform_R[14][3] = r_cell_wire[13];							inform_R[11][3] = r_cell_wire[14];							inform_R[15][3] = r_cell_wire[15];							inform_R[16][3] = r_cell_wire[16];							inform_R[20][3] = r_cell_wire[17];							inform_R[17][3] = r_cell_wire[18];							inform_R[21][3] = r_cell_wire[19];							inform_R[18][3] = r_cell_wire[20];							inform_R[22][3] = r_cell_wire[21];							inform_R[19][3] = r_cell_wire[22];							inform_R[23][3] = r_cell_wire[23];							inform_R[24][3] = r_cell_wire[24];							inform_R[28][3] = r_cell_wire[25];							inform_R[25][3] = r_cell_wire[26];							inform_R[29][3] = r_cell_wire[27];							inform_R[26][3] = r_cell_wire[28];							inform_R[30][3] = r_cell_wire[29];							inform_R[27][3] = r_cell_wire[30];							inform_R[31][3] = r_cell_wire[31];							inform_R[32][3] = r_cell_wire[32];							inform_R[36][3] = r_cell_wire[33];							inform_R[33][3] = r_cell_wire[34];							inform_R[37][3] = r_cell_wire[35];							inform_R[34][3] = r_cell_wire[36];							inform_R[38][3] = r_cell_wire[37];							inform_R[35][3] = r_cell_wire[38];							inform_R[39][3] = r_cell_wire[39];							inform_R[40][3] = r_cell_wire[40];							inform_R[44][3] = r_cell_wire[41];							inform_R[41][3] = r_cell_wire[42];							inform_R[45][3] = r_cell_wire[43];							inform_R[42][3] = r_cell_wire[44];							inform_R[46][3] = r_cell_wire[45];							inform_R[43][3] = r_cell_wire[46];							inform_R[47][3] = r_cell_wire[47];							inform_R[48][3] = r_cell_wire[48];							inform_R[52][3] = r_cell_wire[49];							inform_R[49][3] = r_cell_wire[50];							inform_R[53][3] = r_cell_wire[51];							inform_R[50][3] = r_cell_wire[52];							inform_R[54][3] = r_cell_wire[53];							inform_R[51][3] = r_cell_wire[54];							inform_R[55][3] = r_cell_wire[55];							inform_R[56][3] = r_cell_wire[56];							inform_R[60][3] = r_cell_wire[57];							inform_R[57][3] = r_cell_wire[58];							inform_R[61][3] = r_cell_wire[59];							inform_R[58][3] = r_cell_wire[60];							inform_R[62][3] = r_cell_wire[61];							inform_R[59][3] = r_cell_wire[62];							inform_R[63][3] = r_cell_wire[63];							inform_R[64][3] = r_cell_wire[64];							inform_R[68][3] = r_cell_wire[65];							inform_R[65][3] = r_cell_wire[66];							inform_R[69][3] = r_cell_wire[67];							inform_R[66][3] = r_cell_wire[68];							inform_R[70][3] = r_cell_wire[69];							inform_R[67][3] = r_cell_wire[70];							inform_R[71][3] = r_cell_wire[71];							inform_R[72][3] = r_cell_wire[72];							inform_R[76][3] = r_cell_wire[73];							inform_R[73][3] = r_cell_wire[74];							inform_R[77][3] = r_cell_wire[75];							inform_R[74][3] = r_cell_wire[76];							inform_R[78][3] = r_cell_wire[77];							inform_R[75][3] = r_cell_wire[78];							inform_R[79][3] = r_cell_wire[79];							inform_R[80][3] = r_cell_wire[80];							inform_R[84][3] = r_cell_wire[81];							inform_R[81][3] = r_cell_wire[82];							inform_R[85][3] = r_cell_wire[83];							inform_R[82][3] = r_cell_wire[84];							inform_R[86][3] = r_cell_wire[85];							inform_R[83][3] = r_cell_wire[86];							inform_R[87][3] = r_cell_wire[87];							inform_R[88][3] = r_cell_wire[88];							inform_R[92][3] = r_cell_wire[89];							inform_R[89][3] = r_cell_wire[90];							inform_R[93][3] = r_cell_wire[91];							inform_R[90][3] = r_cell_wire[92];							inform_R[94][3] = r_cell_wire[93];							inform_R[91][3] = r_cell_wire[94];							inform_R[95][3] = r_cell_wire[95];							inform_R[96][3] = r_cell_wire[96];							inform_R[100][3] = r_cell_wire[97];							inform_R[97][3] = r_cell_wire[98];							inform_R[101][3] = r_cell_wire[99];							inform_R[98][3] = r_cell_wire[100];							inform_R[102][3] = r_cell_wire[101];							inform_R[99][3] = r_cell_wire[102];							inform_R[103][3] = r_cell_wire[103];							inform_R[104][3] = r_cell_wire[104];							inform_R[108][3] = r_cell_wire[105];							inform_R[105][3] = r_cell_wire[106];							inform_R[109][3] = r_cell_wire[107];							inform_R[106][3] = r_cell_wire[108];							inform_R[110][3] = r_cell_wire[109];							inform_R[107][3] = r_cell_wire[110];							inform_R[111][3] = r_cell_wire[111];							inform_R[112][3] = r_cell_wire[112];							inform_R[116][3] = r_cell_wire[113];							inform_R[113][3] = r_cell_wire[114];							inform_R[117][3] = r_cell_wire[115];							inform_R[114][3] = r_cell_wire[116];							inform_R[118][3] = r_cell_wire[117];							inform_R[115][3] = r_cell_wire[118];							inform_R[119][3] = r_cell_wire[119];							inform_R[120][3] = r_cell_wire[120];							inform_R[124][3] = r_cell_wire[121];							inform_R[121][3] = r_cell_wire[122];							inform_R[125][3] = r_cell_wire[123];							inform_R[122][3] = r_cell_wire[124];							inform_R[126][3] = r_cell_wire[125];							inform_R[123][3] = r_cell_wire[126];							inform_R[127][3] = r_cell_wire[127];							inform_L[0][2] = l_cell_wire[0];							inform_L[4][2] = l_cell_wire[1];							inform_L[1][2] = l_cell_wire[2];							inform_L[5][2] = l_cell_wire[3];							inform_L[2][2] = l_cell_wire[4];							inform_L[6][2] = l_cell_wire[5];							inform_L[3][2] = l_cell_wire[6];							inform_L[7][2] = l_cell_wire[7];							inform_L[8][2] = l_cell_wire[8];							inform_L[12][2] = l_cell_wire[9];							inform_L[9][2] = l_cell_wire[10];							inform_L[13][2] = l_cell_wire[11];							inform_L[10][2] = l_cell_wire[12];							inform_L[14][2] = l_cell_wire[13];							inform_L[11][2] = l_cell_wire[14];							inform_L[15][2] = l_cell_wire[15];							inform_L[16][2] = l_cell_wire[16];							inform_L[20][2] = l_cell_wire[17];							inform_L[17][2] = l_cell_wire[18];							inform_L[21][2] = l_cell_wire[19];							inform_L[18][2] = l_cell_wire[20];							inform_L[22][2] = l_cell_wire[21];							inform_L[19][2] = l_cell_wire[22];							inform_L[23][2] = l_cell_wire[23];							inform_L[24][2] = l_cell_wire[24];							inform_L[28][2] = l_cell_wire[25];							inform_L[25][2] = l_cell_wire[26];							inform_L[29][2] = l_cell_wire[27];							inform_L[26][2] = l_cell_wire[28];							inform_L[30][2] = l_cell_wire[29];							inform_L[27][2] = l_cell_wire[30];							inform_L[31][2] = l_cell_wire[31];							inform_L[32][2] = l_cell_wire[32];							inform_L[36][2] = l_cell_wire[33];							inform_L[33][2] = l_cell_wire[34];							inform_L[37][2] = l_cell_wire[35];							inform_L[34][2] = l_cell_wire[36];							inform_L[38][2] = l_cell_wire[37];							inform_L[35][2] = l_cell_wire[38];							inform_L[39][2] = l_cell_wire[39];							inform_L[40][2] = l_cell_wire[40];							inform_L[44][2] = l_cell_wire[41];							inform_L[41][2] = l_cell_wire[42];							inform_L[45][2] = l_cell_wire[43];							inform_L[42][2] = l_cell_wire[44];							inform_L[46][2] = l_cell_wire[45];							inform_L[43][2] = l_cell_wire[46];							inform_L[47][2] = l_cell_wire[47];							inform_L[48][2] = l_cell_wire[48];							inform_L[52][2] = l_cell_wire[49];							inform_L[49][2] = l_cell_wire[50];							inform_L[53][2] = l_cell_wire[51];							inform_L[50][2] = l_cell_wire[52];							inform_L[54][2] = l_cell_wire[53];							inform_L[51][2] = l_cell_wire[54];							inform_L[55][2] = l_cell_wire[55];							inform_L[56][2] = l_cell_wire[56];							inform_L[60][2] = l_cell_wire[57];							inform_L[57][2] = l_cell_wire[58];							inform_L[61][2] = l_cell_wire[59];							inform_L[58][2] = l_cell_wire[60];							inform_L[62][2] = l_cell_wire[61];							inform_L[59][2] = l_cell_wire[62];							inform_L[63][2] = l_cell_wire[63];							inform_L[64][2] = l_cell_wire[64];							inform_L[68][2] = l_cell_wire[65];							inform_L[65][2] = l_cell_wire[66];							inform_L[69][2] = l_cell_wire[67];							inform_L[66][2] = l_cell_wire[68];							inform_L[70][2] = l_cell_wire[69];							inform_L[67][2] = l_cell_wire[70];							inform_L[71][2] = l_cell_wire[71];							inform_L[72][2] = l_cell_wire[72];							inform_L[76][2] = l_cell_wire[73];							inform_L[73][2] = l_cell_wire[74];							inform_L[77][2] = l_cell_wire[75];							inform_L[74][2] = l_cell_wire[76];							inform_L[78][2] = l_cell_wire[77];							inform_L[75][2] = l_cell_wire[78];							inform_L[79][2] = l_cell_wire[79];							inform_L[80][2] = l_cell_wire[80];							inform_L[84][2] = l_cell_wire[81];							inform_L[81][2] = l_cell_wire[82];							inform_L[85][2] = l_cell_wire[83];							inform_L[82][2] = l_cell_wire[84];							inform_L[86][2] = l_cell_wire[85];							inform_L[83][2] = l_cell_wire[86];							inform_L[87][2] = l_cell_wire[87];							inform_L[88][2] = l_cell_wire[88];							inform_L[92][2] = l_cell_wire[89];							inform_L[89][2] = l_cell_wire[90];							inform_L[93][2] = l_cell_wire[91];							inform_L[90][2] = l_cell_wire[92];							inform_L[94][2] = l_cell_wire[93];							inform_L[91][2] = l_cell_wire[94];							inform_L[95][2] = l_cell_wire[95];							inform_L[96][2] = l_cell_wire[96];							inform_L[100][2] = l_cell_wire[97];							inform_L[97][2] = l_cell_wire[98];							inform_L[101][2] = l_cell_wire[99];							inform_L[98][2] = l_cell_wire[100];							inform_L[102][2] = l_cell_wire[101];							inform_L[99][2] = l_cell_wire[102];							inform_L[103][2] = l_cell_wire[103];							inform_L[104][2] = l_cell_wire[104];							inform_L[108][2] = l_cell_wire[105];							inform_L[105][2] = l_cell_wire[106];							inform_L[109][2] = l_cell_wire[107];							inform_L[106][2] = l_cell_wire[108];							inform_L[110][2] = l_cell_wire[109];							inform_L[107][2] = l_cell_wire[110];							inform_L[111][2] = l_cell_wire[111];							inform_L[112][2] = l_cell_wire[112];							inform_L[116][2] = l_cell_wire[113];							inform_L[113][2] = l_cell_wire[114];							inform_L[117][2] = l_cell_wire[115];							inform_L[114][2] = l_cell_wire[116];							inform_L[118][2] = l_cell_wire[117];							inform_L[115][2] = l_cell_wire[118];							inform_L[119][2] = l_cell_wire[119];							inform_L[120][2] = l_cell_wire[120];							inform_L[124][2] = l_cell_wire[121];							inform_L[121][2] = l_cell_wire[122];							inform_L[125][2] = l_cell_wire[123];							inform_L[122][2] = l_cell_wire[124];							inform_L[126][2] = l_cell_wire[125];							inform_L[123][2] = l_cell_wire[126];							inform_L[127][2] = l_cell_wire[127];						end
						4:						begin							inform_R[0][4] = r_cell_wire[0];							inform_R[8][4] = r_cell_wire[1];							inform_R[1][4] = r_cell_wire[2];							inform_R[9][4] = r_cell_wire[3];							inform_R[2][4] = r_cell_wire[4];							inform_R[10][4] = r_cell_wire[5];							inform_R[3][4] = r_cell_wire[6];							inform_R[11][4] = r_cell_wire[7];							inform_R[4][4] = r_cell_wire[8];							inform_R[12][4] = r_cell_wire[9];							inform_R[5][4] = r_cell_wire[10];							inform_R[13][4] = r_cell_wire[11];							inform_R[6][4] = r_cell_wire[12];							inform_R[14][4] = r_cell_wire[13];							inform_R[7][4] = r_cell_wire[14];							inform_R[15][4] = r_cell_wire[15];							inform_R[16][4] = r_cell_wire[16];							inform_R[24][4] = r_cell_wire[17];							inform_R[17][4] = r_cell_wire[18];							inform_R[25][4] = r_cell_wire[19];							inform_R[18][4] = r_cell_wire[20];							inform_R[26][4] = r_cell_wire[21];							inform_R[19][4] = r_cell_wire[22];							inform_R[27][4] = r_cell_wire[23];							inform_R[20][4] = r_cell_wire[24];							inform_R[28][4] = r_cell_wire[25];							inform_R[21][4] = r_cell_wire[26];							inform_R[29][4] = r_cell_wire[27];							inform_R[22][4] = r_cell_wire[28];							inform_R[30][4] = r_cell_wire[29];							inform_R[23][4] = r_cell_wire[30];							inform_R[31][4] = r_cell_wire[31];							inform_R[32][4] = r_cell_wire[32];							inform_R[40][4] = r_cell_wire[33];							inform_R[33][4] = r_cell_wire[34];							inform_R[41][4] = r_cell_wire[35];							inform_R[34][4] = r_cell_wire[36];							inform_R[42][4] = r_cell_wire[37];							inform_R[35][4] = r_cell_wire[38];							inform_R[43][4] = r_cell_wire[39];							inform_R[36][4] = r_cell_wire[40];							inform_R[44][4] = r_cell_wire[41];							inform_R[37][4] = r_cell_wire[42];							inform_R[45][4] = r_cell_wire[43];							inform_R[38][4] = r_cell_wire[44];							inform_R[46][4] = r_cell_wire[45];							inform_R[39][4] = r_cell_wire[46];							inform_R[47][4] = r_cell_wire[47];							inform_R[48][4] = r_cell_wire[48];							inform_R[56][4] = r_cell_wire[49];							inform_R[49][4] = r_cell_wire[50];							inform_R[57][4] = r_cell_wire[51];							inform_R[50][4] = r_cell_wire[52];							inform_R[58][4] = r_cell_wire[53];							inform_R[51][4] = r_cell_wire[54];							inform_R[59][4] = r_cell_wire[55];							inform_R[52][4] = r_cell_wire[56];							inform_R[60][4] = r_cell_wire[57];							inform_R[53][4] = r_cell_wire[58];							inform_R[61][4] = r_cell_wire[59];							inform_R[54][4] = r_cell_wire[60];							inform_R[62][4] = r_cell_wire[61];							inform_R[55][4] = r_cell_wire[62];							inform_R[63][4] = r_cell_wire[63];							inform_R[64][4] = r_cell_wire[64];							inform_R[72][4] = r_cell_wire[65];							inform_R[65][4] = r_cell_wire[66];							inform_R[73][4] = r_cell_wire[67];							inform_R[66][4] = r_cell_wire[68];							inform_R[74][4] = r_cell_wire[69];							inform_R[67][4] = r_cell_wire[70];							inform_R[75][4] = r_cell_wire[71];							inform_R[68][4] = r_cell_wire[72];							inform_R[76][4] = r_cell_wire[73];							inform_R[69][4] = r_cell_wire[74];							inform_R[77][4] = r_cell_wire[75];							inform_R[70][4] = r_cell_wire[76];							inform_R[78][4] = r_cell_wire[77];							inform_R[71][4] = r_cell_wire[78];							inform_R[79][4] = r_cell_wire[79];							inform_R[80][4] = r_cell_wire[80];							inform_R[88][4] = r_cell_wire[81];							inform_R[81][4] = r_cell_wire[82];							inform_R[89][4] = r_cell_wire[83];							inform_R[82][4] = r_cell_wire[84];							inform_R[90][4] = r_cell_wire[85];							inform_R[83][4] = r_cell_wire[86];							inform_R[91][4] = r_cell_wire[87];							inform_R[84][4] = r_cell_wire[88];							inform_R[92][4] = r_cell_wire[89];							inform_R[85][4] = r_cell_wire[90];							inform_R[93][4] = r_cell_wire[91];							inform_R[86][4] = r_cell_wire[92];							inform_R[94][4] = r_cell_wire[93];							inform_R[87][4] = r_cell_wire[94];							inform_R[95][4] = r_cell_wire[95];							inform_R[96][4] = r_cell_wire[96];							inform_R[104][4] = r_cell_wire[97];							inform_R[97][4] = r_cell_wire[98];							inform_R[105][4] = r_cell_wire[99];							inform_R[98][4] = r_cell_wire[100];							inform_R[106][4] = r_cell_wire[101];							inform_R[99][4] = r_cell_wire[102];							inform_R[107][4] = r_cell_wire[103];							inform_R[100][4] = r_cell_wire[104];							inform_R[108][4] = r_cell_wire[105];							inform_R[101][4] = r_cell_wire[106];							inform_R[109][4] = r_cell_wire[107];							inform_R[102][4] = r_cell_wire[108];							inform_R[110][4] = r_cell_wire[109];							inform_R[103][4] = r_cell_wire[110];							inform_R[111][4] = r_cell_wire[111];							inform_R[112][4] = r_cell_wire[112];							inform_R[120][4] = r_cell_wire[113];							inform_R[113][4] = r_cell_wire[114];							inform_R[121][4] = r_cell_wire[115];							inform_R[114][4] = r_cell_wire[116];							inform_R[122][4] = r_cell_wire[117];							inform_R[115][4] = r_cell_wire[118];							inform_R[123][4] = r_cell_wire[119];							inform_R[116][4] = r_cell_wire[120];							inform_R[124][4] = r_cell_wire[121];							inform_R[117][4] = r_cell_wire[122];							inform_R[125][4] = r_cell_wire[123];							inform_R[118][4] = r_cell_wire[124];							inform_R[126][4] = r_cell_wire[125];							inform_R[119][4] = r_cell_wire[126];							inform_R[127][4] = r_cell_wire[127];							inform_L[0][3] = l_cell_wire[0];							inform_L[8][3] = l_cell_wire[1];							inform_L[1][3] = l_cell_wire[2];							inform_L[9][3] = l_cell_wire[3];							inform_L[2][3] = l_cell_wire[4];							inform_L[10][3] = l_cell_wire[5];							inform_L[3][3] = l_cell_wire[6];							inform_L[11][3] = l_cell_wire[7];							inform_L[4][3] = l_cell_wire[8];							inform_L[12][3] = l_cell_wire[9];							inform_L[5][3] = l_cell_wire[10];							inform_L[13][3] = l_cell_wire[11];							inform_L[6][3] = l_cell_wire[12];							inform_L[14][3] = l_cell_wire[13];							inform_L[7][3] = l_cell_wire[14];							inform_L[15][3] = l_cell_wire[15];							inform_L[16][3] = l_cell_wire[16];							inform_L[24][3] = l_cell_wire[17];							inform_L[17][3] = l_cell_wire[18];							inform_L[25][3] = l_cell_wire[19];							inform_L[18][3] = l_cell_wire[20];							inform_L[26][3] = l_cell_wire[21];							inform_L[19][3] = l_cell_wire[22];							inform_L[27][3] = l_cell_wire[23];							inform_L[20][3] = l_cell_wire[24];							inform_L[28][3] = l_cell_wire[25];							inform_L[21][3] = l_cell_wire[26];							inform_L[29][3] = l_cell_wire[27];							inform_L[22][3] = l_cell_wire[28];							inform_L[30][3] = l_cell_wire[29];							inform_L[23][3] = l_cell_wire[30];							inform_L[31][3] = l_cell_wire[31];							inform_L[32][3] = l_cell_wire[32];							inform_L[40][3] = l_cell_wire[33];							inform_L[33][3] = l_cell_wire[34];							inform_L[41][3] = l_cell_wire[35];							inform_L[34][3] = l_cell_wire[36];							inform_L[42][3] = l_cell_wire[37];							inform_L[35][3] = l_cell_wire[38];							inform_L[43][3] = l_cell_wire[39];							inform_L[36][3] = l_cell_wire[40];							inform_L[44][3] = l_cell_wire[41];							inform_L[37][3] = l_cell_wire[42];							inform_L[45][3] = l_cell_wire[43];							inform_L[38][3] = l_cell_wire[44];							inform_L[46][3] = l_cell_wire[45];							inform_L[39][3] = l_cell_wire[46];							inform_L[47][3] = l_cell_wire[47];							inform_L[48][3] = l_cell_wire[48];							inform_L[56][3] = l_cell_wire[49];							inform_L[49][3] = l_cell_wire[50];							inform_L[57][3] = l_cell_wire[51];							inform_L[50][3] = l_cell_wire[52];							inform_L[58][3] = l_cell_wire[53];							inform_L[51][3] = l_cell_wire[54];							inform_L[59][3] = l_cell_wire[55];							inform_L[52][3] = l_cell_wire[56];							inform_L[60][3] = l_cell_wire[57];							inform_L[53][3] = l_cell_wire[58];							inform_L[61][3] = l_cell_wire[59];							inform_L[54][3] = l_cell_wire[60];							inform_L[62][3] = l_cell_wire[61];							inform_L[55][3] = l_cell_wire[62];							inform_L[63][3] = l_cell_wire[63];							inform_L[64][3] = l_cell_wire[64];							inform_L[72][3] = l_cell_wire[65];							inform_L[65][3] = l_cell_wire[66];							inform_L[73][3] = l_cell_wire[67];							inform_L[66][3] = l_cell_wire[68];							inform_L[74][3] = l_cell_wire[69];							inform_L[67][3] = l_cell_wire[70];							inform_L[75][3] = l_cell_wire[71];							inform_L[68][3] = l_cell_wire[72];							inform_L[76][3] = l_cell_wire[73];							inform_L[69][3] = l_cell_wire[74];							inform_L[77][3] = l_cell_wire[75];							inform_L[70][3] = l_cell_wire[76];							inform_L[78][3] = l_cell_wire[77];							inform_L[71][3] = l_cell_wire[78];							inform_L[79][3] = l_cell_wire[79];							inform_L[80][3] = l_cell_wire[80];							inform_L[88][3] = l_cell_wire[81];							inform_L[81][3] = l_cell_wire[82];							inform_L[89][3] = l_cell_wire[83];							inform_L[82][3] = l_cell_wire[84];							inform_L[90][3] = l_cell_wire[85];							inform_L[83][3] = l_cell_wire[86];							inform_L[91][3] = l_cell_wire[87];							inform_L[84][3] = l_cell_wire[88];							inform_L[92][3] = l_cell_wire[89];							inform_L[85][3] = l_cell_wire[90];							inform_L[93][3] = l_cell_wire[91];							inform_L[86][3] = l_cell_wire[92];							inform_L[94][3] = l_cell_wire[93];							inform_L[87][3] = l_cell_wire[94];							inform_L[95][3] = l_cell_wire[95];							inform_L[96][3] = l_cell_wire[96];							inform_L[104][3] = l_cell_wire[97];							inform_L[97][3] = l_cell_wire[98];							inform_L[105][3] = l_cell_wire[99];							inform_L[98][3] = l_cell_wire[100];							inform_L[106][3] = l_cell_wire[101];							inform_L[99][3] = l_cell_wire[102];							inform_L[107][3] = l_cell_wire[103];							inform_L[100][3] = l_cell_wire[104];							inform_L[108][3] = l_cell_wire[105];							inform_L[101][3] = l_cell_wire[106];							inform_L[109][3] = l_cell_wire[107];							inform_L[102][3] = l_cell_wire[108];							inform_L[110][3] = l_cell_wire[109];							inform_L[103][3] = l_cell_wire[110];							inform_L[111][3] = l_cell_wire[111];							inform_L[112][3] = l_cell_wire[112];							inform_L[120][3] = l_cell_wire[113];							inform_L[113][3] = l_cell_wire[114];							inform_L[121][3] = l_cell_wire[115];							inform_L[114][3] = l_cell_wire[116];							inform_L[122][3] = l_cell_wire[117];							inform_L[115][3] = l_cell_wire[118];							inform_L[123][3] = l_cell_wire[119];							inform_L[116][3] = l_cell_wire[120];							inform_L[124][3] = l_cell_wire[121];							inform_L[117][3] = l_cell_wire[122];							inform_L[125][3] = l_cell_wire[123];							inform_L[118][3] = l_cell_wire[124];							inform_L[126][3] = l_cell_wire[125];							inform_L[119][3] = l_cell_wire[126];							inform_L[127][3] = l_cell_wire[127];						end
						5:						begin							inform_R[0][5] = r_cell_wire[0];							inform_R[16][5] = r_cell_wire[1];							inform_R[1][5] = r_cell_wire[2];							inform_R[17][5] = r_cell_wire[3];							inform_R[2][5] = r_cell_wire[4];							inform_R[18][5] = r_cell_wire[5];							inform_R[3][5] = r_cell_wire[6];							inform_R[19][5] = r_cell_wire[7];							inform_R[4][5] = r_cell_wire[8];							inform_R[20][5] = r_cell_wire[9];							inform_R[5][5] = r_cell_wire[10];							inform_R[21][5] = r_cell_wire[11];							inform_R[6][5] = r_cell_wire[12];							inform_R[22][5] = r_cell_wire[13];							inform_R[7][5] = r_cell_wire[14];							inform_R[23][5] = r_cell_wire[15];							inform_R[8][5] = r_cell_wire[16];							inform_R[24][5] = r_cell_wire[17];							inform_R[9][5] = r_cell_wire[18];							inform_R[25][5] = r_cell_wire[19];							inform_R[10][5] = r_cell_wire[20];							inform_R[26][5] = r_cell_wire[21];							inform_R[11][5] = r_cell_wire[22];							inform_R[27][5] = r_cell_wire[23];							inform_R[12][5] = r_cell_wire[24];							inform_R[28][5] = r_cell_wire[25];							inform_R[13][5] = r_cell_wire[26];							inform_R[29][5] = r_cell_wire[27];							inform_R[14][5] = r_cell_wire[28];							inform_R[30][5] = r_cell_wire[29];							inform_R[15][5] = r_cell_wire[30];							inform_R[31][5] = r_cell_wire[31];							inform_R[32][5] = r_cell_wire[32];							inform_R[48][5] = r_cell_wire[33];							inform_R[33][5] = r_cell_wire[34];							inform_R[49][5] = r_cell_wire[35];							inform_R[34][5] = r_cell_wire[36];							inform_R[50][5] = r_cell_wire[37];							inform_R[35][5] = r_cell_wire[38];							inform_R[51][5] = r_cell_wire[39];							inform_R[36][5] = r_cell_wire[40];							inform_R[52][5] = r_cell_wire[41];							inform_R[37][5] = r_cell_wire[42];							inform_R[53][5] = r_cell_wire[43];							inform_R[38][5] = r_cell_wire[44];							inform_R[54][5] = r_cell_wire[45];							inform_R[39][5] = r_cell_wire[46];							inform_R[55][5] = r_cell_wire[47];							inform_R[40][5] = r_cell_wire[48];							inform_R[56][5] = r_cell_wire[49];							inform_R[41][5] = r_cell_wire[50];							inform_R[57][5] = r_cell_wire[51];							inform_R[42][5] = r_cell_wire[52];							inform_R[58][5] = r_cell_wire[53];							inform_R[43][5] = r_cell_wire[54];							inform_R[59][5] = r_cell_wire[55];							inform_R[44][5] = r_cell_wire[56];							inform_R[60][5] = r_cell_wire[57];							inform_R[45][5] = r_cell_wire[58];							inform_R[61][5] = r_cell_wire[59];							inform_R[46][5] = r_cell_wire[60];							inform_R[62][5] = r_cell_wire[61];							inform_R[47][5] = r_cell_wire[62];							inform_R[63][5] = r_cell_wire[63];							inform_R[64][5] = r_cell_wire[64];							inform_R[80][5] = r_cell_wire[65];							inform_R[65][5] = r_cell_wire[66];							inform_R[81][5] = r_cell_wire[67];							inform_R[66][5] = r_cell_wire[68];							inform_R[82][5] = r_cell_wire[69];							inform_R[67][5] = r_cell_wire[70];							inform_R[83][5] = r_cell_wire[71];							inform_R[68][5] = r_cell_wire[72];							inform_R[84][5] = r_cell_wire[73];							inform_R[69][5] = r_cell_wire[74];							inform_R[85][5] = r_cell_wire[75];							inform_R[70][5] = r_cell_wire[76];							inform_R[86][5] = r_cell_wire[77];							inform_R[71][5] = r_cell_wire[78];							inform_R[87][5] = r_cell_wire[79];							inform_R[72][5] = r_cell_wire[80];							inform_R[88][5] = r_cell_wire[81];							inform_R[73][5] = r_cell_wire[82];							inform_R[89][5] = r_cell_wire[83];							inform_R[74][5] = r_cell_wire[84];							inform_R[90][5] = r_cell_wire[85];							inform_R[75][5] = r_cell_wire[86];							inform_R[91][5] = r_cell_wire[87];							inform_R[76][5] = r_cell_wire[88];							inform_R[92][5] = r_cell_wire[89];							inform_R[77][5] = r_cell_wire[90];							inform_R[93][5] = r_cell_wire[91];							inform_R[78][5] = r_cell_wire[92];							inform_R[94][5] = r_cell_wire[93];							inform_R[79][5] = r_cell_wire[94];							inform_R[95][5] = r_cell_wire[95];							inform_R[96][5] = r_cell_wire[96];							inform_R[112][5] = r_cell_wire[97];							inform_R[97][5] = r_cell_wire[98];							inform_R[113][5] = r_cell_wire[99];							inform_R[98][5] = r_cell_wire[100];							inform_R[114][5] = r_cell_wire[101];							inform_R[99][5] = r_cell_wire[102];							inform_R[115][5] = r_cell_wire[103];							inform_R[100][5] = r_cell_wire[104];							inform_R[116][5] = r_cell_wire[105];							inform_R[101][5] = r_cell_wire[106];							inform_R[117][5] = r_cell_wire[107];							inform_R[102][5] = r_cell_wire[108];							inform_R[118][5] = r_cell_wire[109];							inform_R[103][5] = r_cell_wire[110];							inform_R[119][5] = r_cell_wire[111];							inform_R[104][5] = r_cell_wire[112];							inform_R[120][5] = r_cell_wire[113];							inform_R[105][5] = r_cell_wire[114];							inform_R[121][5] = r_cell_wire[115];							inform_R[106][5] = r_cell_wire[116];							inform_R[122][5] = r_cell_wire[117];							inform_R[107][5] = r_cell_wire[118];							inform_R[123][5] = r_cell_wire[119];							inform_R[108][5] = r_cell_wire[120];							inform_R[124][5] = r_cell_wire[121];							inform_R[109][5] = r_cell_wire[122];							inform_R[125][5] = r_cell_wire[123];							inform_R[110][5] = r_cell_wire[124];							inform_R[126][5] = r_cell_wire[125];							inform_R[111][5] = r_cell_wire[126];							inform_R[127][5] = r_cell_wire[127];							inform_L[0][4] = l_cell_wire[0];							inform_L[16][4] = l_cell_wire[1];							inform_L[1][4] = l_cell_wire[2];							inform_L[17][4] = l_cell_wire[3];							inform_L[2][4] = l_cell_wire[4];							inform_L[18][4] = l_cell_wire[5];							inform_L[3][4] = l_cell_wire[6];							inform_L[19][4] = l_cell_wire[7];							inform_L[4][4] = l_cell_wire[8];							inform_L[20][4] = l_cell_wire[9];							inform_L[5][4] = l_cell_wire[10];							inform_L[21][4] = l_cell_wire[11];							inform_L[6][4] = l_cell_wire[12];							inform_L[22][4] = l_cell_wire[13];							inform_L[7][4] = l_cell_wire[14];							inform_L[23][4] = l_cell_wire[15];							inform_L[8][4] = l_cell_wire[16];							inform_L[24][4] = l_cell_wire[17];							inform_L[9][4] = l_cell_wire[18];							inform_L[25][4] = l_cell_wire[19];							inform_L[10][4] = l_cell_wire[20];							inform_L[26][4] = l_cell_wire[21];							inform_L[11][4] = l_cell_wire[22];							inform_L[27][4] = l_cell_wire[23];							inform_L[12][4] = l_cell_wire[24];							inform_L[28][4] = l_cell_wire[25];							inform_L[13][4] = l_cell_wire[26];							inform_L[29][4] = l_cell_wire[27];							inform_L[14][4] = l_cell_wire[28];							inform_L[30][4] = l_cell_wire[29];							inform_L[15][4] = l_cell_wire[30];							inform_L[31][4] = l_cell_wire[31];							inform_L[32][4] = l_cell_wire[32];							inform_L[48][4] = l_cell_wire[33];							inform_L[33][4] = l_cell_wire[34];							inform_L[49][4] = l_cell_wire[35];							inform_L[34][4] = l_cell_wire[36];							inform_L[50][4] = l_cell_wire[37];							inform_L[35][4] = l_cell_wire[38];							inform_L[51][4] = l_cell_wire[39];							inform_L[36][4] = l_cell_wire[40];							inform_L[52][4] = l_cell_wire[41];							inform_L[37][4] = l_cell_wire[42];							inform_L[53][4] = l_cell_wire[43];							inform_L[38][4] = l_cell_wire[44];							inform_L[54][4] = l_cell_wire[45];							inform_L[39][4] = l_cell_wire[46];							inform_L[55][4] = l_cell_wire[47];							inform_L[40][4] = l_cell_wire[48];							inform_L[56][4] = l_cell_wire[49];							inform_L[41][4] = l_cell_wire[50];							inform_L[57][4] = l_cell_wire[51];							inform_L[42][4] = l_cell_wire[52];							inform_L[58][4] = l_cell_wire[53];							inform_L[43][4] = l_cell_wire[54];							inform_L[59][4] = l_cell_wire[55];							inform_L[44][4] = l_cell_wire[56];							inform_L[60][4] = l_cell_wire[57];							inform_L[45][4] = l_cell_wire[58];							inform_L[61][4] = l_cell_wire[59];							inform_L[46][4] = l_cell_wire[60];							inform_L[62][4] = l_cell_wire[61];							inform_L[47][4] = l_cell_wire[62];							inform_L[63][4] = l_cell_wire[63];							inform_L[64][4] = l_cell_wire[64];							inform_L[80][4] = l_cell_wire[65];							inform_L[65][4] = l_cell_wire[66];							inform_L[81][4] = l_cell_wire[67];							inform_L[66][4] = l_cell_wire[68];							inform_L[82][4] = l_cell_wire[69];							inform_L[67][4] = l_cell_wire[70];							inform_L[83][4] = l_cell_wire[71];							inform_L[68][4] = l_cell_wire[72];							inform_L[84][4] = l_cell_wire[73];							inform_L[69][4] = l_cell_wire[74];							inform_L[85][4] = l_cell_wire[75];							inform_L[70][4] = l_cell_wire[76];							inform_L[86][4] = l_cell_wire[77];							inform_L[71][4] = l_cell_wire[78];							inform_L[87][4] = l_cell_wire[79];							inform_L[72][4] = l_cell_wire[80];							inform_L[88][4] = l_cell_wire[81];							inform_L[73][4] = l_cell_wire[82];							inform_L[89][4] = l_cell_wire[83];							inform_L[74][4] = l_cell_wire[84];							inform_L[90][4] = l_cell_wire[85];							inform_L[75][4] = l_cell_wire[86];							inform_L[91][4] = l_cell_wire[87];							inform_L[76][4] = l_cell_wire[88];							inform_L[92][4] = l_cell_wire[89];							inform_L[77][4] = l_cell_wire[90];							inform_L[93][4] = l_cell_wire[91];							inform_L[78][4] = l_cell_wire[92];							inform_L[94][4] = l_cell_wire[93];							inform_L[79][4] = l_cell_wire[94];							inform_L[95][4] = l_cell_wire[95];							inform_L[96][4] = l_cell_wire[96];							inform_L[112][4] = l_cell_wire[97];							inform_L[97][4] = l_cell_wire[98];							inform_L[113][4] = l_cell_wire[99];							inform_L[98][4] = l_cell_wire[100];							inform_L[114][4] = l_cell_wire[101];							inform_L[99][4] = l_cell_wire[102];							inform_L[115][4] = l_cell_wire[103];							inform_L[100][4] = l_cell_wire[104];							inform_L[116][4] = l_cell_wire[105];							inform_L[101][4] = l_cell_wire[106];							inform_L[117][4] = l_cell_wire[107];							inform_L[102][4] = l_cell_wire[108];							inform_L[118][4] = l_cell_wire[109];							inform_L[103][4] = l_cell_wire[110];							inform_L[119][4] = l_cell_wire[111];							inform_L[104][4] = l_cell_wire[112];							inform_L[120][4] = l_cell_wire[113];							inform_L[105][4] = l_cell_wire[114];							inform_L[121][4] = l_cell_wire[115];							inform_L[106][4] = l_cell_wire[116];							inform_L[122][4] = l_cell_wire[117];							inform_L[107][4] = l_cell_wire[118];							inform_L[123][4] = l_cell_wire[119];							inform_L[108][4] = l_cell_wire[120];							inform_L[124][4] = l_cell_wire[121];							inform_L[109][4] = l_cell_wire[122];							inform_L[125][4] = l_cell_wire[123];							inform_L[110][4] = l_cell_wire[124];							inform_L[126][4] = l_cell_wire[125];							inform_L[111][4] = l_cell_wire[126];							inform_L[127][4] = l_cell_wire[127];						end
						6:						begin							inform_R[0][6] = r_cell_wire[0];							inform_R[32][6] = r_cell_wire[1];							inform_R[1][6] = r_cell_wire[2];							inform_R[33][6] = r_cell_wire[3];							inform_R[2][6] = r_cell_wire[4];							inform_R[34][6] = r_cell_wire[5];							inform_R[3][6] = r_cell_wire[6];							inform_R[35][6] = r_cell_wire[7];							inform_R[4][6] = r_cell_wire[8];							inform_R[36][6] = r_cell_wire[9];							inform_R[5][6] = r_cell_wire[10];							inform_R[37][6] = r_cell_wire[11];							inform_R[6][6] = r_cell_wire[12];							inform_R[38][6] = r_cell_wire[13];							inform_R[7][6] = r_cell_wire[14];							inform_R[39][6] = r_cell_wire[15];							inform_R[8][6] = r_cell_wire[16];							inform_R[40][6] = r_cell_wire[17];							inform_R[9][6] = r_cell_wire[18];							inform_R[41][6] = r_cell_wire[19];							inform_R[10][6] = r_cell_wire[20];							inform_R[42][6] = r_cell_wire[21];							inform_R[11][6] = r_cell_wire[22];							inform_R[43][6] = r_cell_wire[23];							inform_R[12][6] = r_cell_wire[24];							inform_R[44][6] = r_cell_wire[25];							inform_R[13][6] = r_cell_wire[26];							inform_R[45][6] = r_cell_wire[27];							inform_R[14][6] = r_cell_wire[28];							inform_R[46][6] = r_cell_wire[29];							inform_R[15][6] = r_cell_wire[30];							inform_R[47][6] = r_cell_wire[31];							inform_R[16][6] = r_cell_wire[32];							inform_R[48][6] = r_cell_wire[33];							inform_R[17][6] = r_cell_wire[34];							inform_R[49][6] = r_cell_wire[35];							inform_R[18][6] = r_cell_wire[36];							inform_R[50][6] = r_cell_wire[37];							inform_R[19][6] = r_cell_wire[38];							inform_R[51][6] = r_cell_wire[39];							inform_R[20][6] = r_cell_wire[40];							inform_R[52][6] = r_cell_wire[41];							inform_R[21][6] = r_cell_wire[42];							inform_R[53][6] = r_cell_wire[43];							inform_R[22][6] = r_cell_wire[44];							inform_R[54][6] = r_cell_wire[45];							inform_R[23][6] = r_cell_wire[46];							inform_R[55][6] = r_cell_wire[47];							inform_R[24][6] = r_cell_wire[48];							inform_R[56][6] = r_cell_wire[49];							inform_R[25][6] = r_cell_wire[50];							inform_R[57][6] = r_cell_wire[51];							inform_R[26][6] = r_cell_wire[52];							inform_R[58][6] = r_cell_wire[53];							inform_R[27][6] = r_cell_wire[54];							inform_R[59][6] = r_cell_wire[55];							inform_R[28][6] = r_cell_wire[56];							inform_R[60][6] = r_cell_wire[57];							inform_R[29][6] = r_cell_wire[58];							inform_R[61][6] = r_cell_wire[59];							inform_R[30][6] = r_cell_wire[60];							inform_R[62][6] = r_cell_wire[61];							inform_R[31][6] = r_cell_wire[62];							inform_R[63][6] = r_cell_wire[63];							inform_R[64][6] = r_cell_wire[64];							inform_R[96][6] = r_cell_wire[65];							inform_R[65][6] = r_cell_wire[66];							inform_R[97][6] = r_cell_wire[67];							inform_R[66][6] = r_cell_wire[68];							inform_R[98][6] = r_cell_wire[69];							inform_R[67][6] = r_cell_wire[70];							inform_R[99][6] = r_cell_wire[71];							inform_R[68][6] = r_cell_wire[72];							inform_R[100][6] = r_cell_wire[73];							inform_R[69][6] = r_cell_wire[74];							inform_R[101][6] = r_cell_wire[75];							inform_R[70][6] = r_cell_wire[76];							inform_R[102][6] = r_cell_wire[77];							inform_R[71][6] = r_cell_wire[78];							inform_R[103][6] = r_cell_wire[79];							inform_R[72][6] = r_cell_wire[80];							inform_R[104][6] = r_cell_wire[81];							inform_R[73][6] = r_cell_wire[82];							inform_R[105][6] = r_cell_wire[83];							inform_R[74][6] = r_cell_wire[84];							inform_R[106][6] = r_cell_wire[85];							inform_R[75][6] = r_cell_wire[86];							inform_R[107][6] = r_cell_wire[87];							inform_R[76][6] = r_cell_wire[88];							inform_R[108][6] = r_cell_wire[89];							inform_R[77][6] = r_cell_wire[90];							inform_R[109][6] = r_cell_wire[91];							inform_R[78][6] = r_cell_wire[92];							inform_R[110][6] = r_cell_wire[93];							inform_R[79][6] = r_cell_wire[94];							inform_R[111][6] = r_cell_wire[95];							inform_R[80][6] = r_cell_wire[96];							inform_R[112][6] = r_cell_wire[97];							inform_R[81][6] = r_cell_wire[98];							inform_R[113][6] = r_cell_wire[99];							inform_R[82][6] = r_cell_wire[100];							inform_R[114][6] = r_cell_wire[101];							inform_R[83][6] = r_cell_wire[102];							inform_R[115][6] = r_cell_wire[103];							inform_R[84][6] = r_cell_wire[104];							inform_R[116][6] = r_cell_wire[105];							inform_R[85][6] = r_cell_wire[106];							inform_R[117][6] = r_cell_wire[107];							inform_R[86][6] = r_cell_wire[108];							inform_R[118][6] = r_cell_wire[109];							inform_R[87][6] = r_cell_wire[110];							inform_R[119][6] = r_cell_wire[111];							inform_R[88][6] = r_cell_wire[112];							inform_R[120][6] = r_cell_wire[113];							inform_R[89][6] = r_cell_wire[114];							inform_R[121][6] = r_cell_wire[115];							inform_R[90][6] = r_cell_wire[116];							inform_R[122][6] = r_cell_wire[117];							inform_R[91][6] = r_cell_wire[118];							inform_R[123][6] = r_cell_wire[119];							inform_R[92][6] = r_cell_wire[120];							inform_R[124][6] = r_cell_wire[121];							inform_R[93][6] = r_cell_wire[122];							inform_R[125][6] = r_cell_wire[123];							inform_R[94][6] = r_cell_wire[124];							inform_R[126][6] = r_cell_wire[125];							inform_R[95][6] = r_cell_wire[126];							inform_R[127][6] = r_cell_wire[127];							inform_L[0][5] = l_cell_wire[0];							inform_L[32][5] = l_cell_wire[1];							inform_L[1][5] = l_cell_wire[2];							inform_L[33][5] = l_cell_wire[3];							inform_L[2][5] = l_cell_wire[4];							inform_L[34][5] = l_cell_wire[5];							inform_L[3][5] = l_cell_wire[6];							inform_L[35][5] = l_cell_wire[7];							inform_L[4][5] = l_cell_wire[8];							inform_L[36][5] = l_cell_wire[9];							inform_L[5][5] = l_cell_wire[10];							inform_L[37][5] = l_cell_wire[11];							inform_L[6][5] = l_cell_wire[12];							inform_L[38][5] = l_cell_wire[13];							inform_L[7][5] = l_cell_wire[14];							inform_L[39][5] = l_cell_wire[15];							inform_L[8][5] = l_cell_wire[16];							inform_L[40][5] = l_cell_wire[17];							inform_L[9][5] = l_cell_wire[18];							inform_L[41][5] = l_cell_wire[19];							inform_L[10][5] = l_cell_wire[20];							inform_L[42][5] = l_cell_wire[21];							inform_L[11][5] = l_cell_wire[22];							inform_L[43][5] = l_cell_wire[23];							inform_L[12][5] = l_cell_wire[24];							inform_L[44][5] = l_cell_wire[25];							inform_L[13][5] = l_cell_wire[26];							inform_L[45][5] = l_cell_wire[27];							inform_L[14][5] = l_cell_wire[28];							inform_L[46][5] = l_cell_wire[29];							inform_L[15][5] = l_cell_wire[30];							inform_L[47][5] = l_cell_wire[31];							inform_L[16][5] = l_cell_wire[32];							inform_L[48][5] = l_cell_wire[33];							inform_L[17][5] = l_cell_wire[34];							inform_L[49][5] = l_cell_wire[35];							inform_L[18][5] = l_cell_wire[36];							inform_L[50][5] = l_cell_wire[37];							inform_L[19][5] = l_cell_wire[38];							inform_L[51][5] = l_cell_wire[39];							inform_L[20][5] = l_cell_wire[40];							inform_L[52][5] = l_cell_wire[41];							inform_L[21][5] = l_cell_wire[42];							inform_L[53][5] = l_cell_wire[43];							inform_L[22][5] = l_cell_wire[44];							inform_L[54][5] = l_cell_wire[45];							inform_L[23][5] = l_cell_wire[46];							inform_L[55][5] = l_cell_wire[47];							inform_L[24][5] = l_cell_wire[48];							inform_L[56][5] = l_cell_wire[49];							inform_L[25][5] = l_cell_wire[50];							inform_L[57][5] = l_cell_wire[51];							inform_L[26][5] = l_cell_wire[52];							inform_L[58][5] = l_cell_wire[53];							inform_L[27][5] = l_cell_wire[54];							inform_L[59][5] = l_cell_wire[55];							inform_L[28][5] = l_cell_wire[56];							inform_L[60][5] = l_cell_wire[57];							inform_L[29][5] = l_cell_wire[58];							inform_L[61][5] = l_cell_wire[59];							inform_L[30][5] = l_cell_wire[60];							inform_L[62][5] = l_cell_wire[61];							inform_L[31][5] = l_cell_wire[62];							inform_L[63][5] = l_cell_wire[63];							inform_L[64][5] = l_cell_wire[64];							inform_L[96][5] = l_cell_wire[65];							inform_L[65][5] = l_cell_wire[66];							inform_L[97][5] = l_cell_wire[67];							inform_L[66][5] = l_cell_wire[68];							inform_L[98][5] = l_cell_wire[69];							inform_L[67][5] = l_cell_wire[70];							inform_L[99][5] = l_cell_wire[71];							inform_L[68][5] = l_cell_wire[72];							inform_L[100][5] = l_cell_wire[73];							inform_L[69][5] = l_cell_wire[74];							inform_L[101][5] = l_cell_wire[75];							inform_L[70][5] = l_cell_wire[76];							inform_L[102][5] = l_cell_wire[77];							inform_L[71][5] = l_cell_wire[78];							inform_L[103][5] = l_cell_wire[79];							inform_L[72][5] = l_cell_wire[80];							inform_L[104][5] = l_cell_wire[81];							inform_L[73][5] = l_cell_wire[82];							inform_L[105][5] = l_cell_wire[83];							inform_L[74][5] = l_cell_wire[84];							inform_L[106][5] = l_cell_wire[85];							inform_L[75][5] = l_cell_wire[86];							inform_L[107][5] = l_cell_wire[87];							inform_L[76][5] = l_cell_wire[88];							inform_L[108][5] = l_cell_wire[89];							inform_L[77][5] = l_cell_wire[90];							inform_L[109][5] = l_cell_wire[91];							inform_L[78][5] = l_cell_wire[92];							inform_L[110][5] = l_cell_wire[93];							inform_L[79][5] = l_cell_wire[94];							inform_L[111][5] = l_cell_wire[95];							inform_L[80][5] = l_cell_wire[96];							inform_L[112][5] = l_cell_wire[97];							inform_L[81][5] = l_cell_wire[98];							inform_L[113][5] = l_cell_wire[99];							inform_L[82][5] = l_cell_wire[100];							inform_L[114][5] = l_cell_wire[101];							inform_L[83][5] = l_cell_wire[102];							inform_L[115][5] = l_cell_wire[103];							inform_L[84][5] = l_cell_wire[104];							inform_L[116][5] = l_cell_wire[105];							inform_L[85][5] = l_cell_wire[106];							inform_L[117][5] = l_cell_wire[107];							inform_L[86][5] = l_cell_wire[108];							inform_L[118][5] = l_cell_wire[109];							inform_L[87][5] = l_cell_wire[110];							inform_L[119][5] = l_cell_wire[111];							inform_L[88][5] = l_cell_wire[112];							inform_L[120][5] = l_cell_wire[113];							inform_L[89][5] = l_cell_wire[114];							inform_L[121][5] = l_cell_wire[115];							inform_L[90][5] = l_cell_wire[116];							inform_L[122][5] = l_cell_wire[117];							inform_L[91][5] = l_cell_wire[118];							inform_L[123][5] = l_cell_wire[119];							inform_L[92][5] = l_cell_wire[120];							inform_L[124][5] = l_cell_wire[121];							inform_L[93][5] = l_cell_wire[122];							inform_L[125][5] = l_cell_wire[123];							inform_L[94][5] = l_cell_wire[124];							inform_L[126][5] = l_cell_wire[125];							inform_L[95][5] = l_cell_wire[126];							inform_L[127][5] = l_cell_wire[127];						end
						7:						begin							inform_R[0][7] = r_cell_wire[0];							inform_R[64][7] = r_cell_wire[1];							inform_R[1][7] = r_cell_wire[2];							inform_R[65][7] = r_cell_wire[3];							inform_R[2][7] = r_cell_wire[4];							inform_R[66][7] = r_cell_wire[5];							inform_R[3][7] = r_cell_wire[6];							inform_R[67][7] = r_cell_wire[7];							inform_R[4][7] = r_cell_wire[8];							inform_R[68][7] = r_cell_wire[9];							inform_R[5][7] = r_cell_wire[10];							inform_R[69][7] = r_cell_wire[11];							inform_R[6][7] = r_cell_wire[12];							inform_R[70][7] = r_cell_wire[13];							inform_R[7][7] = r_cell_wire[14];							inform_R[71][7] = r_cell_wire[15];							inform_R[8][7] = r_cell_wire[16];							inform_R[72][7] = r_cell_wire[17];							inform_R[9][7] = r_cell_wire[18];							inform_R[73][7] = r_cell_wire[19];							inform_R[10][7] = r_cell_wire[20];							inform_R[74][7] = r_cell_wire[21];							inform_R[11][7] = r_cell_wire[22];							inform_R[75][7] = r_cell_wire[23];							inform_R[12][7] = r_cell_wire[24];							inform_R[76][7] = r_cell_wire[25];							inform_R[13][7] = r_cell_wire[26];							inform_R[77][7] = r_cell_wire[27];							inform_R[14][7] = r_cell_wire[28];							inform_R[78][7] = r_cell_wire[29];							inform_R[15][7] = r_cell_wire[30];							inform_R[79][7] = r_cell_wire[31];							inform_R[16][7] = r_cell_wire[32];							inform_R[80][7] = r_cell_wire[33];							inform_R[17][7] = r_cell_wire[34];							inform_R[81][7] = r_cell_wire[35];							inform_R[18][7] = r_cell_wire[36];							inform_R[82][7] = r_cell_wire[37];							inform_R[19][7] = r_cell_wire[38];							inform_R[83][7] = r_cell_wire[39];							inform_R[20][7] = r_cell_wire[40];							inform_R[84][7] = r_cell_wire[41];							inform_R[21][7] = r_cell_wire[42];							inform_R[85][7] = r_cell_wire[43];							inform_R[22][7] = r_cell_wire[44];							inform_R[86][7] = r_cell_wire[45];							inform_R[23][7] = r_cell_wire[46];							inform_R[87][7] = r_cell_wire[47];							inform_R[24][7] = r_cell_wire[48];							inform_R[88][7] = r_cell_wire[49];							inform_R[25][7] = r_cell_wire[50];							inform_R[89][7] = r_cell_wire[51];							inform_R[26][7] = r_cell_wire[52];							inform_R[90][7] = r_cell_wire[53];							inform_R[27][7] = r_cell_wire[54];							inform_R[91][7] = r_cell_wire[55];							inform_R[28][7] = r_cell_wire[56];							inform_R[92][7] = r_cell_wire[57];							inform_R[29][7] = r_cell_wire[58];							inform_R[93][7] = r_cell_wire[59];							inform_R[30][7] = r_cell_wire[60];							inform_R[94][7] = r_cell_wire[61];							inform_R[31][7] = r_cell_wire[62];							inform_R[95][7] = r_cell_wire[63];							inform_R[32][7] = r_cell_wire[64];							inform_R[96][7] = r_cell_wire[65];							inform_R[33][7] = r_cell_wire[66];							inform_R[97][7] = r_cell_wire[67];							inform_R[34][7] = r_cell_wire[68];							inform_R[98][7] = r_cell_wire[69];							inform_R[35][7] = r_cell_wire[70];							inform_R[99][7] = r_cell_wire[71];							inform_R[36][7] = r_cell_wire[72];							inform_R[100][7] = r_cell_wire[73];							inform_R[37][7] = r_cell_wire[74];							inform_R[101][7] = r_cell_wire[75];							inform_R[38][7] = r_cell_wire[76];							inform_R[102][7] = r_cell_wire[77];							inform_R[39][7] = r_cell_wire[78];							inform_R[103][7] = r_cell_wire[79];							inform_R[40][7] = r_cell_wire[80];							inform_R[104][7] = r_cell_wire[81];							inform_R[41][7] = r_cell_wire[82];							inform_R[105][7] = r_cell_wire[83];							inform_R[42][7] = r_cell_wire[84];							inform_R[106][7] = r_cell_wire[85];							inform_R[43][7] = r_cell_wire[86];							inform_R[107][7] = r_cell_wire[87];							inform_R[44][7] = r_cell_wire[88];							inform_R[108][7] = r_cell_wire[89];							inform_R[45][7] = r_cell_wire[90];							inform_R[109][7] = r_cell_wire[91];							inform_R[46][7] = r_cell_wire[92];							inform_R[110][7] = r_cell_wire[93];							inform_R[47][7] = r_cell_wire[94];							inform_R[111][7] = r_cell_wire[95];							inform_R[48][7] = r_cell_wire[96];							inform_R[112][7] = r_cell_wire[97];							inform_R[49][7] = r_cell_wire[98];							inform_R[113][7] = r_cell_wire[99];							inform_R[50][7] = r_cell_wire[100];							inform_R[114][7] = r_cell_wire[101];							inform_R[51][7] = r_cell_wire[102];							inform_R[115][7] = r_cell_wire[103];							inform_R[52][7] = r_cell_wire[104];							inform_R[116][7] = r_cell_wire[105];							inform_R[53][7] = r_cell_wire[106];							inform_R[117][7] = r_cell_wire[107];							inform_R[54][7] = r_cell_wire[108];							inform_R[118][7] = r_cell_wire[109];							inform_R[55][7] = r_cell_wire[110];							inform_R[119][7] = r_cell_wire[111];							inform_R[56][7] = r_cell_wire[112];							inform_R[120][7] = r_cell_wire[113];							inform_R[57][7] = r_cell_wire[114];							inform_R[121][7] = r_cell_wire[115];							inform_R[58][7] = r_cell_wire[116];							inform_R[122][7] = r_cell_wire[117];							inform_R[59][7] = r_cell_wire[118];							inform_R[123][7] = r_cell_wire[119];							inform_R[60][7] = r_cell_wire[120];							inform_R[124][7] = r_cell_wire[121];							inform_R[61][7] = r_cell_wire[122];							inform_R[125][7] = r_cell_wire[123];							inform_R[62][7] = r_cell_wire[124];							inform_R[126][7] = r_cell_wire[125];							inform_R[63][7] = r_cell_wire[126];							inform_R[127][7] = r_cell_wire[127];							inform_L[0][6] = l_cell_wire[0];							inform_L[64][6] = l_cell_wire[1];							inform_L[1][6] = l_cell_wire[2];							inform_L[65][6] = l_cell_wire[3];							inform_L[2][6] = l_cell_wire[4];							inform_L[66][6] = l_cell_wire[5];							inform_L[3][6] = l_cell_wire[6];							inform_L[67][6] = l_cell_wire[7];							inform_L[4][6] = l_cell_wire[8];							inform_L[68][6] = l_cell_wire[9];							inform_L[5][6] = l_cell_wire[10];							inform_L[69][6] = l_cell_wire[11];							inform_L[6][6] = l_cell_wire[12];							inform_L[70][6] = l_cell_wire[13];							inform_L[7][6] = l_cell_wire[14];							inform_L[71][6] = l_cell_wire[15];							inform_L[8][6] = l_cell_wire[16];							inform_L[72][6] = l_cell_wire[17];							inform_L[9][6] = l_cell_wire[18];							inform_L[73][6] = l_cell_wire[19];							inform_L[10][6] = l_cell_wire[20];							inform_L[74][6] = l_cell_wire[21];							inform_L[11][6] = l_cell_wire[22];							inform_L[75][6] = l_cell_wire[23];							inform_L[12][6] = l_cell_wire[24];							inform_L[76][6] = l_cell_wire[25];							inform_L[13][6] = l_cell_wire[26];							inform_L[77][6] = l_cell_wire[27];							inform_L[14][6] = l_cell_wire[28];							inform_L[78][6] = l_cell_wire[29];							inform_L[15][6] = l_cell_wire[30];							inform_L[79][6] = l_cell_wire[31];							inform_L[16][6] = l_cell_wire[32];							inform_L[80][6] = l_cell_wire[33];							inform_L[17][6] = l_cell_wire[34];							inform_L[81][6] = l_cell_wire[35];							inform_L[18][6] = l_cell_wire[36];							inform_L[82][6] = l_cell_wire[37];							inform_L[19][6] = l_cell_wire[38];							inform_L[83][6] = l_cell_wire[39];							inform_L[20][6] = l_cell_wire[40];							inform_L[84][6] = l_cell_wire[41];							inform_L[21][6] = l_cell_wire[42];							inform_L[85][6] = l_cell_wire[43];							inform_L[22][6] = l_cell_wire[44];							inform_L[86][6] = l_cell_wire[45];							inform_L[23][6] = l_cell_wire[46];							inform_L[87][6] = l_cell_wire[47];							inform_L[24][6] = l_cell_wire[48];							inform_L[88][6] = l_cell_wire[49];							inform_L[25][6] = l_cell_wire[50];							inform_L[89][6] = l_cell_wire[51];							inform_L[26][6] = l_cell_wire[52];							inform_L[90][6] = l_cell_wire[53];							inform_L[27][6] = l_cell_wire[54];							inform_L[91][6] = l_cell_wire[55];							inform_L[28][6] = l_cell_wire[56];							inform_L[92][6] = l_cell_wire[57];							inform_L[29][6] = l_cell_wire[58];							inform_L[93][6] = l_cell_wire[59];							inform_L[30][6] = l_cell_wire[60];							inform_L[94][6] = l_cell_wire[61];							inform_L[31][6] = l_cell_wire[62];							inform_L[95][6] = l_cell_wire[63];							inform_L[32][6] = l_cell_wire[64];							inform_L[96][6] = l_cell_wire[65];							inform_L[33][6] = l_cell_wire[66];							inform_L[97][6] = l_cell_wire[67];							inform_L[34][6] = l_cell_wire[68];							inform_L[98][6] = l_cell_wire[69];							inform_L[35][6] = l_cell_wire[70];							inform_L[99][6] = l_cell_wire[71];							inform_L[36][6] = l_cell_wire[72];							inform_L[100][6] = l_cell_wire[73];							inform_L[37][6] = l_cell_wire[74];							inform_L[101][6] = l_cell_wire[75];							inform_L[38][6] = l_cell_wire[76];							inform_L[102][6] = l_cell_wire[77];							inform_L[39][6] = l_cell_wire[78];							inform_L[103][6] = l_cell_wire[79];							inform_L[40][6] = l_cell_wire[80];							inform_L[104][6] = l_cell_wire[81];							inform_L[41][6] = l_cell_wire[82];							inform_L[105][6] = l_cell_wire[83];							inform_L[42][6] = l_cell_wire[84];							inform_L[106][6] = l_cell_wire[85];							inform_L[43][6] = l_cell_wire[86];							inform_L[107][6] = l_cell_wire[87];							inform_L[44][6] = l_cell_wire[88];							inform_L[108][6] = l_cell_wire[89];							inform_L[45][6] = l_cell_wire[90];							inform_L[109][6] = l_cell_wire[91];							inform_L[46][6] = l_cell_wire[92];							inform_L[110][6] = l_cell_wire[93];							inform_L[47][6] = l_cell_wire[94];							inform_L[111][6] = l_cell_wire[95];							inform_L[48][6] = l_cell_wire[96];							inform_L[112][6] = l_cell_wire[97];							inform_L[49][6] = l_cell_wire[98];							inform_L[113][6] = l_cell_wire[99];							inform_L[50][6] = l_cell_wire[100];							inform_L[114][6] = l_cell_wire[101];							inform_L[51][6] = l_cell_wire[102];							inform_L[115][6] = l_cell_wire[103];							inform_L[52][6] = l_cell_wire[104];							inform_L[116][6] = l_cell_wire[105];							inform_L[53][6] = l_cell_wire[106];							inform_L[117][6] = l_cell_wire[107];							inform_L[54][6] = l_cell_wire[108];							inform_L[118][6] = l_cell_wire[109];							inform_L[55][6] = l_cell_wire[110];							inform_L[119][6] = l_cell_wire[111];							inform_L[56][6] = l_cell_wire[112];							inform_L[120][6] = l_cell_wire[113];							inform_L[57][6] = l_cell_wire[114];							inform_L[121][6] = l_cell_wire[115];							inform_L[58][6] = l_cell_wire[116];							inform_L[122][6] = l_cell_wire[117];							inform_L[59][6] = l_cell_wire[118];							inform_L[123][6] = l_cell_wire[119];							inform_L[60][6] = l_cell_wire[120];							inform_L[124][6] = l_cell_wire[121];							inform_L[61][6] = l_cell_wire[122];							inform_L[125][6] = l_cell_wire[123];							inform_L[62][6] = l_cell_wire[124];							inform_L[126][6] = l_cell_wire[125];							inform_L[63][6] = l_cell_wire[126];							inform_L[127][6] = l_cell_wire[127];						end
						default:							for (x = 0; x < 128; x = x + 1)								for (y = 0; y < 7; y = y + 1)								begin									inform_R[x][y+1] <= 8'd0;									inform_L[x][y] <= 8'd0;								end					endcase				end			end
				default:				begin				if (start) begin					inform_R [0][0] <= 8'b0111_1111;					inform_R [1][0] <= 8'b0111_1111;					inform_R [2][0] <= 8'b0111_1111;					inform_R [3][0] <= 8'b0111_1111;					inform_R [4][0] <= 8'b0111_1111;					inform_R [5][0] <= 8'b0111_1111;					inform_R [6][0] <= 8'b0111_1111;					inform_R [7][0] <= 8'b0111_1111;					inform_R [8][0] <= 8'b0111_1111;					inform_R [9][0] <= 8'b0111_1111;					inform_R [10][0] <= 8'b0111_1111;					inform_R [11][0] <= 8'b0111_1111;					inform_R [12][0] <= 8'b0111_1111;					inform_R [13][0] <= 8'b0111_1111;					inform_R [14][0] <= 8'b0111_1111;					inform_R [15][0] <= 8'b0111_1111;					inform_R [16][0] <= 8'b0111_1111;					inform_R [17][0] <= 8'b0111_1111;					inform_R [18][0] <= 8'b0111_1111;					inform_R [19][0] <= 8'b0111_1111;					inform_R [20][0] <= 8'b0111_1111;					inform_R [21][0] <= 8'b0111_1111;					inform_R [22][0] <= 8'b0111_1111;					inform_R [23][0] <= 8'b0111_1111;					inform_R [24][0] <= 8'b0111_1111;					inform_R [25][0] <= 8'b0111_1111;					inform_R [26][0] <= 8'b0111_1111;					inform_R [27][0] <= 8'b0111_1111;					inform_R [28][0] <= 8'b0111_1111;					inform_R [29][0] <= 8'b0111_1111;					inform_R [30][0] <= 8'b0111_1111;					inform_R [31][0] <= 8'b0000_0000;					inform_R [32][0] <= 8'b0111_1111;					inform_R [33][0] <= 8'b0111_1111;					inform_R [34][0] <= 8'b0111_1111;					inform_R [35][0] <= 8'b0111_1111;					inform_R [36][0] <= 8'b0111_1111;					inform_R [37][0] <= 8'b0111_1111;					inform_R [38][0] <= 8'b0111_1111;					inform_R [39][0] <= 8'b0111_1111;					inform_R [40][0] <= 8'b0111_1111;					inform_R [41][0] <= 8'b0111_1111;					inform_R [42][0] <= 8'b0111_1111;					inform_R [43][0] <= 8'b0111_1111;					inform_R [44][0] <= 8'b0111_1111;					inform_R [45][0] <= 8'b0000_0000;					inform_R [46][0] <= 8'b0000_0000;					inform_R [47][0] <= 8'b0000_0000;					inform_R [48][0] <= 8'b0111_1111;					inform_R [49][0] <= 8'b0111_1111;					inform_R [50][0] <= 8'b0111_1111;					inform_R [51][0] <= 8'b0000_0000;					inform_R [52][0] <= 8'b0111_1111;					inform_R [53][0] <= 8'b0000_0000;					inform_R [54][0] <= 8'b0000_0000;					inform_R [55][0] <= 8'b0000_0000;					inform_R [56][0] <= 8'b0111_1111;					inform_R [57][0] <= 8'b0000_0000;					inform_R [58][0] <= 8'b0000_0000;					inform_R [59][0] <= 8'b0000_0000;					inform_R [60][0] <= 8'b0000_0000;					inform_R [61][0] <= 8'b0000_0000;					inform_R [62][0] <= 8'b0000_0000;					inform_R [63][0] <= 8'b0000_0000;					inform_R [64][0] <= 8'b0111_1111;					inform_R [65][0] <= 8'b0111_1111;					inform_R [66][0] <= 8'b0111_1111;					inform_R [67][0] <= 8'b0111_1111;					inform_R [68][0] <= 8'b0111_1111;					inform_R [69][0] <= 8'b0111_1111;					inform_R [70][0] <= 8'b0111_1111;					inform_R [71][0] <= 8'b0000_0000;					inform_R [72][0] <= 8'b0111_1111;					inform_R [73][0] <= 8'b0111_1111;					inform_R [74][0] <= 8'b0111_1111;					inform_R [75][0] <= 8'b0000_0000;					inform_R [76][0] <= 8'b0111_1111;					inform_R [77][0] <= 8'b0000_0000;					inform_R [78][0] <= 8'b0000_0000;					inform_R [79][0] <= 8'b0000_0000;					inform_R [80][0] <= 8'b0111_1111;					inform_R [81][0] <= 8'b0111_1111;					inform_R [82][0] <= 8'b0111_1111;					inform_R [83][0] <= 8'b0000_0000;					inform_R [84][0] <= 8'b0000_0000;					inform_R [85][0] <= 8'b0000_0000;					inform_R [86][0] <= 8'b0000_0000;					inform_R [87][0] <= 8'b0000_0000;					inform_R [88][0] <= 8'b0000_0000;					inform_R [89][0] <= 8'b0000_0000;					inform_R [90][0] <= 8'b0000_0000;					inform_R [91][0] <= 8'b0000_0000;					inform_R [92][0] <= 8'b0000_0000;					inform_R [93][0] <= 8'b0000_0000;					inform_R [94][0] <= 8'b0000_0000;					inform_R [95][0] <= 8'b0000_0000;					inform_R [96][0] <= 8'b0111_1111;					inform_R [97][0] <= 8'b0000_0000;					inform_R [98][0] <= 8'b0000_0000;					inform_R [99][0] <= 8'b0000_0000;					inform_R [100][0] <= 8'b0000_0000;					inform_R [101][0] <= 8'b0000_0000;					inform_R [102][0] <= 8'b0000_0000;					inform_R [103][0] <= 8'b0000_0000;					inform_R [104][0] <= 8'b0000_0000;					inform_R [105][0] <= 8'b0000_0000;					inform_R [106][0] <= 8'b0000_0000;					inform_R [107][0] <= 8'b0000_0000;					inform_R [108][0] <= 8'b0000_0000;					inform_R [109][0] <= 8'b0000_0000;					inform_R [110][0] <= 8'b0000_0000;					inform_R [111][0] <= 8'b0000_0000;					inform_R [112][0] <= 8'b0000_0000;					inform_R [113][0] <= 8'b0000_0000;					inform_R [114][0] <= 8'b0000_0000;					inform_R [115][0] <= 8'b0000_0000;					inform_R [116][0] <= 8'b0000_0000;					inform_R [117][0] <= 8'b0000_0000;					inform_R [118][0] <= 8'b0000_0000;					inform_R [119][0] <= 8'b0000_0000;					inform_R [120][0] <= 8'b0000_0000;					inform_R [121][0] <= 8'b0000_0000;					inform_R [122][0] <= 8'b0000_0000;					inform_R [123][0] <= 8'b0000_0000;					inform_R [124][0] <= 8'b0000_0000;					inform_R [125][0] <= 8'b0000_0000;					inform_R [126][0] <= 8'b0000_0000;					inform_R [127][0] <= 8'b0000_0000;					inform_L [0][7] <= LLR_1;					inform_L [1][7] <= LLR_2;					inform_L [2][7] <= LLR_3;					inform_L [3][7] <= LLR_4;					inform_L [4][7] <= LLR_5;					inform_L [5][7] <= LLR_6;					inform_L [6][7] <= LLR_7;					inform_L [7][7] <= LLR_8;					inform_L [8][7] <= LLR_9;					inform_L [9][7] <= LLR_10;					inform_L [10][7] <= LLR_11;					inform_L [11][7] <= LLR_12;					inform_L [12][7] <= LLR_13;					inform_L [13][7] <= LLR_14;					inform_L [14][7] <= LLR_15;					inform_L [15][7] <= LLR_16;					inform_L [16][7] <= LLR_17;					inform_L [17][7] <= LLR_18;					inform_L [18][7] <= LLR_19;					inform_L [19][7] <= LLR_20;					inform_L [20][7] <= LLR_21;					inform_L [21][7] <= LLR_22;					inform_L [22][7] <= LLR_23;					inform_L [23][7] <= LLR_24;					inform_L [24][7] <= LLR_25;					inform_L [25][7] <= LLR_26;					inform_L [26][7] <= LLR_27;					inform_L [27][7] <= LLR_28;					inform_L [28][7] <= LLR_29;					inform_L [29][7] <= LLR_30;					inform_L [30][7] <= LLR_31;					inform_L [31][7] <= LLR_32;					inform_L [32][7] <= LLR_33;					inform_L [33][7] <= LLR_34;					inform_L [34][7] <= LLR_35;					inform_L [35][7] <= LLR_36;					inform_L [36][7] <= LLR_37;					inform_L [37][7] <= LLR_38;					inform_L [38][7] <= LLR_39;					inform_L [39][7] <= LLR_40;					inform_L [40][7] <= LLR_41;					inform_L [41][7] <= LLR_42;					inform_L [42][7] <= LLR_43;					inform_L [43][7] <= LLR_44;					inform_L [44][7] <= LLR_45;					inform_L [45][7] <= LLR_46;					inform_L [46][7] <= LLR_47;					inform_L [47][7] <= LLR_48;					inform_L [48][7] <= LLR_49;					inform_L [49][7] <= LLR_50;					inform_L [50][7] <= LLR_51;					inform_L [51][7] <= LLR_52;					inform_L [52][7] <= LLR_53;					inform_L [53][7] <= LLR_54;					inform_L [54][7] <= LLR_55;					inform_L [55][7] <= LLR_56;					inform_L [56][7] <= LLR_57;					inform_L [57][7] <= LLR_58;					inform_L [58][7] <= LLR_59;					inform_L [59][7] <= LLR_60;					inform_L [60][7] <= LLR_61;					inform_L [61][7] <= LLR_62;					inform_L [62][7] <= LLR_63;					inform_L [63][7] <= LLR_64;					inform_L [64][7] <= LLR_65;					inform_L [65][7] <= LLR_66;					inform_L [66][7] <= LLR_67;					inform_L [67][7] <= LLR_68;					inform_L [68][7] <= LLR_69;					inform_L [69][7] <= LLR_70;					inform_L [70][7] <= LLR_71;					inform_L [71][7] <= LLR_72;					inform_L [72][7] <= LLR_73;					inform_L [73][7] <= LLR_74;					inform_L [74][7] <= LLR_75;					inform_L [75][7] <= LLR_76;					inform_L [76][7] <= LLR_77;					inform_L [77][7] <= LLR_78;					inform_L [78][7] <= LLR_79;					inform_L [79][7] <= LLR_80;					inform_L [80][7] <= LLR_81;					inform_L [81][7] <= LLR_82;					inform_L [82][7] <= LLR_83;					inform_L [83][7] <= LLR_84;					inform_L [84][7] <= LLR_85;					inform_L [85][7] <= LLR_86;					inform_L [86][7] <= LLR_87;					inform_L [87][7] <= LLR_88;					inform_L [88][7] <= LLR_89;					inform_L [89][7] <= LLR_90;					inform_L [90][7] <= LLR_91;					inform_L [91][7] <= LLR_92;					inform_L [92][7] <= LLR_93;					inform_L [93][7] <= LLR_94;					inform_L [94][7] <= LLR_95;					inform_L [95][7] <= LLR_96;					inform_L [96][7] <= LLR_97;					inform_L [97][7] <= LLR_98;					inform_L [98][7] <= LLR_99;					inform_L [99][7] <= LLR_100;					inform_L [100][7] <= LLR_101;					inform_L [101][7] <= LLR_102;					inform_L [102][7] <= LLR_103;					inform_L [103][7] <= LLR_104;					inform_L [104][7] <= LLR_105;					inform_L [105][7] <= LLR_106;					inform_L [106][7] <= LLR_107;					inform_L [107][7] <= LLR_108;					inform_L [108][7] <= LLR_109;					inform_L [109][7] <= LLR_110;					inform_L [110][7] <= LLR_111;					inform_L [111][7] <= LLR_112;					inform_L [112][7] <= LLR_113;					inform_L [113][7] <= LLR_114;					inform_L [114][7] <= LLR_115;					inform_L [115][7] <= LLR_116;					inform_L [116][7] <= LLR_117;					inform_L [117][7] <= LLR_118;					inform_L [118][7] <= LLR_119;					inform_L [119][7] <= LLR_120;					inform_L [120][7] <= LLR_121;					inform_L [121][7] <= LLR_122;					inform_L [122][7] <= LLR_123;					inform_L [123][7] <= LLR_124;					inform_L [124][7] <= LLR_125;					inform_L [125][7] <= LLR_126;					inform_L [126][7] <= LLR_127;					inform_L [127][7] <= LLR_128;				end				for (x = 0; x < 128; x = x + 1)					for (y = 0; y < 7; y = y + 1)					begin						inform_R[x][y+1] <= 8'd0;						inform_L[x][y] <= 8'd0;					end			end
		endcase	end
	assign bp_over_flag = (itera_time == `iteration_times + 1) ? 1 : 0;
	always @(*)	begin		case (w2r)			1:			begin				r_cell_reg[0] = inform_R[0][0];				r_cell_reg[1] = inform_R[1][0];				r_cell_reg[2] = inform_R[2][0];				r_cell_reg[3] = inform_R[3][0];				r_cell_reg[4] = inform_R[4][0];				r_cell_reg[5] = inform_R[5][0];				r_cell_reg[6] = inform_R[6][0];				r_cell_reg[7] = inform_R[7][0];				r_cell_reg[8] = inform_R[8][0];				r_cell_reg[9] = inform_R[9][0];				r_cell_reg[10] = inform_R[10][0];				r_cell_reg[11] = inform_R[11][0];				r_cell_reg[12] = inform_R[12][0];				r_cell_reg[13] = inform_R[13][0];				r_cell_reg[14] = inform_R[14][0];				r_cell_reg[15] = inform_R[15][0];				r_cell_reg[16] = inform_R[16][0];				r_cell_reg[17] = inform_R[17][0];				r_cell_reg[18] = inform_R[18][0];				r_cell_reg[19] = inform_R[19][0];				r_cell_reg[20] = inform_R[20][0];				r_cell_reg[21] = inform_R[21][0];				r_cell_reg[22] = inform_R[22][0];				r_cell_reg[23] = inform_R[23][0];				r_cell_reg[24] = inform_R[24][0];				r_cell_reg[25] = inform_R[25][0];				r_cell_reg[26] = inform_R[26][0];				r_cell_reg[27] = inform_R[27][0];				r_cell_reg[28] = inform_R[28][0];				r_cell_reg[29] = inform_R[29][0];				r_cell_reg[30] = inform_R[30][0];				r_cell_reg[31] = inform_R[31][0];				r_cell_reg[32] = inform_R[32][0];				r_cell_reg[33] = inform_R[33][0];				r_cell_reg[34] = inform_R[34][0];				r_cell_reg[35] = inform_R[35][0];				r_cell_reg[36] = inform_R[36][0];				r_cell_reg[37] = inform_R[37][0];				r_cell_reg[38] = inform_R[38][0];				r_cell_reg[39] = inform_R[39][0];				r_cell_reg[40] = inform_R[40][0];				r_cell_reg[41] = inform_R[41][0];				r_cell_reg[42] = inform_R[42][0];				r_cell_reg[43] = inform_R[43][0];				r_cell_reg[44] = inform_R[44][0];				r_cell_reg[45] = inform_R[45][0];				r_cell_reg[46] = inform_R[46][0];				r_cell_reg[47] = inform_R[47][0];				r_cell_reg[48] = inform_R[48][0];				r_cell_reg[49] = inform_R[49][0];				r_cell_reg[50] = inform_R[50][0];				r_cell_reg[51] = inform_R[51][0];				r_cell_reg[52] = inform_R[52][0];				r_cell_reg[53] = inform_R[53][0];				r_cell_reg[54] = inform_R[54][0];				r_cell_reg[55] = inform_R[55][0];				r_cell_reg[56] = inform_R[56][0];				r_cell_reg[57] = inform_R[57][0];				r_cell_reg[58] = inform_R[58][0];				r_cell_reg[59] = inform_R[59][0];				r_cell_reg[60] = inform_R[60][0];				r_cell_reg[61] = inform_R[61][0];				r_cell_reg[62] = inform_R[62][0];				r_cell_reg[63] = inform_R[63][0];				r_cell_reg[64] = inform_R[64][0];				r_cell_reg[65] = inform_R[65][0];				r_cell_reg[66] = inform_R[66][0];				r_cell_reg[67] = inform_R[67][0];				r_cell_reg[68] = inform_R[68][0];				r_cell_reg[69] = inform_R[69][0];				r_cell_reg[70] = inform_R[70][0];				r_cell_reg[71] = inform_R[71][0];				r_cell_reg[72] = inform_R[72][0];				r_cell_reg[73] = inform_R[73][0];				r_cell_reg[74] = inform_R[74][0];				r_cell_reg[75] = inform_R[75][0];				r_cell_reg[76] = inform_R[76][0];				r_cell_reg[77] = inform_R[77][0];				r_cell_reg[78] = inform_R[78][0];				r_cell_reg[79] = inform_R[79][0];				r_cell_reg[80] = inform_R[80][0];				r_cell_reg[81] = inform_R[81][0];				r_cell_reg[82] = inform_R[82][0];				r_cell_reg[83] = inform_R[83][0];				r_cell_reg[84] = inform_R[84][0];				r_cell_reg[85] = inform_R[85][0];				r_cell_reg[86] = inform_R[86][0];				r_cell_reg[87] = inform_R[87][0];				r_cell_reg[88] = inform_R[88][0];				r_cell_reg[89] = inform_R[89][0];				r_cell_reg[90] = inform_R[90][0];				r_cell_reg[91] = inform_R[91][0];				r_cell_reg[92] = inform_R[92][0];				r_cell_reg[93] = inform_R[93][0];				r_cell_reg[94] = inform_R[94][0];				r_cell_reg[95] = inform_R[95][0];				r_cell_reg[96] = inform_R[96][0];				r_cell_reg[97] = inform_R[97][0];				r_cell_reg[98] = inform_R[98][0];				r_cell_reg[99] = inform_R[99][0];				r_cell_reg[100] = inform_R[100][0];				r_cell_reg[101] = inform_R[101][0];				r_cell_reg[102] = inform_R[102][0];				r_cell_reg[103] = inform_R[103][0];				r_cell_reg[104] = inform_R[104][0];				r_cell_reg[105] = inform_R[105][0];				r_cell_reg[106] = inform_R[106][0];				r_cell_reg[107] = inform_R[107][0];				r_cell_reg[108] = inform_R[108][0];				r_cell_reg[109] = inform_R[109][0];				r_cell_reg[110] = inform_R[110][0];				r_cell_reg[111] = inform_R[111][0];				r_cell_reg[112] = inform_R[112][0];				r_cell_reg[113] = inform_R[113][0];				r_cell_reg[114] = inform_R[114][0];				r_cell_reg[115] = inform_R[115][0];				r_cell_reg[116] = inform_R[116][0];				r_cell_reg[117] = inform_R[117][0];				r_cell_reg[118] = inform_R[118][0];				r_cell_reg[119] = inform_R[119][0];				r_cell_reg[120] = inform_R[120][0];				r_cell_reg[121] = inform_R[121][0];				r_cell_reg[122] = inform_R[122][0];				r_cell_reg[123] = inform_R[123][0];				r_cell_reg[124] = inform_R[124][0];				r_cell_reg[125] = inform_R[125][0];				r_cell_reg[126] = inform_R[126][0];				r_cell_reg[127] = inform_R[127][0];				l_cell_reg[0] = inform_L[0][1];				l_cell_reg[1] = inform_L[1][1];				l_cell_reg[2] = inform_L[2][1];				l_cell_reg[3] = inform_L[3][1];				l_cell_reg[4] = inform_L[4][1];				l_cell_reg[5] = inform_L[5][1];				l_cell_reg[6] = inform_L[6][1];				l_cell_reg[7] = inform_L[7][1];				l_cell_reg[8] = inform_L[8][1];				l_cell_reg[9] = inform_L[9][1];				l_cell_reg[10] = inform_L[10][1];				l_cell_reg[11] = inform_L[11][1];				l_cell_reg[12] = inform_L[12][1];				l_cell_reg[13] = inform_L[13][1];				l_cell_reg[14] = inform_L[14][1];				l_cell_reg[15] = inform_L[15][1];				l_cell_reg[16] = inform_L[16][1];				l_cell_reg[17] = inform_L[17][1];				l_cell_reg[18] = inform_L[18][1];				l_cell_reg[19] = inform_L[19][1];				l_cell_reg[20] = inform_L[20][1];				l_cell_reg[21] = inform_L[21][1];				l_cell_reg[22] = inform_L[22][1];				l_cell_reg[23] = inform_L[23][1];				l_cell_reg[24] = inform_L[24][1];				l_cell_reg[25] = inform_L[25][1];				l_cell_reg[26] = inform_L[26][1];				l_cell_reg[27] = inform_L[27][1];				l_cell_reg[28] = inform_L[28][1];				l_cell_reg[29] = inform_L[29][1];				l_cell_reg[30] = inform_L[30][1];				l_cell_reg[31] = inform_L[31][1];				l_cell_reg[32] = inform_L[32][1];				l_cell_reg[33] = inform_L[33][1];				l_cell_reg[34] = inform_L[34][1];				l_cell_reg[35] = inform_L[35][1];				l_cell_reg[36] = inform_L[36][1];				l_cell_reg[37] = inform_L[37][1];				l_cell_reg[38] = inform_L[38][1];				l_cell_reg[39] = inform_L[39][1];				l_cell_reg[40] = inform_L[40][1];				l_cell_reg[41] = inform_L[41][1];				l_cell_reg[42] = inform_L[42][1];				l_cell_reg[43] = inform_L[43][1];				l_cell_reg[44] = inform_L[44][1];				l_cell_reg[45] = inform_L[45][1];				l_cell_reg[46] = inform_L[46][1];				l_cell_reg[47] = inform_L[47][1];				l_cell_reg[48] = inform_L[48][1];				l_cell_reg[49] = inform_L[49][1];				l_cell_reg[50] = inform_L[50][1];				l_cell_reg[51] = inform_L[51][1];				l_cell_reg[52] = inform_L[52][1];				l_cell_reg[53] = inform_L[53][1];				l_cell_reg[54] = inform_L[54][1];				l_cell_reg[55] = inform_L[55][1];				l_cell_reg[56] = inform_L[56][1];				l_cell_reg[57] = inform_L[57][1];				l_cell_reg[58] = inform_L[58][1];				l_cell_reg[59] = inform_L[59][1];				l_cell_reg[60] = inform_L[60][1];				l_cell_reg[61] = inform_L[61][1];				l_cell_reg[62] = inform_L[62][1];				l_cell_reg[63] = inform_L[63][1];				l_cell_reg[64] = inform_L[64][1];				l_cell_reg[65] = inform_L[65][1];				l_cell_reg[66] = inform_L[66][1];				l_cell_reg[67] = inform_L[67][1];				l_cell_reg[68] = inform_L[68][1];				l_cell_reg[69] = inform_L[69][1];				l_cell_reg[70] = inform_L[70][1];				l_cell_reg[71] = inform_L[71][1];				l_cell_reg[72] = inform_L[72][1];				l_cell_reg[73] = inform_L[73][1];				l_cell_reg[74] = inform_L[74][1];				l_cell_reg[75] = inform_L[75][1];				l_cell_reg[76] = inform_L[76][1];				l_cell_reg[77] = inform_L[77][1];				l_cell_reg[78] = inform_L[78][1];				l_cell_reg[79] = inform_L[79][1];				l_cell_reg[80] = inform_L[80][1];				l_cell_reg[81] = inform_L[81][1];				l_cell_reg[82] = inform_L[82][1];				l_cell_reg[83] = inform_L[83][1];				l_cell_reg[84] = inform_L[84][1];				l_cell_reg[85] = inform_L[85][1];				l_cell_reg[86] = inform_L[86][1];				l_cell_reg[87] = inform_L[87][1];				l_cell_reg[88] = inform_L[88][1];				l_cell_reg[89] = inform_L[89][1];				l_cell_reg[90] = inform_L[90][1];				l_cell_reg[91] = inform_L[91][1];				l_cell_reg[92] = inform_L[92][1];				l_cell_reg[93] = inform_L[93][1];				l_cell_reg[94] = inform_L[94][1];				l_cell_reg[95] = inform_L[95][1];				l_cell_reg[96] = inform_L[96][1];				l_cell_reg[97] = inform_L[97][1];				l_cell_reg[98] = inform_L[98][1];				l_cell_reg[99] = inform_L[99][1];				l_cell_reg[100] = inform_L[100][1];				l_cell_reg[101] = inform_L[101][1];				l_cell_reg[102] = inform_L[102][1];				l_cell_reg[103] = inform_L[103][1];				l_cell_reg[104] = inform_L[104][1];				l_cell_reg[105] = inform_L[105][1];				l_cell_reg[106] = inform_L[106][1];				l_cell_reg[107] = inform_L[107][1];				l_cell_reg[108] = inform_L[108][1];				l_cell_reg[109] = inform_L[109][1];				l_cell_reg[110] = inform_L[110][1];				l_cell_reg[111] = inform_L[111][1];				l_cell_reg[112] = inform_L[112][1];				l_cell_reg[113] = inform_L[113][1];				l_cell_reg[114] = inform_L[114][1];				l_cell_reg[115] = inform_L[115][1];				l_cell_reg[116] = inform_L[116][1];				l_cell_reg[117] = inform_L[117][1];				l_cell_reg[118] = inform_L[118][1];				l_cell_reg[119] = inform_L[119][1];				l_cell_reg[120] = inform_L[120][1];				l_cell_reg[121] = inform_L[121][1];				l_cell_reg[122] = inform_L[122][1];				l_cell_reg[123] = inform_L[123][1];				l_cell_reg[124] = inform_L[124][1];				l_cell_reg[125] = inform_L[125][1];				l_cell_reg[126] = inform_L[126][1];				l_cell_reg[127] = inform_L[127][1];			end
			2:			begin				r_cell_reg[0] = inform_R[0][1];				r_cell_reg[1] = inform_R[2][1];				r_cell_reg[2] = inform_R[1][1];				r_cell_reg[3] = inform_R[3][1];				r_cell_reg[4] = inform_R[4][1];				r_cell_reg[5] = inform_R[6][1];				r_cell_reg[6] = inform_R[5][1];				r_cell_reg[7] = inform_R[7][1];				r_cell_reg[8] = inform_R[8][1];				r_cell_reg[9] = inform_R[10][1];				r_cell_reg[10] = inform_R[9][1];				r_cell_reg[11] = inform_R[11][1];				r_cell_reg[12] = inform_R[12][1];				r_cell_reg[13] = inform_R[14][1];				r_cell_reg[14] = inform_R[13][1];				r_cell_reg[15] = inform_R[15][1];				r_cell_reg[16] = inform_R[16][1];				r_cell_reg[17] = inform_R[18][1];				r_cell_reg[18] = inform_R[17][1];				r_cell_reg[19] = inform_R[19][1];				r_cell_reg[20] = inform_R[20][1];				r_cell_reg[21] = inform_R[22][1];				r_cell_reg[22] = inform_R[21][1];				r_cell_reg[23] = inform_R[23][1];				r_cell_reg[24] = inform_R[24][1];				r_cell_reg[25] = inform_R[26][1];				r_cell_reg[26] = inform_R[25][1];				r_cell_reg[27] = inform_R[27][1];				r_cell_reg[28] = inform_R[28][1];				r_cell_reg[29] = inform_R[30][1];				r_cell_reg[30] = inform_R[29][1];				r_cell_reg[31] = inform_R[31][1];				r_cell_reg[32] = inform_R[32][1];				r_cell_reg[33] = inform_R[34][1];				r_cell_reg[34] = inform_R[33][1];				r_cell_reg[35] = inform_R[35][1];				r_cell_reg[36] = inform_R[36][1];				r_cell_reg[37] = inform_R[38][1];				r_cell_reg[38] = inform_R[37][1];				r_cell_reg[39] = inform_R[39][1];				r_cell_reg[40] = inform_R[40][1];				r_cell_reg[41] = inform_R[42][1];				r_cell_reg[42] = inform_R[41][1];				r_cell_reg[43] = inform_R[43][1];				r_cell_reg[44] = inform_R[44][1];				r_cell_reg[45] = inform_R[46][1];				r_cell_reg[46] = inform_R[45][1];				r_cell_reg[47] = inform_R[47][1];				r_cell_reg[48] = inform_R[48][1];				r_cell_reg[49] = inform_R[50][1];				r_cell_reg[50] = inform_R[49][1];				r_cell_reg[51] = inform_R[51][1];				r_cell_reg[52] = inform_R[52][1];				r_cell_reg[53] = inform_R[54][1];				r_cell_reg[54] = inform_R[53][1];				r_cell_reg[55] = inform_R[55][1];				r_cell_reg[56] = inform_R[56][1];				r_cell_reg[57] = inform_R[58][1];				r_cell_reg[58] = inform_R[57][1];				r_cell_reg[59] = inform_R[59][1];				r_cell_reg[60] = inform_R[60][1];				r_cell_reg[61] = inform_R[62][1];				r_cell_reg[62] = inform_R[61][1];				r_cell_reg[63] = inform_R[63][1];				r_cell_reg[64] = inform_R[64][1];				r_cell_reg[65] = inform_R[66][1];				r_cell_reg[66] = inform_R[65][1];				r_cell_reg[67] = inform_R[67][1];				r_cell_reg[68] = inform_R[68][1];				r_cell_reg[69] = inform_R[70][1];				r_cell_reg[70] = inform_R[69][1];				r_cell_reg[71] = inform_R[71][1];				r_cell_reg[72] = inform_R[72][1];				r_cell_reg[73] = inform_R[74][1];				r_cell_reg[74] = inform_R[73][1];				r_cell_reg[75] = inform_R[75][1];				r_cell_reg[76] = inform_R[76][1];				r_cell_reg[77] = inform_R[78][1];				r_cell_reg[78] = inform_R[77][1];				r_cell_reg[79] = inform_R[79][1];				r_cell_reg[80] = inform_R[80][1];				r_cell_reg[81] = inform_R[82][1];				r_cell_reg[82] = inform_R[81][1];				r_cell_reg[83] = inform_R[83][1];				r_cell_reg[84] = inform_R[84][1];				r_cell_reg[85] = inform_R[86][1];				r_cell_reg[86] = inform_R[85][1];				r_cell_reg[87] = inform_R[87][1];				r_cell_reg[88] = inform_R[88][1];				r_cell_reg[89] = inform_R[90][1];				r_cell_reg[90] = inform_R[89][1];				r_cell_reg[91] = inform_R[91][1];				r_cell_reg[92] = inform_R[92][1];				r_cell_reg[93] = inform_R[94][1];				r_cell_reg[94] = inform_R[93][1];				r_cell_reg[95] = inform_R[95][1];				r_cell_reg[96] = inform_R[96][1];				r_cell_reg[97] = inform_R[98][1];				r_cell_reg[98] = inform_R[97][1];				r_cell_reg[99] = inform_R[99][1];				r_cell_reg[100] = inform_R[100][1];				r_cell_reg[101] = inform_R[102][1];				r_cell_reg[102] = inform_R[101][1];				r_cell_reg[103] = inform_R[103][1];				r_cell_reg[104] = inform_R[104][1];				r_cell_reg[105] = inform_R[106][1];				r_cell_reg[106] = inform_R[105][1];				r_cell_reg[107] = inform_R[107][1];				r_cell_reg[108] = inform_R[108][1];				r_cell_reg[109] = inform_R[110][1];				r_cell_reg[110] = inform_R[109][1];				r_cell_reg[111] = inform_R[111][1];				r_cell_reg[112] = inform_R[112][1];				r_cell_reg[113] = inform_R[114][1];				r_cell_reg[114] = inform_R[113][1];				r_cell_reg[115] = inform_R[115][1];				r_cell_reg[116] = inform_R[116][1];				r_cell_reg[117] = inform_R[118][1];				r_cell_reg[118] = inform_R[117][1];				r_cell_reg[119] = inform_R[119][1];				r_cell_reg[120] = inform_R[120][1];				r_cell_reg[121] = inform_R[122][1];				r_cell_reg[122] = inform_R[121][1];				r_cell_reg[123] = inform_R[123][1];				r_cell_reg[124] = inform_R[124][1];				r_cell_reg[125] = inform_R[126][1];				r_cell_reg[126] = inform_R[125][1];				r_cell_reg[127] = inform_R[127][1];				l_cell_reg[0] = inform_L[0][2];				l_cell_reg[1] = inform_L[2][2];				l_cell_reg[2] = inform_L[1][2];				l_cell_reg[3] = inform_L[3][2];				l_cell_reg[4] = inform_L[4][2];				l_cell_reg[5] = inform_L[6][2];				l_cell_reg[6] = inform_L[5][2];				l_cell_reg[7] = inform_L[7][2];				l_cell_reg[8] = inform_L[8][2];				l_cell_reg[9] = inform_L[10][2];				l_cell_reg[10] = inform_L[9][2];				l_cell_reg[11] = inform_L[11][2];				l_cell_reg[12] = inform_L[12][2];				l_cell_reg[13] = inform_L[14][2];				l_cell_reg[14] = inform_L[13][2];				l_cell_reg[15] = inform_L[15][2];				l_cell_reg[16] = inform_L[16][2];				l_cell_reg[17] = inform_L[18][2];				l_cell_reg[18] = inform_L[17][2];				l_cell_reg[19] = inform_L[19][2];				l_cell_reg[20] = inform_L[20][2];				l_cell_reg[21] = inform_L[22][2];				l_cell_reg[22] = inform_L[21][2];				l_cell_reg[23] = inform_L[23][2];				l_cell_reg[24] = inform_L[24][2];				l_cell_reg[25] = inform_L[26][2];				l_cell_reg[26] = inform_L[25][2];				l_cell_reg[27] = inform_L[27][2];				l_cell_reg[28] = inform_L[28][2];				l_cell_reg[29] = inform_L[30][2];				l_cell_reg[30] = inform_L[29][2];				l_cell_reg[31] = inform_L[31][2];				l_cell_reg[32] = inform_L[32][2];				l_cell_reg[33] = inform_L[34][2];				l_cell_reg[34] = inform_L[33][2];				l_cell_reg[35] = inform_L[35][2];				l_cell_reg[36] = inform_L[36][2];				l_cell_reg[37] = inform_L[38][2];				l_cell_reg[38] = inform_L[37][2];				l_cell_reg[39] = inform_L[39][2];				l_cell_reg[40] = inform_L[40][2];				l_cell_reg[41] = inform_L[42][2];				l_cell_reg[42] = inform_L[41][2];				l_cell_reg[43] = inform_L[43][2];				l_cell_reg[44] = inform_L[44][2];				l_cell_reg[45] = inform_L[46][2];				l_cell_reg[46] = inform_L[45][2];				l_cell_reg[47] = inform_L[47][2];				l_cell_reg[48] = inform_L[48][2];				l_cell_reg[49] = inform_L[50][2];				l_cell_reg[50] = inform_L[49][2];				l_cell_reg[51] = inform_L[51][2];				l_cell_reg[52] = inform_L[52][2];				l_cell_reg[53] = inform_L[54][2];				l_cell_reg[54] = inform_L[53][2];				l_cell_reg[55] = inform_L[55][2];				l_cell_reg[56] = inform_L[56][2];				l_cell_reg[57] = inform_L[58][2];				l_cell_reg[58] = inform_L[57][2];				l_cell_reg[59] = inform_L[59][2];				l_cell_reg[60] = inform_L[60][2];				l_cell_reg[61] = inform_L[62][2];				l_cell_reg[62] = inform_L[61][2];				l_cell_reg[63] = inform_L[63][2];				l_cell_reg[64] = inform_L[64][2];				l_cell_reg[65] = inform_L[66][2];				l_cell_reg[66] = inform_L[65][2];				l_cell_reg[67] = inform_L[67][2];				l_cell_reg[68] = inform_L[68][2];				l_cell_reg[69] = inform_L[70][2];				l_cell_reg[70] = inform_L[69][2];				l_cell_reg[71] = inform_L[71][2];				l_cell_reg[72] = inform_L[72][2];				l_cell_reg[73] = inform_L[74][2];				l_cell_reg[74] = inform_L[73][2];				l_cell_reg[75] = inform_L[75][2];				l_cell_reg[76] = inform_L[76][2];				l_cell_reg[77] = inform_L[78][2];				l_cell_reg[78] = inform_L[77][2];				l_cell_reg[79] = inform_L[79][2];				l_cell_reg[80] = inform_L[80][2];				l_cell_reg[81] = inform_L[82][2];				l_cell_reg[82] = inform_L[81][2];				l_cell_reg[83] = inform_L[83][2];				l_cell_reg[84] = inform_L[84][2];				l_cell_reg[85] = inform_L[86][2];				l_cell_reg[86] = inform_L[85][2];				l_cell_reg[87] = inform_L[87][2];				l_cell_reg[88] = inform_L[88][2];				l_cell_reg[89] = inform_L[90][2];				l_cell_reg[90] = inform_L[89][2];				l_cell_reg[91] = inform_L[91][2];				l_cell_reg[92] = inform_L[92][2];				l_cell_reg[93] = inform_L[94][2];				l_cell_reg[94] = inform_L[93][2];				l_cell_reg[95] = inform_L[95][2];				l_cell_reg[96] = inform_L[96][2];				l_cell_reg[97] = inform_L[98][2];				l_cell_reg[98] = inform_L[97][2];				l_cell_reg[99] = inform_L[99][2];				l_cell_reg[100] = inform_L[100][2];				l_cell_reg[101] = inform_L[102][2];				l_cell_reg[102] = inform_L[101][2];				l_cell_reg[103] = inform_L[103][2];				l_cell_reg[104] = inform_L[104][2];				l_cell_reg[105] = inform_L[106][2];				l_cell_reg[106] = inform_L[105][2];				l_cell_reg[107] = inform_L[107][2];				l_cell_reg[108] = inform_L[108][2];				l_cell_reg[109] = inform_L[110][2];				l_cell_reg[110] = inform_L[109][2];				l_cell_reg[111] = inform_L[111][2];				l_cell_reg[112] = inform_L[112][2];				l_cell_reg[113] = inform_L[114][2];				l_cell_reg[114] = inform_L[113][2];				l_cell_reg[115] = inform_L[115][2];				l_cell_reg[116] = inform_L[116][2];				l_cell_reg[117] = inform_L[118][2];				l_cell_reg[118] = inform_L[117][2];				l_cell_reg[119] = inform_L[119][2];				l_cell_reg[120] = inform_L[120][2];				l_cell_reg[121] = inform_L[122][2];				l_cell_reg[122] = inform_L[121][2];				l_cell_reg[123] = inform_L[123][2];				l_cell_reg[124] = inform_L[124][2];				l_cell_reg[125] = inform_L[126][2];				l_cell_reg[126] = inform_L[125][2];				l_cell_reg[127] = inform_L[127][2];			end
			3:			begin				r_cell_reg[0] = inform_R[0][2];				r_cell_reg[1] = inform_R[4][2];				r_cell_reg[2] = inform_R[1][2];				r_cell_reg[3] = inform_R[5][2];				r_cell_reg[4] = inform_R[2][2];				r_cell_reg[5] = inform_R[6][2];				r_cell_reg[6] = inform_R[3][2];				r_cell_reg[7] = inform_R[7][2];				r_cell_reg[8] = inform_R[8][2];				r_cell_reg[9] = inform_R[12][2];				r_cell_reg[10] = inform_R[9][2];				r_cell_reg[11] = inform_R[13][2];				r_cell_reg[12] = inform_R[10][2];				r_cell_reg[13] = inform_R[14][2];				r_cell_reg[14] = inform_R[11][2];				r_cell_reg[15] = inform_R[15][2];				r_cell_reg[16] = inform_R[16][2];				r_cell_reg[17] = inform_R[20][2];				r_cell_reg[18] = inform_R[17][2];				r_cell_reg[19] = inform_R[21][2];				r_cell_reg[20] = inform_R[18][2];				r_cell_reg[21] = inform_R[22][2];				r_cell_reg[22] = inform_R[19][2];				r_cell_reg[23] = inform_R[23][2];				r_cell_reg[24] = inform_R[24][2];				r_cell_reg[25] = inform_R[28][2];				r_cell_reg[26] = inform_R[25][2];				r_cell_reg[27] = inform_R[29][2];				r_cell_reg[28] = inform_R[26][2];				r_cell_reg[29] = inform_R[30][2];				r_cell_reg[30] = inform_R[27][2];				r_cell_reg[31] = inform_R[31][2];				r_cell_reg[32] = inform_R[32][2];				r_cell_reg[33] = inform_R[36][2];				r_cell_reg[34] = inform_R[33][2];				r_cell_reg[35] = inform_R[37][2];				r_cell_reg[36] = inform_R[34][2];				r_cell_reg[37] = inform_R[38][2];				r_cell_reg[38] = inform_R[35][2];				r_cell_reg[39] = inform_R[39][2];				r_cell_reg[40] = inform_R[40][2];				r_cell_reg[41] = inform_R[44][2];				r_cell_reg[42] = inform_R[41][2];				r_cell_reg[43] = inform_R[45][2];				r_cell_reg[44] = inform_R[42][2];				r_cell_reg[45] = inform_R[46][2];				r_cell_reg[46] = inform_R[43][2];				r_cell_reg[47] = inform_R[47][2];				r_cell_reg[48] = inform_R[48][2];				r_cell_reg[49] = inform_R[52][2];				r_cell_reg[50] = inform_R[49][2];				r_cell_reg[51] = inform_R[53][2];				r_cell_reg[52] = inform_R[50][2];				r_cell_reg[53] = inform_R[54][2];				r_cell_reg[54] = inform_R[51][2];				r_cell_reg[55] = inform_R[55][2];				r_cell_reg[56] = inform_R[56][2];				r_cell_reg[57] = inform_R[60][2];				r_cell_reg[58] = inform_R[57][2];				r_cell_reg[59] = inform_R[61][2];				r_cell_reg[60] = inform_R[58][2];				r_cell_reg[61] = inform_R[62][2];				r_cell_reg[62] = inform_R[59][2];				r_cell_reg[63] = inform_R[63][2];				r_cell_reg[64] = inform_R[64][2];				r_cell_reg[65] = inform_R[68][2];				r_cell_reg[66] = inform_R[65][2];				r_cell_reg[67] = inform_R[69][2];				r_cell_reg[68] = inform_R[66][2];				r_cell_reg[69] = inform_R[70][2];				r_cell_reg[70] = inform_R[67][2];				r_cell_reg[71] = inform_R[71][2];				r_cell_reg[72] = inform_R[72][2];				r_cell_reg[73] = inform_R[76][2];				r_cell_reg[74] = inform_R[73][2];				r_cell_reg[75] = inform_R[77][2];				r_cell_reg[76] = inform_R[74][2];				r_cell_reg[77] = inform_R[78][2];				r_cell_reg[78] = inform_R[75][2];				r_cell_reg[79] = inform_R[79][2];				r_cell_reg[80] = inform_R[80][2];				r_cell_reg[81] = inform_R[84][2];				r_cell_reg[82] = inform_R[81][2];				r_cell_reg[83] = inform_R[85][2];				r_cell_reg[84] = inform_R[82][2];				r_cell_reg[85] = inform_R[86][2];				r_cell_reg[86] = inform_R[83][2];				r_cell_reg[87] = inform_R[87][2];				r_cell_reg[88] = inform_R[88][2];				r_cell_reg[89] = inform_R[92][2];				r_cell_reg[90] = inform_R[89][2];				r_cell_reg[91] = inform_R[93][2];				r_cell_reg[92] = inform_R[90][2];				r_cell_reg[93] = inform_R[94][2];				r_cell_reg[94] = inform_R[91][2];				r_cell_reg[95] = inform_R[95][2];				r_cell_reg[96] = inform_R[96][2];				r_cell_reg[97] = inform_R[100][2];				r_cell_reg[98] = inform_R[97][2];				r_cell_reg[99] = inform_R[101][2];				r_cell_reg[100] = inform_R[98][2];				r_cell_reg[101] = inform_R[102][2];				r_cell_reg[102] = inform_R[99][2];				r_cell_reg[103] = inform_R[103][2];				r_cell_reg[104] = inform_R[104][2];				r_cell_reg[105] = inform_R[108][2];				r_cell_reg[106] = inform_R[105][2];				r_cell_reg[107] = inform_R[109][2];				r_cell_reg[108] = inform_R[106][2];				r_cell_reg[109] = inform_R[110][2];				r_cell_reg[110] = inform_R[107][2];				r_cell_reg[111] = inform_R[111][2];				r_cell_reg[112] = inform_R[112][2];				r_cell_reg[113] = inform_R[116][2];				r_cell_reg[114] = inform_R[113][2];				r_cell_reg[115] = inform_R[117][2];				r_cell_reg[116] = inform_R[114][2];				r_cell_reg[117] = inform_R[118][2];				r_cell_reg[118] = inform_R[115][2];				r_cell_reg[119] = inform_R[119][2];				r_cell_reg[120] = inform_R[120][2];				r_cell_reg[121] = inform_R[124][2];				r_cell_reg[122] = inform_R[121][2];				r_cell_reg[123] = inform_R[125][2];				r_cell_reg[124] = inform_R[122][2];				r_cell_reg[125] = inform_R[126][2];				r_cell_reg[126] = inform_R[123][2];				r_cell_reg[127] = inform_R[127][2];				l_cell_reg[0] = inform_L[0][3];				l_cell_reg[1] = inform_L[4][3];				l_cell_reg[2] = inform_L[1][3];				l_cell_reg[3] = inform_L[5][3];				l_cell_reg[4] = inform_L[2][3];				l_cell_reg[5] = inform_L[6][3];				l_cell_reg[6] = inform_L[3][3];				l_cell_reg[7] = inform_L[7][3];				l_cell_reg[8] = inform_L[8][3];				l_cell_reg[9] = inform_L[12][3];				l_cell_reg[10] = inform_L[9][3];				l_cell_reg[11] = inform_L[13][3];				l_cell_reg[12] = inform_L[10][3];				l_cell_reg[13] = inform_L[14][3];				l_cell_reg[14] = inform_L[11][3];				l_cell_reg[15] = inform_L[15][3];				l_cell_reg[16] = inform_L[16][3];				l_cell_reg[17] = inform_L[20][3];				l_cell_reg[18] = inform_L[17][3];				l_cell_reg[19] = inform_L[21][3];				l_cell_reg[20] = inform_L[18][3];				l_cell_reg[21] = inform_L[22][3];				l_cell_reg[22] = inform_L[19][3];				l_cell_reg[23] = inform_L[23][3];				l_cell_reg[24] = inform_L[24][3];				l_cell_reg[25] = inform_L[28][3];				l_cell_reg[26] = inform_L[25][3];				l_cell_reg[27] = inform_L[29][3];				l_cell_reg[28] = inform_L[26][3];				l_cell_reg[29] = inform_L[30][3];				l_cell_reg[30] = inform_L[27][3];				l_cell_reg[31] = inform_L[31][3];				l_cell_reg[32] = inform_L[32][3];				l_cell_reg[33] = inform_L[36][3];				l_cell_reg[34] = inform_L[33][3];				l_cell_reg[35] = inform_L[37][3];				l_cell_reg[36] = inform_L[34][3];				l_cell_reg[37] = inform_L[38][3];				l_cell_reg[38] = inform_L[35][3];				l_cell_reg[39] = inform_L[39][3];				l_cell_reg[40] = inform_L[40][3];				l_cell_reg[41] = inform_L[44][3];				l_cell_reg[42] = inform_L[41][3];				l_cell_reg[43] = inform_L[45][3];				l_cell_reg[44] = inform_L[42][3];				l_cell_reg[45] = inform_L[46][3];				l_cell_reg[46] = inform_L[43][3];				l_cell_reg[47] = inform_L[47][3];				l_cell_reg[48] = inform_L[48][3];				l_cell_reg[49] = inform_L[52][3];				l_cell_reg[50] = inform_L[49][3];				l_cell_reg[51] = inform_L[53][3];				l_cell_reg[52] = inform_L[50][3];				l_cell_reg[53] = inform_L[54][3];				l_cell_reg[54] = inform_L[51][3];				l_cell_reg[55] = inform_L[55][3];				l_cell_reg[56] = inform_L[56][3];				l_cell_reg[57] = inform_L[60][3];				l_cell_reg[58] = inform_L[57][3];				l_cell_reg[59] = inform_L[61][3];				l_cell_reg[60] = inform_L[58][3];				l_cell_reg[61] = inform_L[62][3];				l_cell_reg[62] = inform_L[59][3];				l_cell_reg[63] = inform_L[63][3];				l_cell_reg[64] = inform_L[64][3];				l_cell_reg[65] = inform_L[68][3];				l_cell_reg[66] = inform_L[65][3];				l_cell_reg[67] = inform_L[69][3];				l_cell_reg[68] = inform_L[66][3];				l_cell_reg[69] = inform_L[70][3];				l_cell_reg[70] = inform_L[67][3];				l_cell_reg[71] = inform_L[71][3];				l_cell_reg[72] = inform_L[72][3];				l_cell_reg[73] = inform_L[76][3];				l_cell_reg[74] = inform_L[73][3];				l_cell_reg[75] = inform_L[77][3];				l_cell_reg[76] = inform_L[74][3];				l_cell_reg[77] = inform_L[78][3];				l_cell_reg[78] = inform_L[75][3];				l_cell_reg[79] = inform_L[79][3];				l_cell_reg[80] = inform_L[80][3];				l_cell_reg[81] = inform_L[84][3];				l_cell_reg[82] = inform_L[81][3];				l_cell_reg[83] = inform_L[85][3];				l_cell_reg[84] = inform_L[82][3];				l_cell_reg[85] = inform_L[86][3];				l_cell_reg[86] = inform_L[83][3];				l_cell_reg[87] = inform_L[87][3];				l_cell_reg[88] = inform_L[88][3];				l_cell_reg[89] = inform_L[92][3];				l_cell_reg[90] = inform_L[89][3];				l_cell_reg[91] = inform_L[93][3];				l_cell_reg[92] = inform_L[90][3];				l_cell_reg[93] = inform_L[94][3];				l_cell_reg[94] = inform_L[91][3];				l_cell_reg[95] = inform_L[95][3];				l_cell_reg[96] = inform_L[96][3];				l_cell_reg[97] = inform_L[100][3];				l_cell_reg[98] = inform_L[97][3];				l_cell_reg[99] = inform_L[101][3];				l_cell_reg[100] = inform_L[98][3];				l_cell_reg[101] = inform_L[102][3];				l_cell_reg[102] = inform_L[99][3];				l_cell_reg[103] = inform_L[103][3];				l_cell_reg[104] = inform_L[104][3];				l_cell_reg[105] = inform_L[108][3];				l_cell_reg[106] = inform_L[105][3];				l_cell_reg[107] = inform_L[109][3];				l_cell_reg[108] = inform_L[106][3];				l_cell_reg[109] = inform_L[110][3];				l_cell_reg[110] = inform_L[107][3];				l_cell_reg[111] = inform_L[111][3];				l_cell_reg[112] = inform_L[112][3];				l_cell_reg[113] = inform_L[116][3];				l_cell_reg[114] = inform_L[113][3];				l_cell_reg[115] = inform_L[117][3];				l_cell_reg[116] = inform_L[114][3];				l_cell_reg[117] = inform_L[118][3];				l_cell_reg[118] = inform_L[115][3];				l_cell_reg[119] = inform_L[119][3];				l_cell_reg[120] = inform_L[120][3];				l_cell_reg[121] = inform_L[124][3];				l_cell_reg[122] = inform_L[121][3];				l_cell_reg[123] = inform_L[125][3];				l_cell_reg[124] = inform_L[122][3];				l_cell_reg[125] = inform_L[126][3];				l_cell_reg[126] = inform_L[123][3];				l_cell_reg[127] = inform_L[127][3];			end
			4:			begin				r_cell_reg[0] = inform_R[0][3];				r_cell_reg[1] = inform_R[8][3];				r_cell_reg[2] = inform_R[1][3];				r_cell_reg[3] = inform_R[9][3];				r_cell_reg[4] = inform_R[2][3];				r_cell_reg[5] = inform_R[10][3];				r_cell_reg[6] = inform_R[3][3];				r_cell_reg[7] = inform_R[11][3];				r_cell_reg[8] = inform_R[4][3];				r_cell_reg[9] = inform_R[12][3];				r_cell_reg[10] = inform_R[5][3];				r_cell_reg[11] = inform_R[13][3];				r_cell_reg[12] = inform_R[6][3];				r_cell_reg[13] = inform_R[14][3];				r_cell_reg[14] = inform_R[7][3];				r_cell_reg[15] = inform_R[15][3];				r_cell_reg[16] = inform_R[16][3];				r_cell_reg[17] = inform_R[24][3];				r_cell_reg[18] = inform_R[17][3];				r_cell_reg[19] = inform_R[25][3];				r_cell_reg[20] = inform_R[18][3];				r_cell_reg[21] = inform_R[26][3];				r_cell_reg[22] = inform_R[19][3];				r_cell_reg[23] = inform_R[27][3];				r_cell_reg[24] = inform_R[20][3];				r_cell_reg[25] = inform_R[28][3];				r_cell_reg[26] = inform_R[21][3];				r_cell_reg[27] = inform_R[29][3];				r_cell_reg[28] = inform_R[22][3];				r_cell_reg[29] = inform_R[30][3];				r_cell_reg[30] = inform_R[23][3];				r_cell_reg[31] = inform_R[31][3];				r_cell_reg[32] = inform_R[32][3];				r_cell_reg[33] = inform_R[40][3];				r_cell_reg[34] = inform_R[33][3];				r_cell_reg[35] = inform_R[41][3];				r_cell_reg[36] = inform_R[34][3];				r_cell_reg[37] = inform_R[42][3];				r_cell_reg[38] = inform_R[35][3];				r_cell_reg[39] = inform_R[43][3];				r_cell_reg[40] = inform_R[36][3];				r_cell_reg[41] = inform_R[44][3];				r_cell_reg[42] = inform_R[37][3];				r_cell_reg[43] = inform_R[45][3];				r_cell_reg[44] = inform_R[38][3];				r_cell_reg[45] = inform_R[46][3];				r_cell_reg[46] = inform_R[39][3];				r_cell_reg[47] = inform_R[47][3];				r_cell_reg[48] = inform_R[48][3];				r_cell_reg[49] = inform_R[56][3];				r_cell_reg[50] = inform_R[49][3];				r_cell_reg[51] = inform_R[57][3];				r_cell_reg[52] = inform_R[50][3];				r_cell_reg[53] = inform_R[58][3];				r_cell_reg[54] = inform_R[51][3];				r_cell_reg[55] = inform_R[59][3];				r_cell_reg[56] = inform_R[52][3];				r_cell_reg[57] = inform_R[60][3];				r_cell_reg[58] = inform_R[53][3];				r_cell_reg[59] = inform_R[61][3];				r_cell_reg[60] = inform_R[54][3];				r_cell_reg[61] = inform_R[62][3];				r_cell_reg[62] = inform_R[55][3];				r_cell_reg[63] = inform_R[63][3];				r_cell_reg[64] = inform_R[64][3];				r_cell_reg[65] = inform_R[72][3];				r_cell_reg[66] = inform_R[65][3];				r_cell_reg[67] = inform_R[73][3];				r_cell_reg[68] = inform_R[66][3];				r_cell_reg[69] = inform_R[74][3];				r_cell_reg[70] = inform_R[67][3];				r_cell_reg[71] = inform_R[75][3];				r_cell_reg[72] = inform_R[68][3];				r_cell_reg[73] = inform_R[76][3];				r_cell_reg[74] = inform_R[69][3];				r_cell_reg[75] = inform_R[77][3];				r_cell_reg[76] = inform_R[70][3];				r_cell_reg[77] = inform_R[78][3];				r_cell_reg[78] = inform_R[71][3];				r_cell_reg[79] = inform_R[79][3];				r_cell_reg[80] = inform_R[80][3];				r_cell_reg[81] = inform_R[88][3];				r_cell_reg[82] = inform_R[81][3];				r_cell_reg[83] = inform_R[89][3];				r_cell_reg[84] = inform_R[82][3];				r_cell_reg[85] = inform_R[90][3];				r_cell_reg[86] = inform_R[83][3];				r_cell_reg[87] = inform_R[91][3];				r_cell_reg[88] = inform_R[84][3];				r_cell_reg[89] = inform_R[92][3];				r_cell_reg[90] = inform_R[85][3];				r_cell_reg[91] = inform_R[93][3];				r_cell_reg[92] = inform_R[86][3];				r_cell_reg[93] = inform_R[94][3];				r_cell_reg[94] = inform_R[87][3];				r_cell_reg[95] = inform_R[95][3];				r_cell_reg[96] = inform_R[96][3];				r_cell_reg[97] = inform_R[104][3];				r_cell_reg[98] = inform_R[97][3];				r_cell_reg[99] = inform_R[105][3];				r_cell_reg[100] = inform_R[98][3];				r_cell_reg[101] = inform_R[106][3];				r_cell_reg[102] = inform_R[99][3];				r_cell_reg[103] = inform_R[107][3];				r_cell_reg[104] = inform_R[100][3];				r_cell_reg[105] = inform_R[108][3];				r_cell_reg[106] = inform_R[101][3];				r_cell_reg[107] = inform_R[109][3];				r_cell_reg[108] = inform_R[102][3];				r_cell_reg[109] = inform_R[110][3];				r_cell_reg[110] = inform_R[103][3];				r_cell_reg[111] = inform_R[111][3];				r_cell_reg[112] = inform_R[112][3];				r_cell_reg[113] = inform_R[120][3];				r_cell_reg[114] = inform_R[113][3];				r_cell_reg[115] = inform_R[121][3];				r_cell_reg[116] = inform_R[114][3];				r_cell_reg[117] = inform_R[122][3];				r_cell_reg[118] = inform_R[115][3];				r_cell_reg[119] = inform_R[123][3];				r_cell_reg[120] = inform_R[116][3];				r_cell_reg[121] = inform_R[124][3];				r_cell_reg[122] = inform_R[117][3];				r_cell_reg[123] = inform_R[125][3];				r_cell_reg[124] = inform_R[118][3];				r_cell_reg[125] = inform_R[126][3];				r_cell_reg[126] = inform_R[119][3];				r_cell_reg[127] = inform_R[127][3];				l_cell_reg[0] = inform_L[0][4];				l_cell_reg[1] = inform_L[8][4];				l_cell_reg[2] = inform_L[1][4];				l_cell_reg[3] = inform_L[9][4];				l_cell_reg[4] = inform_L[2][4];				l_cell_reg[5] = inform_L[10][4];				l_cell_reg[6] = inform_L[3][4];				l_cell_reg[7] = inform_L[11][4];				l_cell_reg[8] = inform_L[4][4];				l_cell_reg[9] = inform_L[12][4];				l_cell_reg[10] = inform_L[5][4];				l_cell_reg[11] = inform_L[13][4];				l_cell_reg[12] = inform_L[6][4];				l_cell_reg[13] = inform_L[14][4];				l_cell_reg[14] = inform_L[7][4];				l_cell_reg[15] = inform_L[15][4];				l_cell_reg[16] = inform_L[16][4];				l_cell_reg[17] = inform_L[24][4];				l_cell_reg[18] = inform_L[17][4];				l_cell_reg[19] = inform_L[25][4];				l_cell_reg[20] = inform_L[18][4];				l_cell_reg[21] = inform_L[26][4];				l_cell_reg[22] = inform_L[19][4];				l_cell_reg[23] = inform_L[27][4];				l_cell_reg[24] = inform_L[20][4];				l_cell_reg[25] = inform_L[28][4];				l_cell_reg[26] = inform_L[21][4];				l_cell_reg[27] = inform_L[29][4];				l_cell_reg[28] = inform_L[22][4];				l_cell_reg[29] = inform_L[30][4];				l_cell_reg[30] = inform_L[23][4];				l_cell_reg[31] = inform_L[31][4];				l_cell_reg[32] = inform_L[32][4];				l_cell_reg[33] = inform_L[40][4];				l_cell_reg[34] = inform_L[33][4];				l_cell_reg[35] = inform_L[41][4];				l_cell_reg[36] = inform_L[34][4];				l_cell_reg[37] = inform_L[42][4];				l_cell_reg[38] = inform_L[35][4];				l_cell_reg[39] = inform_L[43][4];				l_cell_reg[40] = inform_L[36][4];				l_cell_reg[41] = inform_L[44][4];				l_cell_reg[42] = inform_L[37][4];				l_cell_reg[43] = inform_L[45][4];				l_cell_reg[44] = inform_L[38][4];				l_cell_reg[45] = inform_L[46][4];				l_cell_reg[46] = inform_L[39][4];				l_cell_reg[47] = inform_L[47][4];				l_cell_reg[48] = inform_L[48][4];				l_cell_reg[49] = inform_L[56][4];				l_cell_reg[50] = inform_L[49][4];				l_cell_reg[51] = inform_L[57][4];				l_cell_reg[52] = inform_L[50][4];				l_cell_reg[53] = inform_L[58][4];				l_cell_reg[54] = inform_L[51][4];				l_cell_reg[55] = inform_L[59][4];				l_cell_reg[56] = inform_L[52][4];				l_cell_reg[57] = inform_L[60][4];				l_cell_reg[58] = inform_L[53][4];				l_cell_reg[59] = inform_L[61][4];				l_cell_reg[60] = inform_L[54][4];				l_cell_reg[61] = inform_L[62][4];				l_cell_reg[62] = inform_L[55][4];				l_cell_reg[63] = inform_L[63][4];				l_cell_reg[64] = inform_L[64][4];				l_cell_reg[65] = inform_L[72][4];				l_cell_reg[66] = inform_L[65][4];				l_cell_reg[67] = inform_L[73][4];				l_cell_reg[68] = inform_L[66][4];				l_cell_reg[69] = inform_L[74][4];				l_cell_reg[70] = inform_L[67][4];				l_cell_reg[71] = inform_L[75][4];				l_cell_reg[72] = inform_L[68][4];				l_cell_reg[73] = inform_L[76][4];				l_cell_reg[74] = inform_L[69][4];				l_cell_reg[75] = inform_L[77][4];				l_cell_reg[76] = inform_L[70][4];				l_cell_reg[77] = inform_L[78][4];				l_cell_reg[78] = inform_L[71][4];				l_cell_reg[79] = inform_L[79][4];				l_cell_reg[80] = inform_L[80][4];				l_cell_reg[81] = inform_L[88][4];				l_cell_reg[82] = inform_L[81][4];				l_cell_reg[83] = inform_L[89][4];				l_cell_reg[84] = inform_L[82][4];				l_cell_reg[85] = inform_L[90][4];				l_cell_reg[86] = inform_L[83][4];				l_cell_reg[87] = inform_L[91][4];				l_cell_reg[88] = inform_L[84][4];				l_cell_reg[89] = inform_L[92][4];				l_cell_reg[90] = inform_L[85][4];				l_cell_reg[91] = inform_L[93][4];				l_cell_reg[92] = inform_L[86][4];				l_cell_reg[93] = inform_L[94][4];				l_cell_reg[94] = inform_L[87][4];				l_cell_reg[95] = inform_L[95][4];				l_cell_reg[96] = inform_L[96][4];				l_cell_reg[97] = inform_L[104][4];				l_cell_reg[98] = inform_L[97][4];				l_cell_reg[99] = inform_L[105][4];				l_cell_reg[100] = inform_L[98][4];				l_cell_reg[101] = inform_L[106][4];				l_cell_reg[102] = inform_L[99][4];				l_cell_reg[103] = inform_L[107][4];				l_cell_reg[104] = inform_L[100][4];				l_cell_reg[105] = inform_L[108][4];				l_cell_reg[106] = inform_L[101][4];				l_cell_reg[107] = inform_L[109][4];				l_cell_reg[108] = inform_L[102][4];				l_cell_reg[109] = inform_L[110][4];				l_cell_reg[110] = inform_L[103][4];				l_cell_reg[111] = inform_L[111][4];				l_cell_reg[112] = inform_L[112][4];				l_cell_reg[113] = inform_L[120][4];				l_cell_reg[114] = inform_L[113][4];				l_cell_reg[115] = inform_L[121][4];				l_cell_reg[116] = inform_L[114][4];				l_cell_reg[117] = inform_L[122][4];				l_cell_reg[118] = inform_L[115][4];				l_cell_reg[119] = inform_L[123][4];				l_cell_reg[120] = inform_L[116][4];				l_cell_reg[121] = inform_L[124][4];				l_cell_reg[122] = inform_L[117][4];				l_cell_reg[123] = inform_L[125][4];				l_cell_reg[124] = inform_L[118][4];				l_cell_reg[125] = inform_L[126][4];				l_cell_reg[126] = inform_L[119][4];				l_cell_reg[127] = inform_L[127][4];			end
			5:			begin				r_cell_reg[0] = inform_R[0][4];				r_cell_reg[1] = inform_R[16][4];				r_cell_reg[2] = inform_R[1][4];				r_cell_reg[3] = inform_R[17][4];				r_cell_reg[4] = inform_R[2][4];				r_cell_reg[5] = inform_R[18][4];				r_cell_reg[6] = inform_R[3][4];				r_cell_reg[7] = inform_R[19][4];				r_cell_reg[8] = inform_R[4][4];				r_cell_reg[9] = inform_R[20][4];				r_cell_reg[10] = inform_R[5][4];				r_cell_reg[11] = inform_R[21][4];				r_cell_reg[12] = inform_R[6][4];				r_cell_reg[13] = inform_R[22][4];				r_cell_reg[14] = inform_R[7][4];				r_cell_reg[15] = inform_R[23][4];				r_cell_reg[16] = inform_R[8][4];				r_cell_reg[17] = inform_R[24][4];				r_cell_reg[18] = inform_R[9][4];				r_cell_reg[19] = inform_R[25][4];				r_cell_reg[20] = inform_R[10][4];				r_cell_reg[21] = inform_R[26][4];				r_cell_reg[22] = inform_R[11][4];				r_cell_reg[23] = inform_R[27][4];				r_cell_reg[24] = inform_R[12][4];				r_cell_reg[25] = inform_R[28][4];				r_cell_reg[26] = inform_R[13][4];				r_cell_reg[27] = inform_R[29][4];				r_cell_reg[28] = inform_R[14][4];				r_cell_reg[29] = inform_R[30][4];				r_cell_reg[30] = inform_R[15][4];				r_cell_reg[31] = inform_R[31][4];				r_cell_reg[32] = inform_R[32][4];				r_cell_reg[33] = inform_R[48][4];				r_cell_reg[34] = inform_R[33][4];				r_cell_reg[35] = inform_R[49][4];				r_cell_reg[36] = inform_R[34][4];				r_cell_reg[37] = inform_R[50][4];				r_cell_reg[38] = inform_R[35][4];				r_cell_reg[39] = inform_R[51][4];				r_cell_reg[40] = inform_R[36][4];				r_cell_reg[41] = inform_R[52][4];				r_cell_reg[42] = inform_R[37][4];				r_cell_reg[43] = inform_R[53][4];				r_cell_reg[44] = inform_R[38][4];				r_cell_reg[45] = inform_R[54][4];				r_cell_reg[46] = inform_R[39][4];				r_cell_reg[47] = inform_R[55][4];				r_cell_reg[48] = inform_R[40][4];				r_cell_reg[49] = inform_R[56][4];				r_cell_reg[50] = inform_R[41][4];				r_cell_reg[51] = inform_R[57][4];				r_cell_reg[52] = inform_R[42][4];				r_cell_reg[53] = inform_R[58][4];				r_cell_reg[54] = inform_R[43][4];				r_cell_reg[55] = inform_R[59][4];				r_cell_reg[56] = inform_R[44][4];				r_cell_reg[57] = inform_R[60][4];				r_cell_reg[58] = inform_R[45][4];				r_cell_reg[59] = inform_R[61][4];				r_cell_reg[60] = inform_R[46][4];				r_cell_reg[61] = inform_R[62][4];				r_cell_reg[62] = inform_R[47][4];				r_cell_reg[63] = inform_R[63][4];				r_cell_reg[64] = inform_R[64][4];				r_cell_reg[65] = inform_R[80][4];				r_cell_reg[66] = inform_R[65][4];				r_cell_reg[67] = inform_R[81][4];				r_cell_reg[68] = inform_R[66][4];				r_cell_reg[69] = inform_R[82][4];				r_cell_reg[70] = inform_R[67][4];				r_cell_reg[71] = inform_R[83][4];				r_cell_reg[72] = inform_R[68][4];				r_cell_reg[73] = inform_R[84][4];				r_cell_reg[74] = inform_R[69][4];				r_cell_reg[75] = inform_R[85][4];				r_cell_reg[76] = inform_R[70][4];				r_cell_reg[77] = inform_R[86][4];				r_cell_reg[78] = inform_R[71][4];				r_cell_reg[79] = inform_R[87][4];				r_cell_reg[80] = inform_R[72][4];				r_cell_reg[81] = inform_R[88][4];				r_cell_reg[82] = inform_R[73][4];				r_cell_reg[83] = inform_R[89][4];				r_cell_reg[84] = inform_R[74][4];				r_cell_reg[85] = inform_R[90][4];				r_cell_reg[86] = inform_R[75][4];				r_cell_reg[87] = inform_R[91][4];				r_cell_reg[88] = inform_R[76][4];				r_cell_reg[89] = inform_R[92][4];				r_cell_reg[90] = inform_R[77][4];				r_cell_reg[91] = inform_R[93][4];				r_cell_reg[92] = inform_R[78][4];				r_cell_reg[93] = inform_R[94][4];				r_cell_reg[94] = inform_R[79][4];				r_cell_reg[95] = inform_R[95][4];				r_cell_reg[96] = inform_R[96][4];				r_cell_reg[97] = inform_R[112][4];				r_cell_reg[98] = inform_R[97][4];				r_cell_reg[99] = inform_R[113][4];				r_cell_reg[100] = inform_R[98][4];				r_cell_reg[101] = inform_R[114][4];				r_cell_reg[102] = inform_R[99][4];				r_cell_reg[103] = inform_R[115][4];				r_cell_reg[104] = inform_R[100][4];				r_cell_reg[105] = inform_R[116][4];				r_cell_reg[106] = inform_R[101][4];				r_cell_reg[107] = inform_R[117][4];				r_cell_reg[108] = inform_R[102][4];				r_cell_reg[109] = inform_R[118][4];				r_cell_reg[110] = inform_R[103][4];				r_cell_reg[111] = inform_R[119][4];				r_cell_reg[112] = inform_R[104][4];				r_cell_reg[113] = inform_R[120][4];				r_cell_reg[114] = inform_R[105][4];				r_cell_reg[115] = inform_R[121][4];				r_cell_reg[116] = inform_R[106][4];				r_cell_reg[117] = inform_R[122][4];				r_cell_reg[118] = inform_R[107][4];				r_cell_reg[119] = inform_R[123][4];				r_cell_reg[120] = inform_R[108][4];				r_cell_reg[121] = inform_R[124][4];				r_cell_reg[122] = inform_R[109][4];				r_cell_reg[123] = inform_R[125][4];				r_cell_reg[124] = inform_R[110][4];				r_cell_reg[125] = inform_R[126][4];				r_cell_reg[126] = inform_R[111][4];				r_cell_reg[127] = inform_R[127][4];				l_cell_reg[0] = inform_L[0][5];				l_cell_reg[1] = inform_L[16][5];				l_cell_reg[2] = inform_L[1][5];				l_cell_reg[3] = inform_L[17][5];				l_cell_reg[4] = inform_L[2][5];				l_cell_reg[5] = inform_L[18][5];				l_cell_reg[6] = inform_L[3][5];				l_cell_reg[7] = inform_L[19][5];				l_cell_reg[8] = inform_L[4][5];				l_cell_reg[9] = inform_L[20][5];				l_cell_reg[10] = inform_L[5][5];				l_cell_reg[11] = inform_L[21][5];				l_cell_reg[12] = inform_L[6][5];				l_cell_reg[13] = inform_L[22][5];				l_cell_reg[14] = inform_L[7][5];				l_cell_reg[15] = inform_L[23][5];				l_cell_reg[16] = inform_L[8][5];				l_cell_reg[17] = inform_L[24][5];				l_cell_reg[18] = inform_L[9][5];				l_cell_reg[19] = inform_L[25][5];				l_cell_reg[20] = inform_L[10][5];				l_cell_reg[21] = inform_L[26][5];				l_cell_reg[22] = inform_L[11][5];				l_cell_reg[23] = inform_L[27][5];				l_cell_reg[24] = inform_L[12][5];				l_cell_reg[25] = inform_L[28][5];				l_cell_reg[26] = inform_L[13][5];				l_cell_reg[27] = inform_L[29][5];				l_cell_reg[28] = inform_L[14][5];				l_cell_reg[29] = inform_L[30][5];				l_cell_reg[30] = inform_L[15][5];				l_cell_reg[31] = inform_L[31][5];				l_cell_reg[32] = inform_L[32][5];				l_cell_reg[33] = inform_L[48][5];				l_cell_reg[34] = inform_L[33][5];				l_cell_reg[35] = inform_L[49][5];				l_cell_reg[36] = inform_L[34][5];				l_cell_reg[37] = inform_L[50][5];				l_cell_reg[38] = inform_L[35][5];				l_cell_reg[39] = inform_L[51][5];				l_cell_reg[40] = inform_L[36][5];				l_cell_reg[41] = inform_L[52][5];				l_cell_reg[42] = inform_L[37][5];				l_cell_reg[43] = inform_L[53][5];				l_cell_reg[44] = inform_L[38][5];				l_cell_reg[45] = inform_L[54][5];				l_cell_reg[46] = inform_L[39][5];				l_cell_reg[47] = inform_L[55][5];				l_cell_reg[48] = inform_L[40][5];				l_cell_reg[49] = inform_L[56][5];				l_cell_reg[50] = inform_L[41][5];				l_cell_reg[51] = inform_L[57][5];				l_cell_reg[52] = inform_L[42][5];				l_cell_reg[53] = inform_L[58][5];				l_cell_reg[54] = inform_L[43][5];				l_cell_reg[55] = inform_L[59][5];				l_cell_reg[56] = inform_L[44][5];				l_cell_reg[57] = inform_L[60][5];				l_cell_reg[58] = inform_L[45][5];				l_cell_reg[59] = inform_L[61][5];				l_cell_reg[60] = inform_L[46][5];				l_cell_reg[61] = inform_L[62][5];				l_cell_reg[62] = inform_L[47][5];				l_cell_reg[63] = inform_L[63][5];				l_cell_reg[64] = inform_L[64][5];				l_cell_reg[65] = inform_L[80][5];				l_cell_reg[66] = inform_L[65][5];				l_cell_reg[67] = inform_L[81][5];				l_cell_reg[68] = inform_L[66][5];				l_cell_reg[69] = inform_L[82][5];				l_cell_reg[70] = inform_L[67][5];				l_cell_reg[71] = inform_L[83][5];				l_cell_reg[72] = inform_L[68][5];				l_cell_reg[73] = inform_L[84][5];				l_cell_reg[74] = inform_L[69][5];				l_cell_reg[75] = inform_L[85][5];				l_cell_reg[76] = inform_L[70][5];				l_cell_reg[77] = inform_L[86][5];				l_cell_reg[78] = inform_L[71][5];				l_cell_reg[79] = inform_L[87][5];				l_cell_reg[80] = inform_L[72][5];				l_cell_reg[81] = inform_L[88][5];				l_cell_reg[82] = inform_L[73][5];				l_cell_reg[83] = inform_L[89][5];				l_cell_reg[84] = inform_L[74][5];				l_cell_reg[85] = inform_L[90][5];				l_cell_reg[86] = inform_L[75][5];				l_cell_reg[87] = inform_L[91][5];				l_cell_reg[88] = inform_L[76][5];				l_cell_reg[89] = inform_L[92][5];				l_cell_reg[90] = inform_L[77][5];				l_cell_reg[91] = inform_L[93][5];				l_cell_reg[92] = inform_L[78][5];				l_cell_reg[93] = inform_L[94][5];				l_cell_reg[94] = inform_L[79][5];				l_cell_reg[95] = inform_L[95][5];				l_cell_reg[96] = inform_L[96][5];				l_cell_reg[97] = inform_L[112][5];				l_cell_reg[98] = inform_L[97][5];				l_cell_reg[99] = inform_L[113][5];				l_cell_reg[100] = inform_L[98][5];				l_cell_reg[101] = inform_L[114][5];				l_cell_reg[102] = inform_L[99][5];				l_cell_reg[103] = inform_L[115][5];				l_cell_reg[104] = inform_L[100][5];				l_cell_reg[105] = inform_L[116][5];				l_cell_reg[106] = inform_L[101][5];				l_cell_reg[107] = inform_L[117][5];				l_cell_reg[108] = inform_L[102][5];				l_cell_reg[109] = inform_L[118][5];				l_cell_reg[110] = inform_L[103][5];				l_cell_reg[111] = inform_L[119][5];				l_cell_reg[112] = inform_L[104][5];				l_cell_reg[113] = inform_L[120][5];				l_cell_reg[114] = inform_L[105][5];				l_cell_reg[115] = inform_L[121][5];				l_cell_reg[116] = inform_L[106][5];				l_cell_reg[117] = inform_L[122][5];				l_cell_reg[118] = inform_L[107][5];				l_cell_reg[119] = inform_L[123][5];				l_cell_reg[120] = inform_L[108][5];				l_cell_reg[121] = inform_L[124][5];				l_cell_reg[122] = inform_L[109][5];				l_cell_reg[123] = inform_L[125][5];				l_cell_reg[124] = inform_L[110][5];				l_cell_reg[125] = inform_L[126][5];				l_cell_reg[126] = inform_L[111][5];				l_cell_reg[127] = inform_L[127][5];			end
			6:			begin				r_cell_reg[0] = inform_R[0][5];				r_cell_reg[1] = inform_R[32][5];				r_cell_reg[2] = inform_R[1][5];				r_cell_reg[3] = inform_R[33][5];				r_cell_reg[4] = inform_R[2][5];				r_cell_reg[5] = inform_R[34][5];				r_cell_reg[6] = inform_R[3][5];				r_cell_reg[7] = inform_R[35][5];				r_cell_reg[8] = inform_R[4][5];				r_cell_reg[9] = inform_R[36][5];				r_cell_reg[10] = inform_R[5][5];				r_cell_reg[11] = inform_R[37][5];				r_cell_reg[12] = inform_R[6][5];				r_cell_reg[13] = inform_R[38][5];				r_cell_reg[14] = inform_R[7][5];				r_cell_reg[15] = inform_R[39][5];				r_cell_reg[16] = inform_R[8][5];				r_cell_reg[17] = inform_R[40][5];				r_cell_reg[18] = inform_R[9][5];				r_cell_reg[19] = inform_R[41][5];				r_cell_reg[20] = inform_R[10][5];				r_cell_reg[21] = inform_R[42][5];				r_cell_reg[22] = inform_R[11][5];				r_cell_reg[23] = inform_R[43][5];				r_cell_reg[24] = inform_R[12][5];				r_cell_reg[25] = inform_R[44][5];				r_cell_reg[26] = inform_R[13][5];				r_cell_reg[27] = inform_R[45][5];				r_cell_reg[28] = inform_R[14][5];				r_cell_reg[29] = inform_R[46][5];				r_cell_reg[30] = inform_R[15][5];				r_cell_reg[31] = inform_R[47][5];				r_cell_reg[32] = inform_R[16][5];				r_cell_reg[33] = inform_R[48][5];				r_cell_reg[34] = inform_R[17][5];				r_cell_reg[35] = inform_R[49][5];				r_cell_reg[36] = inform_R[18][5];				r_cell_reg[37] = inform_R[50][5];				r_cell_reg[38] = inform_R[19][5];				r_cell_reg[39] = inform_R[51][5];				r_cell_reg[40] = inform_R[20][5];				r_cell_reg[41] = inform_R[52][5];				r_cell_reg[42] = inform_R[21][5];				r_cell_reg[43] = inform_R[53][5];				r_cell_reg[44] = inform_R[22][5];				r_cell_reg[45] = inform_R[54][5];				r_cell_reg[46] = inform_R[23][5];				r_cell_reg[47] = inform_R[55][5];				r_cell_reg[48] = inform_R[24][5];				r_cell_reg[49] = inform_R[56][5];				r_cell_reg[50] = inform_R[25][5];				r_cell_reg[51] = inform_R[57][5];				r_cell_reg[52] = inform_R[26][5];				r_cell_reg[53] = inform_R[58][5];				r_cell_reg[54] = inform_R[27][5];				r_cell_reg[55] = inform_R[59][5];				r_cell_reg[56] = inform_R[28][5];				r_cell_reg[57] = inform_R[60][5];				r_cell_reg[58] = inform_R[29][5];				r_cell_reg[59] = inform_R[61][5];				r_cell_reg[60] = inform_R[30][5];				r_cell_reg[61] = inform_R[62][5];				r_cell_reg[62] = inform_R[31][5];				r_cell_reg[63] = inform_R[63][5];				r_cell_reg[64] = inform_R[64][5];				r_cell_reg[65] = inform_R[96][5];				r_cell_reg[66] = inform_R[65][5];				r_cell_reg[67] = inform_R[97][5];				r_cell_reg[68] = inform_R[66][5];				r_cell_reg[69] = inform_R[98][5];				r_cell_reg[70] = inform_R[67][5];				r_cell_reg[71] = inform_R[99][5];				r_cell_reg[72] = inform_R[68][5];				r_cell_reg[73] = inform_R[100][5];				r_cell_reg[74] = inform_R[69][5];				r_cell_reg[75] = inform_R[101][5];				r_cell_reg[76] = inform_R[70][5];				r_cell_reg[77] = inform_R[102][5];				r_cell_reg[78] = inform_R[71][5];				r_cell_reg[79] = inform_R[103][5];				r_cell_reg[80] = inform_R[72][5];				r_cell_reg[81] = inform_R[104][5];				r_cell_reg[82] = inform_R[73][5];				r_cell_reg[83] = inform_R[105][5];				r_cell_reg[84] = inform_R[74][5];				r_cell_reg[85] = inform_R[106][5];				r_cell_reg[86] = inform_R[75][5];				r_cell_reg[87] = inform_R[107][5];				r_cell_reg[88] = inform_R[76][5];				r_cell_reg[89] = inform_R[108][5];				r_cell_reg[90] = inform_R[77][5];				r_cell_reg[91] = inform_R[109][5];				r_cell_reg[92] = inform_R[78][5];				r_cell_reg[93] = inform_R[110][5];				r_cell_reg[94] = inform_R[79][5];				r_cell_reg[95] = inform_R[111][5];				r_cell_reg[96] = inform_R[80][5];				r_cell_reg[97] = inform_R[112][5];				r_cell_reg[98] = inform_R[81][5];				r_cell_reg[99] = inform_R[113][5];				r_cell_reg[100] = inform_R[82][5];				r_cell_reg[101] = inform_R[114][5];				r_cell_reg[102] = inform_R[83][5];				r_cell_reg[103] = inform_R[115][5];				r_cell_reg[104] = inform_R[84][5];				r_cell_reg[105] = inform_R[116][5];				r_cell_reg[106] = inform_R[85][5];				r_cell_reg[107] = inform_R[117][5];				r_cell_reg[108] = inform_R[86][5];				r_cell_reg[109] = inform_R[118][5];				r_cell_reg[110] = inform_R[87][5];				r_cell_reg[111] = inform_R[119][5];				r_cell_reg[112] = inform_R[88][5];				r_cell_reg[113] = inform_R[120][5];				r_cell_reg[114] = inform_R[89][5];				r_cell_reg[115] = inform_R[121][5];				r_cell_reg[116] = inform_R[90][5];				r_cell_reg[117] = inform_R[122][5];				r_cell_reg[118] = inform_R[91][5];				r_cell_reg[119] = inform_R[123][5];				r_cell_reg[120] = inform_R[92][5];				r_cell_reg[121] = inform_R[124][5];				r_cell_reg[122] = inform_R[93][5];				r_cell_reg[123] = inform_R[125][5];				r_cell_reg[124] = inform_R[94][5];				r_cell_reg[125] = inform_R[126][5];				r_cell_reg[126] = inform_R[95][5];				r_cell_reg[127] = inform_R[127][5];				l_cell_reg[0] = inform_L[0][6];				l_cell_reg[1] = inform_L[32][6];				l_cell_reg[2] = inform_L[1][6];				l_cell_reg[3] = inform_L[33][6];				l_cell_reg[4] = inform_L[2][6];				l_cell_reg[5] = inform_L[34][6];				l_cell_reg[6] = inform_L[3][6];				l_cell_reg[7] = inform_L[35][6];				l_cell_reg[8] = inform_L[4][6];				l_cell_reg[9] = inform_L[36][6];				l_cell_reg[10] = inform_L[5][6];				l_cell_reg[11] = inform_L[37][6];				l_cell_reg[12] = inform_L[6][6];				l_cell_reg[13] = inform_L[38][6];				l_cell_reg[14] = inform_L[7][6];				l_cell_reg[15] = inform_L[39][6];				l_cell_reg[16] = inform_L[8][6];				l_cell_reg[17] = inform_L[40][6];				l_cell_reg[18] = inform_L[9][6];				l_cell_reg[19] = inform_L[41][6];				l_cell_reg[20] = inform_L[10][6];				l_cell_reg[21] = inform_L[42][6];				l_cell_reg[22] = inform_L[11][6];				l_cell_reg[23] = inform_L[43][6];				l_cell_reg[24] = inform_L[12][6];				l_cell_reg[25] = inform_L[44][6];				l_cell_reg[26] = inform_L[13][6];				l_cell_reg[27] = inform_L[45][6];				l_cell_reg[28] = inform_L[14][6];				l_cell_reg[29] = inform_L[46][6];				l_cell_reg[30] = inform_L[15][6];				l_cell_reg[31] = inform_L[47][6];				l_cell_reg[32] = inform_L[16][6];				l_cell_reg[33] = inform_L[48][6];				l_cell_reg[34] = inform_L[17][6];				l_cell_reg[35] = inform_L[49][6];				l_cell_reg[36] = inform_L[18][6];				l_cell_reg[37] = inform_L[50][6];				l_cell_reg[38] = inform_L[19][6];				l_cell_reg[39] = inform_L[51][6];				l_cell_reg[40] = inform_L[20][6];				l_cell_reg[41] = inform_L[52][6];				l_cell_reg[42] = inform_L[21][6];				l_cell_reg[43] = inform_L[53][6];				l_cell_reg[44] = inform_L[22][6];				l_cell_reg[45] = inform_L[54][6];				l_cell_reg[46] = inform_L[23][6];				l_cell_reg[47] = inform_L[55][6];				l_cell_reg[48] = inform_L[24][6];				l_cell_reg[49] = inform_L[56][6];				l_cell_reg[50] = inform_L[25][6];				l_cell_reg[51] = inform_L[57][6];				l_cell_reg[52] = inform_L[26][6];				l_cell_reg[53] = inform_L[58][6];				l_cell_reg[54] = inform_L[27][6];				l_cell_reg[55] = inform_L[59][6];				l_cell_reg[56] = inform_L[28][6];				l_cell_reg[57] = inform_L[60][6];				l_cell_reg[58] = inform_L[29][6];				l_cell_reg[59] = inform_L[61][6];				l_cell_reg[60] = inform_L[30][6];				l_cell_reg[61] = inform_L[62][6];				l_cell_reg[62] = inform_L[31][6];				l_cell_reg[63] = inform_L[63][6];				l_cell_reg[64] = inform_L[64][6];				l_cell_reg[65] = inform_L[96][6];				l_cell_reg[66] = inform_L[65][6];				l_cell_reg[67] = inform_L[97][6];				l_cell_reg[68] = inform_L[66][6];				l_cell_reg[69] = inform_L[98][6];				l_cell_reg[70] = inform_L[67][6];				l_cell_reg[71] = inform_L[99][6];				l_cell_reg[72] = inform_L[68][6];				l_cell_reg[73] = inform_L[100][6];				l_cell_reg[74] = inform_L[69][6];				l_cell_reg[75] = inform_L[101][6];				l_cell_reg[76] = inform_L[70][6];				l_cell_reg[77] = inform_L[102][6];				l_cell_reg[78] = inform_L[71][6];				l_cell_reg[79] = inform_L[103][6];				l_cell_reg[80] = inform_L[72][6];				l_cell_reg[81] = inform_L[104][6];				l_cell_reg[82] = inform_L[73][6];				l_cell_reg[83] = inform_L[105][6];				l_cell_reg[84] = inform_L[74][6];				l_cell_reg[85] = inform_L[106][6];				l_cell_reg[86] = inform_L[75][6];				l_cell_reg[87] = inform_L[107][6];				l_cell_reg[88] = inform_L[76][6];				l_cell_reg[89] = inform_L[108][6];				l_cell_reg[90] = inform_L[77][6];				l_cell_reg[91] = inform_L[109][6];				l_cell_reg[92] = inform_L[78][6];				l_cell_reg[93] = inform_L[110][6];				l_cell_reg[94] = inform_L[79][6];				l_cell_reg[95] = inform_L[111][6];				l_cell_reg[96] = inform_L[80][6];				l_cell_reg[97] = inform_L[112][6];				l_cell_reg[98] = inform_L[81][6];				l_cell_reg[99] = inform_L[113][6];				l_cell_reg[100] = inform_L[82][6];				l_cell_reg[101] = inform_L[114][6];				l_cell_reg[102] = inform_L[83][6];				l_cell_reg[103] = inform_L[115][6];				l_cell_reg[104] = inform_L[84][6];				l_cell_reg[105] = inform_L[116][6];				l_cell_reg[106] = inform_L[85][6];				l_cell_reg[107] = inform_L[117][6];				l_cell_reg[108] = inform_L[86][6];				l_cell_reg[109] = inform_L[118][6];				l_cell_reg[110] = inform_L[87][6];				l_cell_reg[111] = inform_L[119][6];				l_cell_reg[112] = inform_L[88][6];				l_cell_reg[113] = inform_L[120][6];				l_cell_reg[114] = inform_L[89][6];				l_cell_reg[115] = inform_L[121][6];				l_cell_reg[116] = inform_L[90][6];				l_cell_reg[117] = inform_L[122][6];				l_cell_reg[118] = inform_L[91][6];				l_cell_reg[119] = inform_L[123][6];				l_cell_reg[120] = inform_L[92][6];				l_cell_reg[121] = inform_L[124][6];				l_cell_reg[122] = inform_L[93][6];				l_cell_reg[123] = inform_L[125][6];				l_cell_reg[124] = inform_L[94][6];				l_cell_reg[125] = inform_L[126][6];				l_cell_reg[126] = inform_L[95][6];				l_cell_reg[127] = inform_L[127][6];			end
			7:			begin				r_cell_reg[0] = inform_R[0][6];				r_cell_reg[1] = inform_R[64][6];				r_cell_reg[2] = inform_R[1][6];				r_cell_reg[3] = inform_R[65][6];				r_cell_reg[4] = inform_R[2][6];				r_cell_reg[5] = inform_R[66][6];				r_cell_reg[6] = inform_R[3][6];				r_cell_reg[7] = inform_R[67][6];				r_cell_reg[8] = inform_R[4][6];				r_cell_reg[9] = inform_R[68][6];				r_cell_reg[10] = inform_R[5][6];				r_cell_reg[11] = inform_R[69][6];				r_cell_reg[12] = inform_R[6][6];				r_cell_reg[13] = inform_R[70][6];				r_cell_reg[14] = inform_R[7][6];				r_cell_reg[15] = inform_R[71][6];				r_cell_reg[16] = inform_R[8][6];				r_cell_reg[17] = inform_R[72][6];				r_cell_reg[18] = inform_R[9][6];				r_cell_reg[19] = inform_R[73][6];				r_cell_reg[20] = inform_R[10][6];				r_cell_reg[21] = inform_R[74][6];				r_cell_reg[22] = inform_R[11][6];				r_cell_reg[23] = inform_R[75][6];				r_cell_reg[24] = inform_R[12][6];				r_cell_reg[25] = inform_R[76][6];				r_cell_reg[26] = inform_R[13][6];				r_cell_reg[27] = inform_R[77][6];				r_cell_reg[28] = inform_R[14][6];				r_cell_reg[29] = inform_R[78][6];				r_cell_reg[30] = inform_R[15][6];				r_cell_reg[31] = inform_R[79][6];				r_cell_reg[32] = inform_R[16][6];				r_cell_reg[33] = inform_R[80][6];				r_cell_reg[34] = inform_R[17][6];				r_cell_reg[35] = inform_R[81][6];				r_cell_reg[36] = inform_R[18][6];				r_cell_reg[37] = inform_R[82][6];				r_cell_reg[38] = inform_R[19][6];				r_cell_reg[39] = inform_R[83][6];				r_cell_reg[40] = inform_R[20][6];				r_cell_reg[41] = inform_R[84][6];				r_cell_reg[42] = inform_R[21][6];				r_cell_reg[43] = inform_R[85][6];				r_cell_reg[44] = inform_R[22][6];				r_cell_reg[45] = inform_R[86][6];				r_cell_reg[46] = inform_R[23][6];				r_cell_reg[47] = inform_R[87][6];				r_cell_reg[48] = inform_R[24][6];				r_cell_reg[49] = inform_R[88][6];				r_cell_reg[50] = inform_R[25][6];				r_cell_reg[51] = inform_R[89][6];				r_cell_reg[52] = inform_R[26][6];				r_cell_reg[53] = inform_R[90][6];				r_cell_reg[54] = inform_R[27][6];				r_cell_reg[55] = inform_R[91][6];				r_cell_reg[56] = inform_R[28][6];				r_cell_reg[57] = inform_R[92][6];				r_cell_reg[58] = inform_R[29][6];				r_cell_reg[59] = inform_R[93][6];				r_cell_reg[60] = inform_R[30][6];				r_cell_reg[61] = inform_R[94][6];				r_cell_reg[62] = inform_R[31][6];				r_cell_reg[63] = inform_R[95][6];				r_cell_reg[64] = inform_R[32][6];				r_cell_reg[65] = inform_R[96][6];				r_cell_reg[66] = inform_R[33][6];				r_cell_reg[67] = inform_R[97][6];				r_cell_reg[68] = inform_R[34][6];				r_cell_reg[69] = inform_R[98][6];				r_cell_reg[70] = inform_R[35][6];				r_cell_reg[71] = inform_R[99][6];				r_cell_reg[72] = inform_R[36][6];				r_cell_reg[73] = inform_R[100][6];				r_cell_reg[74] = inform_R[37][6];				r_cell_reg[75] = inform_R[101][6];				r_cell_reg[76] = inform_R[38][6];				r_cell_reg[77] = inform_R[102][6];				r_cell_reg[78] = inform_R[39][6];				r_cell_reg[79] = inform_R[103][6];				r_cell_reg[80] = inform_R[40][6];				r_cell_reg[81] = inform_R[104][6];				r_cell_reg[82] = inform_R[41][6];				r_cell_reg[83] = inform_R[105][6];				r_cell_reg[84] = inform_R[42][6];				r_cell_reg[85] = inform_R[106][6];				r_cell_reg[86] = inform_R[43][6];				r_cell_reg[87] = inform_R[107][6];				r_cell_reg[88] = inform_R[44][6];				r_cell_reg[89] = inform_R[108][6];				r_cell_reg[90] = inform_R[45][6];				r_cell_reg[91] = inform_R[109][6];				r_cell_reg[92] = inform_R[46][6];				r_cell_reg[93] = inform_R[110][6];				r_cell_reg[94] = inform_R[47][6];				r_cell_reg[95] = inform_R[111][6];				r_cell_reg[96] = inform_R[48][6];				r_cell_reg[97] = inform_R[112][6];				r_cell_reg[98] = inform_R[49][6];				r_cell_reg[99] = inform_R[113][6];				r_cell_reg[100] = inform_R[50][6];				r_cell_reg[101] = inform_R[114][6];				r_cell_reg[102] = inform_R[51][6];				r_cell_reg[103] = inform_R[115][6];				r_cell_reg[104] = inform_R[52][6];				r_cell_reg[105] = inform_R[116][6];				r_cell_reg[106] = inform_R[53][6];				r_cell_reg[107] = inform_R[117][6];				r_cell_reg[108] = inform_R[54][6];				r_cell_reg[109] = inform_R[118][6];				r_cell_reg[110] = inform_R[55][6];				r_cell_reg[111] = inform_R[119][6];				r_cell_reg[112] = inform_R[56][6];				r_cell_reg[113] = inform_R[120][6];				r_cell_reg[114] = inform_R[57][6];				r_cell_reg[115] = inform_R[121][6];				r_cell_reg[116] = inform_R[58][6];				r_cell_reg[117] = inform_R[122][6];				r_cell_reg[118] = inform_R[59][6];				r_cell_reg[119] = inform_R[123][6];				r_cell_reg[120] = inform_R[60][6];				r_cell_reg[121] = inform_R[124][6];				r_cell_reg[122] = inform_R[61][6];				r_cell_reg[123] = inform_R[125][6];				r_cell_reg[124] = inform_R[62][6];				r_cell_reg[125] = inform_R[126][6];				r_cell_reg[126] = inform_R[63][6];				r_cell_reg[127] = inform_R[127][6];				l_cell_reg[0] = inform_L[0][7];				l_cell_reg[1] = inform_L[64][7];				l_cell_reg[2] = inform_L[1][7];				l_cell_reg[3] = inform_L[65][7];				l_cell_reg[4] = inform_L[2][7];				l_cell_reg[5] = inform_L[66][7];				l_cell_reg[6] = inform_L[3][7];				l_cell_reg[7] = inform_L[67][7];				l_cell_reg[8] = inform_L[4][7];				l_cell_reg[9] = inform_L[68][7];				l_cell_reg[10] = inform_L[5][7];				l_cell_reg[11] = inform_L[69][7];				l_cell_reg[12] = inform_L[6][7];				l_cell_reg[13] = inform_L[70][7];				l_cell_reg[14] = inform_L[7][7];				l_cell_reg[15] = inform_L[71][7];				l_cell_reg[16] = inform_L[8][7];				l_cell_reg[17] = inform_L[72][7];				l_cell_reg[18] = inform_L[9][7];				l_cell_reg[19] = inform_L[73][7];				l_cell_reg[20] = inform_L[10][7];				l_cell_reg[21] = inform_L[74][7];				l_cell_reg[22] = inform_L[11][7];				l_cell_reg[23] = inform_L[75][7];				l_cell_reg[24] = inform_L[12][7];				l_cell_reg[25] = inform_L[76][7];				l_cell_reg[26] = inform_L[13][7];				l_cell_reg[27] = inform_L[77][7];				l_cell_reg[28] = inform_L[14][7];				l_cell_reg[29] = inform_L[78][7];				l_cell_reg[30] = inform_L[15][7];				l_cell_reg[31] = inform_L[79][7];				l_cell_reg[32] = inform_L[16][7];				l_cell_reg[33] = inform_L[80][7];				l_cell_reg[34] = inform_L[17][7];				l_cell_reg[35] = inform_L[81][7];				l_cell_reg[36] = inform_L[18][7];				l_cell_reg[37] = inform_L[82][7];				l_cell_reg[38] = inform_L[19][7];				l_cell_reg[39] = inform_L[83][7];				l_cell_reg[40] = inform_L[20][7];				l_cell_reg[41] = inform_L[84][7];				l_cell_reg[42] = inform_L[21][7];				l_cell_reg[43] = inform_L[85][7];				l_cell_reg[44] = inform_L[22][7];				l_cell_reg[45] = inform_L[86][7];				l_cell_reg[46] = inform_L[23][7];				l_cell_reg[47] = inform_L[87][7];				l_cell_reg[48] = inform_L[24][7];				l_cell_reg[49] = inform_L[88][7];				l_cell_reg[50] = inform_L[25][7];				l_cell_reg[51] = inform_L[89][7];				l_cell_reg[52] = inform_L[26][7];				l_cell_reg[53] = inform_L[90][7];				l_cell_reg[54] = inform_L[27][7];				l_cell_reg[55] = inform_L[91][7];				l_cell_reg[56] = inform_L[28][7];				l_cell_reg[57] = inform_L[92][7];				l_cell_reg[58] = inform_L[29][7];				l_cell_reg[59] = inform_L[93][7];				l_cell_reg[60] = inform_L[30][7];				l_cell_reg[61] = inform_L[94][7];				l_cell_reg[62] = inform_L[31][7];				l_cell_reg[63] = inform_L[95][7];				l_cell_reg[64] = inform_L[32][7];				l_cell_reg[65] = inform_L[96][7];				l_cell_reg[66] = inform_L[33][7];				l_cell_reg[67] = inform_L[97][7];				l_cell_reg[68] = inform_L[34][7];				l_cell_reg[69] = inform_L[98][7];				l_cell_reg[70] = inform_L[35][7];				l_cell_reg[71] = inform_L[99][7];				l_cell_reg[72] = inform_L[36][7];				l_cell_reg[73] = inform_L[100][7];				l_cell_reg[74] = inform_L[37][7];				l_cell_reg[75] = inform_L[101][7];				l_cell_reg[76] = inform_L[38][7];				l_cell_reg[77] = inform_L[102][7];				l_cell_reg[78] = inform_L[39][7];				l_cell_reg[79] = inform_L[103][7];				l_cell_reg[80] = inform_L[40][7];				l_cell_reg[81] = inform_L[104][7];				l_cell_reg[82] = inform_L[41][7];				l_cell_reg[83] = inform_L[105][7];				l_cell_reg[84] = inform_L[42][7];				l_cell_reg[85] = inform_L[106][7];				l_cell_reg[86] = inform_L[43][7];				l_cell_reg[87] = inform_L[107][7];				l_cell_reg[88] = inform_L[44][7];				l_cell_reg[89] = inform_L[108][7];				l_cell_reg[90] = inform_L[45][7];				l_cell_reg[91] = inform_L[109][7];				l_cell_reg[92] = inform_L[46][7];				l_cell_reg[93] = inform_L[110][7];				l_cell_reg[94] = inform_L[47][7];				l_cell_reg[95] = inform_L[111][7];				l_cell_reg[96] = inform_L[48][7];				l_cell_reg[97] = inform_L[112][7];				l_cell_reg[98] = inform_L[49][7];				l_cell_reg[99] = inform_L[113][7];				l_cell_reg[100] = inform_L[50][7];				l_cell_reg[101] = inform_L[114][7];				l_cell_reg[102] = inform_L[51][7];				l_cell_reg[103] = inform_L[115][7];				l_cell_reg[104] = inform_L[52][7];				l_cell_reg[105] = inform_L[116][7];				l_cell_reg[106] = inform_L[53][7];				l_cell_reg[107] = inform_L[117][7];				l_cell_reg[108] = inform_L[54][7];				l_cell_reg[109] = inform_L[118][7];				l_cell_reg[110] = inform_L[55][7];				l_cell_reg[111] = inform_L[119][7];				l_cell_reg[112] = inform_L[56][7];				l_cell_reg[113] = inform_L[120][7];				l_cell_reg[114] = inform_L[57][7];				l_cell_reg[115] = inform_L[121][7];				l_cell_reg[116] = inform_L[58][7];				l_cell_reg[117] = inform_L[122][7];				l_cell_reg[118] = inform_L[59][7];				l_cell_reg[119] = inform_L[123][7];				l_cell_reg[120] = inform_L[60][7];				l_cell_reg[121] = inform_L[124][7];				l_cell_reg[122] = inform_L[61][7];				l_cell_reg[123] = inform_L[125][7];				l_cell_reg[124] = inform_L[62][7];				l_cell_reg[125] = inform_L[126][7];				l_cell_reg[126] = inform_L[63][7];				l_cell_reg[127] = inform_L[127][7];			end
			default:			begin					r_cell_reg[0] <= 0;					r_cell_reg[1] <= 0;					r_cell_reg[2] <= 0;					r_cell_reg[3] <= 0;					r_cell_reg[4] <= 0;					r_cell_reg[5] <= 0;					r_cell_reg[6] <= 0;					r_cell_reg[7] <= 0;					r_cell_reg[8] <= 0;					r_cell_reg[9] <= 0;					r_cell_reg[10] <= 0;					r_cell_reg[11] <= 0;					r_cell_reg[12] <= 0;					r_cell_reg[13] <= 0;					r_cell_reg[14] <= 0;					r_cell_reg[15] <= 0;					r_cell_reg[16] <= 0;					r_cell_reg[17] <= 0;					r_cell_reg[18] <= 0;					r_cell_reg[19] <= 0;					r_cell_reg[20] <= 0;					r_cell_reg[21] <= 0;					r_cell_reg[22] <= 0;					r_cell_reg[23] <= 0;					r_cell_reg[24] <= 0;					r_cell_reg[25] <= 0;					r_cell_reg[26] <= 0;					r_cell_reg[27] <= 0;					r_cell_reg[28] <= 0;					r_cell_reg[29] <= 0;					r_cell_reg[30] <= 0;					r_cell_reg[31] <= 0;					r_cell_reg[32] <= 0;					r_cell_reg[33] <= 0;					r_cell_reg[34] <= 0;					r_cell_reg[35] <= 0;					r_cell_reg[36] <= 0;					r_cell_reg[37] <= 0;					r_cell_reg[38] <= 0;					r_cell_reg[39] <= 0;					r_cell_reg[40] <= 0;					r_cell_reg[41] <= 0;					r_cell_reg[42] <= 0;					r_cell_reg[43] <= 0;					r_cell_reg[44] <= 0;					r_cell_reg[45] <= 0;					r_cell_reg[46] <= 0;					r_cell_reg[47] <= 0;					r_cell_reg[48] <= 0;					r_cell_reg[49] <= 0;					r_cell_reg[50] <= 0;					r_cell_reg[51] <= 0;					r_cell_reg[52] <= 0;					r_cell_reg[53] <= 0;					r_cell_reg[54] <= 0;					r_cell_reg[55] <= 0;					r_cell_reg[56] <= 0;					r_cell_reg[57] <= 0;					r_cell_reg[58] <= 0;					r_cell_reg[59] <= 0;					r_cell_reg[60] <= 0;					r_cell_reg[61] <= 0;					r_cell_reg[62] <= 0;					r_cell_reg[63] <= 0;					r_cell_reg[64] <= 0;					r_cell_reg[65] <= 0;					r_cell_reg[66] <= 0;					r_cell_reg[67] <= 0;					r_cell_reg[68] <= 0;					r_cell_reg[69] <= 0;					r_cell_reg[70] <= 0;					r_cell_reg[71] <= 0;					r_cell_reg[72] <= 0;					r_cell_reg[73] <= 0;					r_cell_reg[74] <= 0;					r_cell_reg[75] <= 0;					r_cell_reg[76] <= 0;					r_cell_reg[77] <= 0;					r_cell_reg[78] <= 0;					r_cell_reg[79] <= 0;					r_cell_reg[80] <= 0;					r_cell_reg[81] <= 0;					r_cell_reg[82] <= 0;					r_cell_reg[83] <= 0;					r_cell_reg[84] <= 0;					r_cell_reg[85] <= 0;					r_cell_reg[86] <= 0;					r_cell_reg[87] <= 0;					r_cell_reg[88] <= 0;					r_cell_reg[89] <= 0;					r_cell_reg[90] <= 0;					r_cell_reg[91] <= 0;					r_cell_reg[92] <= 0;					r_cell_reg[93] <= 0;					r_cell_reg[94] <= 0;					r_cell_reg[95] <= 0;					r_cell_reg[96] <= 0;					r_cell_reg[97] <= 0;					r_cell_reg[98] <= 0;					r_cell_reg[99] <= 0;					r_cell_reg[100] <= 0;					r_cell_reg[101] <= 0;					r_cell_reg[102] <= 0;					r_cell_reg[103] <= 0;					r_cell_reg[104] <= 0;					r_cell_reg[105] <= 0;					r_cell_reg[106] <= 0;					r_cell_reg[107] <= 0;					r_cell_reg[108] <= 0;					r_cell_reg[109] <= 0;					r_cell_reg[110] <= 0;					r_cell_reg[111] <= 0;					r_cell_reg[112] <= 0;					r_cell_reg[113] <= 0;					r_cell_reg[114] <= 0;					r_cell_reg[115] <= 0;					r_cell_reg[116] <= 0;					r_cell_reg[117] <= 0;					r_cell_reg[118] <= 0;					r_cell_reg[119] <= 0;					r_cell_reg[120] <= 0;					r_cell_reg[121] <= 0;					r_cell_reg[122] <= 0;					r_cell_reg[123] <= 0;					r_cell_reg[124] <= 0;					r_cell_reg[125] <= 0;					r_cell_reg[126] <= 0;					r_cell_reg[127] <= 0;					l_cell_reg[0] <= 0;					l_cell_reg[1] <= 0;					l_cell_reg[2] <= 0;					l_cell_reg[3] <= 0;					l_cell_reg[4] <= 0;					l_cell_reg[5] <= 0;					l_cell_reg[6] <= 0;					l_cell_reg[7] <= 0;					l_cell_reg[8] <= 0;					l_cell_reg[9] <= 0;					l_cell_reg[10] <= 0;					l_cell_reg[11] <= 0;					l_cell_reg[12] <= 0;					l_cell_reg[13] <= 0;					l_cell_reg[14] <= 0;					l_cell_reg[15] <= 0;					l_cell_reg[16] <= 0;					l_cell_reg[17] <= 0;					l_cell_reg[18] <= 0;					l_cell_reg[19] <= 0;					l_cell_reg[20] <= 0;					l_cell_reg[21] <= 0;					l_cell_reg[22] <= 0;					l_cell_reg[23] <= 0;					l_cell_reg[24] <= 0;					l_cell_reg[25] <= 0;					l_cell_reg[26] <= 0;					l_cell_reg[27] <= 0;					l_cell_reg[28] <= 0;					l_cell_reg[29] <= 0;					l_cell_reg[30] <= 0;					l_cell_reg[31] <= 0;					l_cell_reg[32] <= 0;					l_cell_reg[33] <= 0;					l_cell_reg[34] <= 0;					l_cell_reg[35] <= 0;					l_cell_reg[36] <= 0;					l_cell_reg[37] <= 0;					l_cell_reg[38] <= 0;					l_cell_reg[39] <= 0;					l_cell_reg[40] <= 0;					l_cell_reg[41] <= 0;					l_cell_reg[42] <= 0;					l_cell_reg[43] <= 0;					l_cell_reg[44] <= 0;					l_cell_reg[45] <= 0;					l_cell_reg[46] <= 0;					l_cell_reg[47] <= 0;					l_cell_reg[48] <= 0;					l_cell_reg[49] <= 0;					l_cell_reg[50] <= 0;					l_cell_reg[51] <= 0;					l_cell_reg[52] <= 0;					l_cell_reg[53] <= 0;					l_cell_reg[54] <= 0;					l_cell_reg[55] <= 0;					l_cell_reg[56] <= 0;					l_cell_reg[57] <= 0;					l_cell_reg[58] <= 0;					l_cell_reg[59] <= 0;					l_cell_reg[60] <= 0;					l_cell_reg[61] <= 0;					l_cell_reg[62] <= 0;					l_cell_reg[63] <= 0;					l_cell_reg[64] <= 0;					l_cell_reg[65] <= 0;					l_cell_reg[66] <= 0;					l_cell_reg[67] <= 0;					l_cell_reg[68] <= 0;					l_cell_reg[69] <= 0;					l_cell_reg[70] <= 0;					l_cell_reg[71] <= 0;					l_cell_reg[72] <= 0;					l_cell_reg[73] <= 0;					l_cell_reg[74] <= 0;					l_cell_reg[75] <= 0;					l_cell_reg[76] <= 0;					l_cell_reg[77] <= 0;					l_cell_reg[78] <= 0;					l_cell_reg[79] <= 0;					l_cell_reg[80] <= 0;					l_cell_reg[81] <= 0;					l_cell_reg[82] <= 0;					l_cell_reg[83] <= 0;					l_cell_reg[84] <= 0;					l_cell_reg[85] <= 0;					l_cell_reg[86] <= 0;					l_cell_reg[87] <= 0;					l_cell_reg[88] <= 0;					l_cell_reg[89] <= 0;					l_cell_reg[90] <= 0;					l_cell_reg[91] <= 0;					l_cell_reg[92] <= 0;					l_cell_reg[93] <= 0;					l_cell_reg[94] <= 0;					l_cell_reg[95] <= 0;					l_cell_reg[96] <= 0;					l_cell_reg[97] <= 0;					l_cell_reg[98] <= 0;					l_cell_reg[99] <= 0;					l_cell_reg[100] <= 0;					l_cell_reg[101] <= 0;					l_cell_reg[102] <= 0;					l_cell_reg[103] <= 0;					l_cell_reg[104] <= 0;					l_cell_reg[105] <= 0;					l_cell_reg[106] <= 0;					l_cell_reg[107] <= 0;					l_cell_reg[108] <= 0;					l_cell_reg[109] <= 0;					l_cell_reg[110] <= 0;					l_cell_reg[111] <= 0;					l_cell_reg[112] <= 0;					l_cell_reg[113] <= 0;					l_cell_reg[114] <= 0;					l_cell_reg[115] <= 0;					l_cell_reg[116] <= 0;					l_cell_reg[117] <= 0;					l_cell_reg[118] <= 0;					l_cell_reg[119] <= 0;					l_cell_reg[120] <= 0;					l_cell_reg[121] <= 0;					l_cell_reg[122] <= 0;					l_cell_reg[123] <= 0;					l_cell_reg[124] <= 0;					l_cell_reg[125] <= 0;					l_cell_reg[126] <= 0;					l_cell_reg[127] <= 0;			end
		endcase	end
	genvar i;	generate		for (i = 0; i < 128 ; i = i+2)			begin :bp_2				bp_2_cell fun(					.clk(clk),					.en(1),					.R_IN1(r_cell_reg[i]),					.R_IN2(r_cell_reg[i+1]),					.L_IN1(l_cell_reg[i]),					.L_IN2(l_cell_reg[i+1]),					.R_OUT1(r_cell_wire[i]),					.R_OUT2(r_cell_wire[i+1]),					.L_OUT1(l_cell_wire[i]),					.L_OUT2(l_cell_wire[i+1])				);			end	endgenerate
	always @(posedge clk) begin		if (bp_over_flag) begin			OUT_1 <= inform_L [0][0] ;			OUT_2 <= inform_L [1][0] ;			OUT_3 <= inform_L [2][0] ;			OUT_4 <= inform_L [3][0] ;			OUT_5 <= inform_L [4][0] ;			OUT_6 <= inform_L [5][0] ;			OUT_7 <= inform_L [6][0] ;			OUT_8 <= inform_L [7][0] ;			OUT_9 <= inform_L [8][0] ;			OUT_10 <= inform_L [9][0] ;			OUT_11 <= inform_L [10][0] ;			OUT_12 <= inform_L [11][0] ;			OUT_13 <= inform_L [12][0] ;			OUT_14 <= inform_L [13][0] ;			OUT_15 <= inform_L [14][0] ;			OUT_16 <= inform_L [15][0] ;			OUT_17 <= inform_L [16][0] ;			OUT_18 <= inform_L [17][0] ;			OUT_19 <= inform_L [18][0] ;			OUT_20 <= inform_L [19][0] ;			OUT_21 <= inform_L [20][0] ;			OUT_22 <= inform_L [21][0] ;			OUT_23 <= inform_L [22][0] ;			OUT_24 <= inform_L [23][0] ;			OUT_25 <= inform_L [24][0] ;			OUT_26 <= inform_L [25][0] ;			OUT_27 <= inform_L [26][0] ;			OUT_28 <= inform_L [27][0] ;			OUT_29 <= inform_L [28][0] ;			OUT_30 <= inform_L [29][0] ;			OUT_31 <= inform_L [30][0] ;			OUT_32 <= inform_L [31][0] ;			OUT_33 <= inform_L [32][0] ;			OUT_34 <= inform_L [33][0] ;			OUT_35 <= inform_L [34][0] ;			OUT_36 <= inform_L [35][0] ;			OUT_37 <= inform_L [36][0] ;			OUT_38 <= inform_L [37][0] ;			OUT_39 <= inform_L [38][0] ;			OUT_40 <= inform_L [39][0] ;			OUT_41 <= inform_L [40][0] ;			OUT_42 <= inform_L [41][0] ;			OUT_43 <= inform_L [42][0] ;			OUT_44 <= inform_L [43][0] ;			OUT_45 <= inform_L [44][0] ;			OUT_46 <= inform_L [45][0] ;			OUT_47 <= inform_L [46][0] ;			OUT_48 <= inform_L [47][0] ;			OUT_49 <= inform_L [48][0] ;			OUT_50 <= inform_L [49][0] ;			OUT_51 <= inform_L [50][0] ;			OUT_52 <= inform_L [51][0] ;			OUT_53 <= inform_L [52][0] ;			OUT_54 <= inform_L [53][0] ;			OUT_55 <= inform_L [54][0] ;			OUT_56 <= inform_L [55][0] ;			OUT_57 <= inform_L [56][0] ;			OUT_58 <= inform_L [57][0] ;			OUT_59 <= inform_L [58][0] ;			OUT_60 <= inform_L [59][0] ;			OUT_61 <= inform_L [60][0] ;			OUT_62 <= inform_L [61][0] ;			OUT_63 <= inform_L [62][0] ;			OUT_64 <= inform_L [63][0] ;			OUT_65 <= inform_L [64][0] ;			OUT_66 <= inform_L [65][0] ;			OUT_67 <= inform_L [66][0] ;			OUT_68 <= inform_L [67][0] ;			OUT_69 <= inform_L [68][0] ;			OUT_70 <= inform_L [69][0] ;			OUT_71 <= inform_L [70][0] ;			OUT_72 <= inform_L [71][0] ;			OUT_73 <= inform_L [72][0] ;			OUT_74 <= inform_L [73][0] ;			OUT_75 <= inform_L [74][0] ;			OUT_76 <= inform_L [75][0] ;			OUT_77 <= inform_L [76][0] ;			OUT_78 <= inform_L [77][0] ;			OUT_79 <= inform_L [78][0] ;			OUT_80 <= inform_L [79][0] ;			OUT_81 <= inform_L [80][0] ;			OUT_82 <= inform_L [81][0] ;			OUT_83 <= inform_L [82][0] ;			OUT_84 <= inform_L [83][0] ;			OUT_85 <= inform_L [84][0] ;			OUT_86 <= inform_L [85][0] ;			OUT_87 <= inform_L [86][0] ;			OUT_88 <= inform_L [87][0] ;			OUT_89 <= inform_L [88][0] ;			OUT_90 <= inform_L [89][0] ;			OUT_91 <= inform_L [90][0] ;			OUT_92 <= inform_L [91][0] ;			OUT_93 <= inform_L [92][0] ;			OUT_94 <= inform_L [93][0] ;			OUT_95 <= inform_L [94][0] ;			OUT_96 <= inform_L [95][0] ;			OUT_97 <= inform_L [96][0] ;			OUT_98 <= inform_L [97][0] ;			OUT_99 <= inform_L [98][0] ;			OUT_100 <= inform_L [99][0] ;			OUT_101 <= inform_L [100][0] ;			OUT_102 <= inform_L [101][0] ;			OUT_103 <= inform_L [102][0] ;			OUT_104 <= inform_L [103][0] ;			OUT_105 <= inform_L [104][0] ;			OUT_106 <= inform_L [105][0] ;			OUT_107 <= inform_L [106][0] ;			OUT_108 <= inform_L [107][0] ;			OUT_109 <= inform_L [108][0] ;			OUT_110 <= inform_L [109][0] ;			OUT_111 <= inform_L [110][0] ;			OUT_112 <= inform_L [111][0] ;			OUT_113 <= inform_L [112][0] ;			OUT_114 <= inform_L [113][0] ;			OUT_115 <= inform_L [114][0] ;			OUT_116 <= inform_L [115][0] ;			OUT_117 <= inform_L [116][0] ;			OUT_118 <= inform_L [117][0] ;			OUT_119 <= inform_L [118][0] ;			OUT_120 <= inform_L [119][0] ;			OUT_121 <= inform_L [120][0] ;			OUT_122 <= inform_L [121][0] ;			OUT_123 <= inform_L [122][0] ;			OUT_124 <= inform_L [123][0] ;			OUT_125 <= inform_L [124][0] ;			OUT_126 <= inform_L [125][0] ;			OUT_127 <= inform_L [126][0] ;			OUT_128 <= inform_L [127][0] ;		end	end
endmodule